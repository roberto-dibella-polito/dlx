
module DLX ( CLK, RST, IRAM_ADDRESS, IRAM_ISSUE, IRAM_READY, IRAM_DATA, 
        DRAM_ADDRESS, DRAM_ISSUE, DRAM_READNOTWRITE, DRAM_READY, DRAM_DATA );
  output [31:0] IRAM_ADDRESS;
  input [31:0] IRAM_DATA;
  output [31:0] DRAM_ADDRESS;
  inout [31:0] DRAM_DATA;
  input CLK, RST, IRAM_READY, DRAM_READY;
  output IRAM_ISSUE, DRAM_ISSUE, DRAM_READNOTWRITE;
  wire   pipe_if_id_en_i, pipe_ex_mem_en_i, pipe_clear_n_i, rf_spill_i,
         rf_fill_i, rf_rs1_en_i, rf_rs2_en_i, imm_isoff_i, imm_uns_i,
         reg31_sel_i, regrd_sel_i, muxA_sel_i, muxB_sel_i, is_zero_i,
         mem_in_en_i, npc_wb_en_i, jump_en_i, wb_mux_sel_i, rf_we_i, CU_I_n291,
         CU_I_n290, CU_I_n289, CU_I_n288, CU_I_n287, CU_I_n286, CU_I_n285,
         CU_I_n284, CU_I_n283, CU_I_n282, CU_I_n281, CU_I_n280, CU_I_n279,
         CU_I_n278, CU_I_n277, CU_I_n276, CU_I_n275, CU_I_n274, CU_I_n273,
         CU_I_n272, CU_I_n271, CU_I_n270, CU_I_n269, CU_I_n268, CU_I_n267,
         CU_I_n266, CU_I_n265, CU_I_n264, CU_I_n263, CU_I_n262, CU_I_n261,
         CU_I_n260, CU_I_n259, CU_I_n258, CU_I_n257, CU_I_n256, CU_I_n76,
         CU_I_n75, CU_I_n74, CU_I_n73, CU_I_n72, CU_I_n71, CU_I_n70, CU_I_n69,
         CU_I_n68, CU_I_n67, CU_I_n66, CU_I_n65, CU_I_n64, CU_I_n63, CU_I_n60,
         CU_I_n59, CU_I_n58, CU_I_n57, CU_I_n56, CU_I_n55, CU_I_n54, CU_I_n53,
         CU_I_n52, CU_I_n51, CU_I_n50, CU_I_n49, CU_I_n48, CU_I_n47, CU_I_n45,
         CU_I_n43, CU_I_n42, CU_I_n41, CU_I_n39, CU_I_n38, CU_I_n29, CU_I_n28,
         CU_I_n26, CU_I_n25, CU_I_n24, CU_I_n20, CU_I_n18, CU_I_n14, CU_I_n1,
         CU_I_n254, CU_I_n253, CU_I_n252, CU_I_n251, CU_I_n250, CU_I_n249,
         CU_I_n248, CU_I_n247, CU_I_n246, CU_I_n245, CU_I_n244, CU_I_n243,
         CU_I_n242, CU_I_n241, CU_I_n240, CU_I_n239, CU_I_n238, CU_I_n237,
         CU_I_n236, CU_I_n235, CU_I_n234, CU_I_n233, CU_I_n232, CU_I_n231,
         CU_I_n230, CU_I_n229, CU_I_n228, CU_I_n227, CU_I_n226, CU_I_n225,
         CU_I_n224, CU_I_n223, CU_I_n222, CU_I_n221, CU_I_n220, CU_I_n219,
         CU_I_n218, CU_I_n217, CU_I_n216, CU_I_n215, CU_I_n214, CU_I_n213,
         CU_I_n212, CU_I_n211, CU_I_n210, CU_I_n209, CU_I_n208, CU_I_n207,
         CU_I_n206, CU_I_n205, CU_I_n204, CU_I_n203, CU_I_n202, CU_I_n201,
         CU_I_n200, CU_I_n199, CU_I_n198, CU_I_n197, CU_I_n196, CU_I_n195,
         CU_I_n194, CU_I_n193, CU_I_n192, CU_I_n191, CU_I_n190, CU_I_n189,
         CU_I_n188, CU_I_n187, CU_I_n186, CU_I_n185, CU_I_n184, CU_I_n183,
         CU_I_n182, CU_I_n181, CU_I_n180, CU_I_n179, CU_I_n178, CU_I_n177,
         CU_I_n176, CU_I_n175, CU_I_n174, CU_I_n173, CU_I_n172, CU_I_n171,
         CU_I_n170, CU_I_n169, CU_I_n168, CU_I_n167, CU_I_n166, CU_I_n165,
         CU_I_n164, CU_I_n163, CU_I_n162, CU_I_n161, CU_I_n160, CU_I_n159,
         CU_I_n158, CU_I_n157, CU_I_n156, CU_I_n155, CU_I_n154, CU_I_n153,
         CU_I_n152, CU_I_n151, CU_I_n150, CU_I_n149, CU_I_n148, CU_I_n147,
         CU_I_n146, CU_I_n145, CU_I_n144, CU_I_n143, CU_I_n142, CU_I_n141,
         CU_I_n140, CU_I_n139, CU_I_n138, CU_I_n137, CU_I_n136, CU_I_n135,
         CU_I_n134, CU_I_n133, CU_I_n132, CU_I_n131, CU_I_n130, CU_I_n129,
         CU_I_n128, CU_I_n127, CU_I_n126, CU_I_n125, CU_I_n124, CU_I_n123,
         CU_I_n122, CU_I_n121, CU_I_n120, CU_I_n119, CU_I_n118, CU_I_n117,
         CU_I_n116, CU_I_n115, CU_I_n114, CU_I_n113, CU_I_n112, CU_I_n111,
         CU_I_n110, CU_I_n109, CU_I_n108, CU_I_n107, CU_I_n106, CU_I_n105,
         CU_I_n104, CU_I_n103, CU_I_n102, CU_I_n101, CU_I_n100, CU_I_n99,
         CU_I_n98, CU_I_n97, CU_I_n96, CU_I_n95, CU_I_n94, CU_I_n93, CU_I_n92,
         CU_I_n91, CU_I_n90, CU_I_n89, CU_I_n88, CU_I_n87, CU_I_n86, CU_I_n85,
         CU_I_n84, CU_I_n83, CU_I_n82, CU_I_n81, CU_I_n80, CU_I_n79, CU_I_n78,
         CU_I_n77, CU_I_n37, CU_I_n36, CU_I_n35, CU_I_n34, CU_I_n33, CU_I_n32,
         CU_I_n31, CU_I_n30, CU_I_n27, CU_I_n23, CU_I_n22, CU_I_n21, CU_I_n19,
         CU_I_n17, CU_I_n16, CU_I_n15, CU_I_n13, CU_I_n12, CU_I_n11, CU_I_n10,
         CU_I_n9, CU_I_n8, CU_I_n7, CU_I_n6, CU_I_n5, CU_I_n4, CU_I_n3,
         CU_I_n2, CU_I_cw3_4_, CU_I_cw3_5_, CU_I_cw1_1_, CU_I_n294, CU_I_n293,
         CU_I_n292, dp_n1055, dp_n1054, dp_n1053, dp_n1052, dp_n1051, dp_n1050,
         dp_n1049, dp_n1048, dp_n1047, dp_n1046, dp_n1045, dp_n1044, dp_n1043,
         dp_n1042, dp_n1041, dp_n1040, dp_n1039, dp_n1038, dp_n1037, dp_n1036,
         dp_n1035, dp_n1034, dp_n1033, dp_n1032, dp_n1031, dp_n1030, dp_n1029,
         dp_n1028, dp_n1027, dp_n1026, dp_n1025, dp_n1024, dp_n1023, dp_n1022,
         dp_n1021, dp_n1020, dp_n1019, dp_n1018, dp_n1017, dp_n1016, dp_n648,
         dp_n647, dp_n646, dp_n645, dp_n644, dp_n643, dp_n642, dp_n641,
         dp_n640, dp_n639, dp_n638, dp_n637, dp_n636, dp_n635, dp_n634,
         dp_n633, dp_n632, dp_n631, dp_n630, dp_n629, dp_n628, dp_n627,
         dp_n626, dp_n625, dp_n624, dp_n623, dp_n622, dp_n621, dp_n620,
         dp_n619, dp_n618, dp_n617, dp_n616, dp_n615, dp_n614, dp_n613,
         dp_n612, dp_n611, dp_n610, dp_n609, dp_n608, dp_n607, dp_n606,
         dp_n605, dp_n604, dp_n603, dp_n602, dp_n601, dp_n600, dp_n599,
         dp_n598, dp_n597, dp_n596, dp_n595, dp_n594, dp_n593, dp_n592,
         dp_n591, dp_n590, dp_n589, dp_n588, dp_n587, dp_n586, dp_n585,
         dp_n584, dp_n525, dp_n523, dp_n521, dp_n519, dp_n517, dp_n413,
         dp_n412, dp_n411, dp_n410, dp_n409, dp_n408, dp_n407, dp_n406,
         dp_n405, dp_n404, dp_n403, dp_n402, dp_n334, dp_n333, dp_n332,
         dp_n331, dp_n330, dp_n329, dp_n328, dp_n327, dp_n326, dp_n325,
         dp_n324, dp_n323, dp_n322, dp_n321, dp_n320, dp_n319, dp_n318,
         dp_n317, dp_n316, dp_n315, dp_n314, dp_n313, dp_n312, dp_n311,
         dp_n310, dp_n309, dp_n308, dp_n307, dp_n306, dp_n305, dp_n304,
         dp_n303, dp_n300, dp_n299, dp_n298, dp_n297, dp_n296, dp_n295,
         dp_n294, dp_n293, dp_n292, dp_n291, dp_n290, dp_n289, dp_n288,
         dp_n287, dp_n286, dp_n285, dp_n284, dp_n283, dp_n282, dp_n281,
         dp_n280, dp_n279, dp_n278, dp_n277, dp_n276, dp_n275, dp_n274,
         dp_n273, dp_n272, dp_n271, dp_n270, dp_n269, dp_n268, dp_n267,
         dp_n266, dp_n265, dp_n264, dp_n263, dp_n262, dp_n261, dp_n260,
         dp_n259, dp_n258, dp_n257, dp_n256, dp_n255, dp_n254, dp_n253,
         dp_n252, dp_n251, dp_n250, dp_n249, dp_n248, dp_n247, dp_n246,
         dp_n245, dp_n244, dp_n243, dp_n242, dp_n241, dp_n240, dp_n239,
         dp_n238, dp_n237, dp_n236, dp_n235, dp_n234, dp_n233, dp_n232,
         dp_n231, dp_n230, dp_n229, dp_n228, dp_n227, dp_n226, dp_n225,
         dp_n224, dp_n223, dp_n222, dp_n221, dp_n220, dp_n219, dp_n218,
         dp_n217, dp_n216, dp_n215, dp_n214, dp_n213, dp_n212, dp_n211,
         dp_n210, dp_n209, dp_n208, dp_n207, dp_n206, dp_n205, dp_n204,
         dp_n203, dp_n202, dp_n201, dp_n200, dp_n199, dp_n198, dp_n197,
         dp_n196, dp_n195, dp_n194, dp_n193, dp_n192, dp_n191, dp_n190,
         dp_n189, dp_n188, dp_n187, dp_n186, dp_n185, dp_n184, dp_n183,
         dp_n182, dp_n181, dp_n180, dp_n179, dp_n178, dp_n177, dp_n176,
         dp_n175, dp_n174, dp_n173, dp_n172, dp_n171, dp_n170, dp_n169,
         dp_n168, dp_n167, dp_n166, dp_n165, dp_n164, dp_n163, dp_n162,
         dp_n161, dp_n160, dp_n159, dp_n158, dp_n157, dp_n156, dp_n155,
         dp_n154, dp_n153, dp_n152, dp_n151, dp_n150, dp_n149, dp_n148,
         dp_n147, dp_n146, dp_n145, dp_n144, dp_n143, dp_n142, dp_n141,
         dp_n140, dp_n139, dp_n138, dp_n137, dp_n136, dp_n135, dp_n134,
         dp_n133, dp_n130, dp_n129, dp_n128, dp_n127, dp_n126, dp_n125,
         dp_n124, dp_n123, dp_n122, dp_n121, dp_n120, dp_n119, dp_n118,
         dp_n117, dp_n116, dp_n115, dp_n114, dp_n113, dp_n112, dp_n111,
         dp_n110, dp_n109, dp_n108, dp_n107, dp_n106, dp_n105, dp_n104,
         dp_n103, dp_n102, dp_n101, dp_n100, dp_n99, dp_n98, dp_n97, dp_n96,
         dp_n95, dp_n94, dp_n93, dp_n92, dp_n91, dp_n90, dp_n89, dp_n88,
         dp_n87, dp_n86, dp_n85, dp_n84, dp_n83, dp_n82, dp_n81, dp_n80,
         dp_n79, dp_n78, dp_n77, dp_n76, dp_n75, dp_n74, dp_n73, dp_n72,
         dp_n71, dp_n70, dp_n67, dp_n66, dp_n65, dp_n64, dp_n63, dp_n62,
         dp_n61, dp_n60, dp_n59, dp_n58, dp_n57, dp_n56, dp_n55, dp_n54,
         dp_n53, dp_n52, dp_n51, dp_n50, dp_n49, dp_n48, dp_n47, dp_n46,
         dp_n45, dp_n44, dp_n43, dp_n42, dp_n41, dp_n40, dp_n39, dp_n38,
         dp_n37, dp_n36, dp_n35, dp_n34, dp_n33, dp_n32, dp_n31, dp_n30,
         dp_n29, dp_n28, dp_n27, dp_n26, dp_n25, dp_n24, dp_n23, dp_n22,
         dp_n21, dp_n20, dp_n19, dp_n18, dp_n17, dp_n16, dp_n15, dp_n14,
         dp_n13, dp_n12, dp_n11, dp_n10, dp_n9, dp_n8, dp_n7, dp_n6, dp_n5,
         dp_n4, dp_n3, dp_n1015, dp_n1014, dp_n1013, dp_n1012, dp_n1011,
         dp_n1010, dp_n1009, dp_n1008, dp_n1007, dp_n1006, dp_n1005, dp_n1004,
         dp_n1003, dp_n1002, dp_n1001, dp_n1000, dp_n999, dp_n998, dp_n997,
         dp_n996, dp_n995, dp_n994, dp_n993, dp_n992, dp_n991, dp_n990,
         dp_n989, dp_n988, dp_n987, dp_n986, dp_n985, dp_n984, dp_n983,
         dp_n982, dp_n981, dp_n980, dp_n979, dp_n978, dp_n977, dp_n976,
         dp_n975, dp_n974, dp_n973, dp_n972, dp_n971, dp_n970, dp_n969,
         dp_n968, dp_n967, dp_n966, dp_n965, dp_n964, dp_n963, dp_n962,
         dp_n961, dp_n960, dp_n959, dp_n958, dp_n957, dp_n956, dp_n955,
         dp_n954, dp_n953, dp_n952, dp_n951, dp_n950, dp_n949, dp_n948,
         dp_n947, dp_n946, dp_n945, dp_n944, dp_n943, dp_n942, dp_n941,
         dp_n940, dp_n939, dp_n938, dp_n937, dp_n936, dp_n935, dp_n934,
         dp_n933, dp_n932, dp_n931, dp_n930, dp_n929, dp_n928, dp_n927,
         dp_n926, dp_n925, dp_n924, dp_n923, dp_n922, dp_n921, dp_n920,
         dp_n919, dp_n918, dp_n917, dp_n916, dp_n915, dp_n914, dp_n913,
         dp_n912, dp_n911, dp_n910, dp_n909, dp_n908, dp_n907, dp_n906,
         dp_n905, dp_n904, dp_n903, dp_n902, dp_n901, dp_n900, dp_n899,
         dp_n898, dp_n897, dp_n896, dp_n895, dp_n894, dp_n893, dp_n892,
         dp_n891, dp_n890, dp_n889, dp_n888, dp_n887, dp_n886, dp_n885,
         dp_n884, dp_n883, dp_n882, dp_n881, dp_n880, dp_n879, dp_n878,
         dp_n877, dp_n876, dp_n875, dp_n874, dp_n873, dp_n872, dp_n871,
         dp_n870, dp_n869, dp_n868, dp_n867, dp_n866, dp_n865, dp_n864,
         dp_n863, dp_n862, dp_n861, dp_n860, dp_n859, dp_n858, dp_n857,
         dp_n856, dp_n855, dp_n854, dp_n853, dp_n852, dp_n851, dp_n850,
         dp_n849, dp_n848, dp_n847, dp_n846, dp_n845, dp_n844, dp_n843,
         dp_n842, dp_n841, dp_n840, dp_n839, dp_n838, dp_n837, dp_n836,
         dp_n835, dp_n834, dp_n833, dp_n832, dp_n831, dp_n830, dp_n829,
         dp_n828, dp_n827, dp_n826, dp_n825, dp_n824, dp_n823, dp_n822,
         dp_n821, dp_n820, dp_n819, dp_n818, dp_n817, dp_n816, dp_n815,
         dp_n814, dp_n813, dp_n812, dp_n811, dp_n810, dp_n809, dp_n808,
         dp_n807, dp_n806, dp_n805, dp_n804, dp_n803, dp_n802, dp_n801,
         dp_n800, dp_n799, dp_n798, dp_n797, dp_n796, dp_n795, dp_n794,
         dp_n793, dp_n792, dp_n791, dp_n790, dp_n789, dp_n788, dp_n787,
         dp_n786, dp_n785, dp_n784, dp_n783, dp_n782, dp_n781, dp_n780,
         dp_n779, dp_n778, dp_n777, dp_n776, dp_n775, dp_n774, dp_n773,
         dp_n772, dp_n771, dp_n770, dp_n769, dp_n768, dp_n767, dp_n766,
         dp_n765, dp_n764, dp_n763, dp_n762, dp_n761, dp_n760, dp_n759,
         dp_n758, dp_n757, dp_n756, dp_n755, dp_n754, dp_n753, dp_n752,
         dp_n751, dp_n750, dp_n749, dp_n748, dp_n747, dp_n746, dp_n745,
         dp_n744, dp_n743, dp_n742, dp_n741, dp_n740, dp_n739, dp_n738,
         dp_n737, dp_n736, dp_n735, dp_n734, dp_n733, dp_n732, dp_n731,
         dp_n730, dp_n729, dp_n728, dp_n727, dp_n726, dp_n725, dp_n724,
         dp_n723, dp_n722, dp_n721, dp_n720, dp_n719, dp_n718, dp_n717,
         dp_n716, dp_n715, dp_n714, dp_n713, dp_n712, dp_n706, dp_n705,
         dp_n704, dp_n703, dp_n702, dp_n701, dp_n700, dp_n699, dp_n698,
         dp_n697, dp_n696, dp_n695, dp_n694, dp_n693, dp_n692, dp_n691,
         dp_n690, dp_n689, dp_n688, dp_n687, dp_n686, dp_n685, dp_n684,
         dp_n683, dp_n682, dp_n681, dp_n680, dp_n679, dp_n678, dp_n677,
         dp_n676, dp_n675, dp_n674, dp_n673, dp_n672, dp_n671, dp_n670,
         dp_n669, dp_n668, dp_n667, dp_n666, dp_n665, dp_n664, dp_n663,
         dp_n662, dp_n661, dp_n660, dp_n659, dp_n658, dp_n657, dp_n656,
         dp_n655, dp_n654, dp_n653, dp_n652, dp_n651, dp_n650, dp_n649,
         dp_n583, dp_n582, dp_n581, dp_n580, dp_n579, dp_n578, dp_n577,
         dp_n576, dp_n575, dp_n574, dp_n573, dp_n572, dp_n571, dp_n570,
         dp_n569, dp_n568, dp_n567, dp_n566, dp_n565, dp_n564, dp_n563,
         dp_n562, dp_n561, dp_n560, dp_n559, dp_n558, dp_n557, dp_n556,
         dp_n555, dp_n554, dp_n553, dp_n552, dp_n551, dp_n550, dp_n549,
         dp_n548, dp_n547, dp_n546, dp_n545, dp_n544, dp_n543, dp_n542,
         dp_n541, dp_n540, dp_n539, dp_n538, dp_n537, dp_n536, dp_n535,
         dp_n534, dp_n533, dp_n532, dp_n531, dp_n530, dp_n529, dp_n528,
         dp_n527, dp_n526, dp_n524, dp_n522, dp_n520, dp_n518, dp_n516,
         dp_n515, dp_n514, dp_n513, dp_n512, dp_n511, dp_n510, dp_n509,
         dp_n508, dp_n507, dp_n506, dp_n505, dp_n504, dp_n503, dp_n502,
         dp_n501, dp_n500, dp_n499, dp_n498, dp_n497, dp_n496, dp_n495,
         dp_n494, dp_n493, dp_n492, dp_n491, dp_n490, dp_n489, dp_n488,
         dp_n487, dp_n486, dp_n485, dp_n484, dp_n483, dp_n482, dp_n481,
         dp_n480, dp_n479, dp_n478, dp_n477, dp_n476, dp_n475, dp_n474,
         dp_n473, dp_n472, dp_n471, dp_n470, dp_n469, dp_n468, dp_n467,
         dp_n466, dp_n465, dp_n464, dp_n463, dp_n462, dp_n461, dp_n460,
         dp_n459, dp_n458, dp_n457, dp_n456, dp_n455, dp_n454, dp_n453,
         dp_n452, dp_n451, dp_n450, dp_n449, dp_n448, dp_n447, dp_n446,
         dp_n445, dp_n444, dp_n443, dp_n442, dp_n441, dp_n440, dp_n439,
         dp_n438, dp_n437, dp_n436, dp_n435, dp_n434, dp_n433, dp_n432,
         dp_n431, dp_n430, dp_n429, dp_n428, dp_n427, dp_n426, dp_n425,
         dp_n424, dp_n423, dp_n422, dp_n421, dp_n420, dp_n419, dp_n418,
         dp_n417, dp_n416, dp_n415, dp_n414, dp_n401, dp_n400, dp_n399,
         dp_n398, dp_n397, dp_n396, dp_n395, dp_n394, dp_n393, dp_n392,
         dp_n391, dp_n390, dp_n389, dp_n388, dp_n387, dp_n386, dp_n385,
         dp_n384, dp_n383, dp_n382, dp_n381, dp_n380, dp_n379, dp_n378,
         dp_n377, dp_n376, dp_n375, dp_n374, dp_n373, dp_n372, dp_n371,
         dp_n370, dp_n369, dp_n368, dp_n367, dp_n366, dp_n365, dp_n364,
         dp_n363, dp_n362, dp_n361, dp_n360, dp_n359, dp_n358, dp_n357,
         dp_n356, dp_n355, dp_n354, dp_n353, dp_n352, dp_n351, dp_n350,
         dp_n349, dp_n348, dp_n347, dp_n346, dp_n345, dp_n344, dp_n343,
         dp_n342, dp_n341, dp_n340, dp_n339, dp_n338, dp_n337, dp_n336,
         dp_n335, dp_n302, dp_n301, dp_n132, dp_n131, dp_n69, dp_n68,
         dp_branch_t_ex_o, dp_ir_0_, dp_ir_1_, dp_ir_2_, dp_ir_3_, dp_ir_4_,
         dp_ir_5_, dp_ir_6_, dp_ir_7_, dp_ir_8_, dp_ir_9_, dp_ir_10_,
         dp_ir_11_, dp_ir_12_, dp_ir_13_, dp_ir_14_, dp_ir_15_, dp_ir_16_,
         dp_ir_17_, dp_ir_18_, dp_ir_19_, dp_ir_20_, dp_ir_21_, dp_ir_22_,
         dp_ir_23_, dp_ir_24_, dp_ir_25_, dp_if_stage_n41, dp_if_stage_n40,
         dp_if_stage_n39, dp_if_stage_n38, dp_if_stage_n37, dp_if_stage_n36,
         dp_if_stage_n35, dp_if_stage_n34, dp_if_stage_n33, dp_if_stage_n16,
         dp_if_stage_n15, dp_if_stage_n14, dp_if_stage_n13, dp_if_stage_n12,
         dp_if_stage_n11, dp_if_stage_n10, dp_if_stage_n9, dp_if_stage_n8,
         dp_if_stage_n7, dp_if_stage_n6, dp_if_stage_n5, dp_if_stage_n4,
         dp_if_stage_n3, dp_if_stage_n2, dp_if_stage_n1, dp_if_stage_n97,
         dp_if_stage_n95, dp_if_stage_n94, dp_if_stage_n93, dp_if_stage_n92,
         dp_if_stage_n91, dp_if_stage_n90, dp_if_stage_n89, dp_if_stage_n88,
         dp_if_stage_n87, dp_if_stage_n86, dp_if_stage_n85, dp_if_stage_n84,
         dp_if_stage_n83, dp_if_stage_n82, dp_if_stage_n81, dp_if_stage_n64,
         dp_if_stage_n63, dp_if_stage_n62, dp_if_stage_n61, dp_if_stage_n60,
         dp_if_stage_n59, dp_if_stage_n58, dp_if_stage_n57, dp_if_stage_n56,
         dp_if_stage_n55, dp_if_stage_n54, dp_if_stage_n53, dp_if_stage_n52,
         dp_if_stage_n51, dp_if_stage_n50, dp_if_stage_n49, dp_if_stage_n32,
         dp_if_stage_n31, dp_if_stage_n30, dp_if_stage_n29, dp_if_stage_n28,
         dp_if_stage_n27, dp_if_stage_n26, dp_if_stage_n25, dp_if_stage_n24,
         dp_if_stage_n23, dp_if_stage_n22, dp_if_stage_n21, dp_if_stage_n20,
         dp_if_stage_n19, dp_if_stage_n18, dp_if_stage_n17,
         dp_if_stage_NPC_4_i_2_, dp_if_stage_NPC_4_i_3_,
         dp_if_stage_NPC_4_i_4_, dp_if_stage_NPC_4_i_5_,
         dp_if_stage_NPC_4_i_6_, dp_if_stage_NPC_4_i_7_,
         dp_if_stage_NPC_4_i_8_, dp_if_stage_NPC_4_i_9_,
         dp_if_stage_NPC_4_i_10_, dp_if_stage_NPC_4_i_11_,
         dp_if_stage_NPC_4_i_12_, dp_if_stage_NPC_4_i_13_,
         dp_if_stage_NPC_4_i_14_, dp_if_stage_NPC_4_i_15_,
         dp_if_stage_NPC_4_i_16_, dp_if_stage_NPC_4_i_17_,
         dp_if_stage_NPC_4_i_18_, dp_if_stage_NPC_4_i_19_,
         dp_if_stage_NPC_4_i_20_, dp_if_stage_NPC_4_i_21_,
         dp_if_stage_NPC_4_i_22_, dp_if_stage_NPC_4_i_23_,
         dp_if_stage_NPC_4_i_24_, dp_if_stage_NPC_4_i_25_,
         dp_if_stage_NPC_4_i_26_, dp_if_stage_NPC_4_i_27_,
         dp_if_stage_NPC_4_i_28_, dp_if_stage_NPC_4_i_29_,
         dp_if_stage_NPC_4_i_30_, dp_if_stage_NPC_4_i_31_, dp_if_stage_mux_n7,
         dp_if_stage_mux_n6, dp_if_stage_mux_n5, dp_if_stage_mux_n4,
         dp_if_stage_mux_n3, dp_if_stage_mux_n2, dp_if_stage_mux_n1,
         dp_if_stage_mux_n65, dp_if_stage_mux_n64, dp_if_stage_mux_n63,
         dp_if_stage_mux_n62, dp_if_stage_mux_n61, dp_if_stage_mux_n60,
         dp_if_stage_mux_n59, dp_if_stage_mux_n54, dp_if_stage_mux_n43,
         dp_if_stage_mux_n40, dp_if_stage_mux_n39, dp_if_stage_mux_n38,
         dp_if_stage_mux_n37, dp_if_stage_mux_n36, dp_if_stage_mux_n35,
         dp_if_stage_mux_n34, dp_if_stage_add_77_n61, dp_if_stage_add_77_n60,
         dp_if_stage_add_77_n59, dp_if_stage_add_77_n58,
         dp_if_stage_add_77_n57, dp_if_stage_add_77_n56,
         dp_if_stage_add_77_n55, dp_if_stage_add_77_n54,
         dp_if_stage_add_77_n53, dp_if_stage_add_77_n52,
         dp_if_stage_add_77_n51, dp_if_stage_add_77_n50,
         dp_if_stage_add_77_n49, dp_if_stage_add_77_n48,
         dp_if_stage_add_77_n47, dp_if_stage_add_77_n46,
         dp_if_stage_add_77_n45, dp_if_stage_add_77_n44,
         dp_if_stage_add_77_n43, dp_if_stage_add_77_n42,
         dp_if_stage_add_77_n41, dp_if_stage_add_77_n40,
         dp_if_stage_add_77_n39, dp_if_stage_add_77_n38,
         dp_if_stage_add_77_n37, dp_if_stage_add_77_n36,
         dp_if_stage_add_77_n35, dp_if_stage_add_77_n34,
         dp_if_stage_add_77_n33, dp_if_stage_add_77_n32,
         dp_if_stage_add_77_n31, dp_if_stage_add_77_n30,
         dp_if_stage_add_77_n29, dp_if_stage_add_77_n28,
         dp_if_stage_add_77_n27, dp_if_stage_add_77_n26,
         dp_if_stage_add_77_n25, dp_if_stage_add_77_n24,
         dp_if_stage_add_77_n23, dp_if_stage_add_77_n22,
         dp_if_stage_add_77_n21, dp_if_stage_add_77_n20,
         dp_if_stage_add_77_n19, dp_if_stage_add_77_n18,
         dp_if_stage_add_77_n16, dp_if_stage_add_77_n15,
         dp_if_stage_add_77_n14, dp_if_stage_add_77_n13,
         dp_if_stage_add_77_n12, dp_if_stage_add_77_n11,
         dp_if_stage_add_77_n10, dp_if_stage_add_77_n9, dp_if_stage_add_77_n8,
         dp_if_stage_add_77_n7, dp_if_stage_add_77_n6, dp_if_stage_add_77_n5,
         dp_if_stage_add_77_n4, dp_if_stage_add_77_n3, dp_if_stage_add_77_n2,
         dp_if_stage_add_77_n1, dp_id_stage_n40, dp_id_stage_n39,
         dp_id_stage_n38, dp_id_stage_n37, dp_id_stage_n36, dp_id_stage_n35,
         dp_id_stage_n34, dp_id_stage_n33, dp_id_stage_n32, dp_id_stage_n31,
         dp_id_stage_n30, dp_id_stage_n29, dp_id_stage_n28, dp_id_stage_n27,
         dp_id_stage_n26, dp_id_stage_n25, dp_id_stage_n24, dp_id_stage_n16,
         dp_id_stage_n15, dp_id_stage_n14, dp_id_stage_n13, dp_id_stage_n12,
         dp_id_stage_n11, dp_id_stage_n10, dp_id_stage_n9, dp_id_stage_n8,
         dp_id_stage_n7, dp_id_stage_n6, dp_id_stage_n5, dp_id_stage_n4,
         dp_id_stage_n3, dp_id_stage_n2, dp_id_stage_n1, dp_id_stage_n23,
         dp_id_stage_n22, dp_id_stage_n21, dp_id_stage_n20, dp_id_stage_n19,
         dp_id_stage_n18, dp_id_stage_n17, dp_id_stage_regfile_cpu_work,
         dp_id_stage_regfile_sel_wp, dp_id_stage_regfile_end_sf,
         dp_id_stage_regfile_canrestore, dp_id_stage_regfile_cansave,
         dp_id_stage_regfile_up_dwn_rest, dp_id_stage_regfile_up_dwn_save,
         dp_id_stage_regfile_up_dwn_cwp, dp_id_stage_regfile_up_dwn_swp,
         dp_id_stage_regfile_rst_spill_fill, dp_id_stage_regfile_rst_swp,
         dp_id_stage_regfile_cnt_save, dp_id_stage_regfile_cnt_cwp,
         dp_id_stage_regfile_cnt_swp, dp_id_stage_regfile_rst_rf,
         dp_id_stage_regfile_rf_enable, dp_id_stage_regfile_wr_cu,
         dp_id_stage_regfile_rd_cu, dp_id_stage_regfile_ControlUnit_n41,
         dp_id_stage_regfile_ControlUnit_n15,
         dp_id_stage_regfile_ControlUnit_n10,
         dp_id_stage_regfile_ControlUnit_n9,
         dp_id_stage_regfile_ControlUnit_n6,
         dp_id_stage_regfile_ControlUnit_n5,
         dp_id_stage_regfile_ControlUnit_n4,
         dp_id_stage_regfile_ControlUnit_n3,
         dp_id_stage_regfile_ControlUnit_n1,
         dp_id_stage_regfile_ControlUnit_n40,
         dp_id_stage_regfile_ControlUnit_n39,
         dp_id_stage_regfile_ControlUnit_n38,
         dp_id_stage_regfile_ControlUnit_n37,
         dp_id_stage_regfile_ControlUnit_n36,
         dp_id_stage_regfile_ControlUnit_n35,
         dp_id_stage_regfile_ControlUnit_n34,
         dp_id_stage_regfile_ControlUnit_n33,
         dp_id_stage_regfile_ControlUnit_n32,
         dp_id_stage_regfile_ControlUnit_n31,
         dp_id_stage_regfile_ControlUnit_n30,
         dp_id_stage_regfile_ControlUnit_n29,
         dp_id_stage_regfile_ControlUnit_n28,
         dp_id_stage_regfile_ControlUnit_n27,
         dp_id_stage_regfile_ControlUnit_n26,
         dp_id_stage_regfile_ControlUnit_n25,
         dp_id_stage_regfile_ControlUnit_n24,
         dp_id_stage_regfile_ControlUnit_n23,
         dp_id_stage_regfile_ControlUnit_n22,
         dp_id_stage_regfile_ControlUnit_n21,
         dp_id_stage_regfile_ControlUnit_n20,
         dp_id_stage_regfile_ControlUnit_n19,
         dp_id_stage_regfile_ControlUnit_n18,
         dp_id_stage_regfile_ControlUnit_n17,
         dp_id_stage_regfile_ControlUnit_n16,
         dp_id_stage_regfile_ControlUnit_n14,
         dp_id_stage_regfile_ControlUnit_n13,
         dp_id_stage_regfile_ControlUnit_n12,
         dp_id_stage_regfile_ControlUnit_current_state_0_,
         dp_id_stage_regfile_ControlUnit_current_state_2_,
         dp_id_stage_regfile_ControlUnit_current_state_3_,
         dp_id_stage_regfile_DataPath_mux_en_control_out,
         dp_id_stage_regfile_DataPath_mux_wr_control_out,
         dp_id_stage_regfile_DataPath_mux_rd2_control_out,
         dp_id_stage_regfile_DataPath_mux_rd1_control_out,
         dp_id_stage_regfile_DataPath_cwp_1_0_,
         dp_id_stage_regfile_DataPath_spill_fill_addr_0_,
         dp_id_stage_regfile_DataPath_spill_fill_addr_1_,
         dp_id_stage_regfile_DataPath_spill_fill_addr_2_,
         dp_id_stage_regfile_DataPath_spill_fill_addr_3_,
         dp_id_stage_regfile_DataPath_spill_fill_addr_4_,
         dp_id_stage_regfile_DataPath_spill_fill_addr_5_,
         dp_id_stage_regfile_DataPath_sf_wp_0_,
         dp_id_stage_regfile_DataPath_addr_sf_in_0_,
         dp_id_stage_regfile_DataPath_addr_sf_in_1_,
         dp_id_stage_regfile_DataPath_addr_sf_in_2_,
         dp_id_stage_regfile_DataPath_CWP_0_,
         dp_id_stage_regfile_DataPath_Conv_RD1_n8,
         dp_id_stage_regfile_DataPath_Conv_RD1_n4,
         dp_id_stage_regfile_DataPath_Conv_RD1_n3,
         dp_id_stage_regfile_DataPath_Conv_RD1_n2,
         dp_id_stage_regfile_DataPath_Conv_RD1_n1,
         dp_id_stage_regfile_DataPath_Conv_RD1_n22,
         dp_id_stage_regfile_DataPath_Conv_RD1_n21,
         dp_id_stage_regfile_DataPath_Conv_RD1_n20,
         dp_id_stage_regfile_DataPath_Conv_RD1_n19,
         dp_id_stage_regfile_DataPath_Conv_RD1_n18,
         dp_id_stage_regfile_DataPath_Conv_RD1_N5,
         dp_id_stage_regfile_DataPath_Conv_RD1_N1,
         dp_id_stage_regfile_DataPath_Conv_RD2_n13,
         dp_id_stage_regfile_DataPath_Conv_RD2_n12,
         dp_id_stage_regfile_DataPath_Conv_RD2_n11,
         dp_id_stage_regfile_DataPath_Conv_RD2_n10,
         dp_id_stage_regfile_DataPath_Conv_RD2_n9,
         dp_id_stage_regfile_DataPath_Conv_RD2_n8,
         dp_id_stage_regfile_DataPath_Conv_RD2_n4,
         dp_id_stage_regfile_DataPath_Conv_RD2_n3,
         dp_id_stage_regfile_DataPath_Conv_RD2_n2,
         dp_id_stage_regfile_DataPath_Conv_RD2_n1,
         dp_id_stage_regfile_DataPath_Conv_RD2_N5,
         dp_id_stage_regfile_DataPath_Conv_RD2_N1,
         dp_id_stage_regfile_DataPath_Conv_W_n13,
         dp_id_stage_regfile_DataPath_Conv_W_n12,
         dp_id_stage_regfile_DataPath_Conv_W_n11,
         dp_id_stage_regfile_DataPath_Conv_W_n10,
         dp_id_stage_regfile_DataPath_Conv_W_n9,
         dp_id_stage_regfile_DataPath_Conv_W_n8,
         dp_id_stage_regfile_DataPath_Conv_W_n4,
         dp_id_stage_regfile_DataPath_Conv_W_n3,
         dp_id_stage_regfile_DataPath_Conv_W_n2,
         dp_id_stage_regfile_DataPath_Conv_W_n1,
         dp_id_stage_regfile_DataPath_Conv_W_N5,
         dp_id_stage_regfile_DataPath_Conv_W_N1,
         dp_id_stage_regfile_DataPath_SF_converter_n10,
         dp_id_stage_regfile_DataPath_SF_converter_n9,
         dp_id_stage_regfile_DataPath_SF_converter_n8,
         dp_id_stage_regfile_DataPath_SF_converter_n7,
         dp_id_stage_regfile_DataPath_SF_converter_n6,
         dp_id_stage_regfile_DataPath_SF_converter_n5,
         dp_id_stage_regfile_DataPath_SF_converter_n4,
         dp_id_stage_regfile_DataPath_SF_converter_n3,
         dp_id_stage_regfile_DataPath_SF_converter_n2,
         dp_id_stage_regfile_DataPath_SF_converter_n1,
         dp_id_stage_regfile_DataPath_SF_converter_N5,
         dp_id_stage_regfile_DataPath_SF_converter_N1,
         dp_id_stage_regfile_DataPath_Cwp_counter_n4,
         dp_id_stage_regfile_DataPath_Cwp_counter_n2,
         dp_id_stage_regfile_DataPath_Cwp_counter_n5,
         dp_id_stage_regfile_DataPath_Cwp_counter_n3,
         dp_id_stage_regfile_DataPath_Cwp_counter_n1,
         dp_id_stage_regfile_DataPath_Swp_counter_n8,
         dp_id_stage_regfile_DataPath_Swp_counter_n7,
         dp_id_stage_regfile_DataPath_Swp_counter_n6,
         dp_id_stage_regfile_DataPath_Swp_counter_n4,
         dp_id_stage_regfile_DataPath_Swp_counter_n2,
         dp_id_stage_regfile_DataPath_Swp_counter_Q_0_,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n16,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n12,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n4,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n3,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n2,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n1,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n21,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n20,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n19,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n18,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n17,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n15,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n14,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n13,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n11,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n10,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n9,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n8,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n7,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n6,
         dp_id_stage_regfile_DataPath_Spill_fill_counter_n5,
         dp_id_stage_regfile_DataPath_CANSAVE_counter_n8,
         dp_id_stage_regfile_DataPath_CANSAVE_counter_n7,
         dp_id_stage_regfile_DataPath_CANSAVE_counter_n6,
         dp_id_stage_regfile_DataPath_CANSAVE_counter_n4,
         dp_id_stage_regfile_DataPath_CANSAVE_counter_n2,
         dp_id_stage_regfile_DataPath_CANRESTORE_counter_n8,
         dp_id_stage_regfile_DataPath_CANRESTORE_counter_n7,
         dp_id_stage_regfile_DataPath_CANRESTORE_counter_n6,
         dp_id_stage_regfile_DataPath_CANRESTORE_counter_n4,
         dp_id_stage_regfile_DataPath_CANRESTORE_counter_n2,
         dp_id_stage_regfile_DataPath_Mux_rd_n1,
         dp_id_stage_regfile_DataPath_Mux_rd_n13,
         dp_id_stage_regfile_DataPath_Mux_rd_n12,
         dp_id_stage_regfile_DataPath_Mux_rd_n11,
         dp_id_stage_regfile_DataPath_Mux_rd_n10,
         dp_id_stage_regfile_DataPath_Mux_rd_n9,
         dp_id_stage_regfile_DataPath_Mux_rd_n8,
         dp_id_stage_regfile_DataPath_Mux_wr_n7,
         dp_id_stage_regfile_DataPath_Mux_wr_n6,
         dp_id_stage_regfile_DataPath_Mux_wr_n5,
         dp_id_stage_regfile_DataPath_Mux_wr_n4,
         dp_id_stage_regfile_DataPath_Mux_wr_n3,
         dp_id_stage_regfile_DataPath_Mux_wr_n2,
         dp_id_stage_regfile_DataPath_Mux_wr_n1,
         dp_id_stage_regfile_DataPath_Mux_sf_n1,
         dp_id_stage_regfile_DataPath_Mux_sf_n3,
         dp_id_stage_regfile_DataPath_Mux_rd1_control_n2,
         dp_id_stage_regfile_DataPath_Mux_rd1_control_n3,
         dp_id_stage_regfile_DataPath_Mux_rd2_control_n4,
         dp_id_stage_regfile_DataPath_Mux_rd2_control_n2,
         dp_id_stage_regfile_DataPath_Mux_wr_control_n4,
         dp_id_stage_regfile_DataPath_Mux_wr_control_n2,
         dp_id_stage_regfile_DataPath_Mux_en_control_n4,
         dp_id_stage_regfile_DataPath_Mux_en_control_n2,
         dp_id_stage_regfile_DataPath_Physical_RF_n4270,
         dp_id_stage_regfile_DataPath_Physical_RF_n4269,
         dp_id_stage_regfile_DataPath_Physical_RF_n4268,
         dp_id_stage_regfile_DataPath_Physical_RF_n4267,
         dp_id_stage_regfile_DataPath_Physical_RF_n4266,
         dp_id_stage_regfile_DataPath_Physical_RF_n4265,
         dp_id_stage_regfile_DataPath_Physical_RF_n4264,
         dp_id_stage_regfile_DataPath_Physical_RF_n4263,
         dp_id_stage_regfile_DataPath_Physical_RF_n4262,
         dp_id_stage_regfile_DataPath_Physical_RF_n4261,
         dp_id_stage_regfile_DataPath_Physical_RF_n4260,
         dp_id_stage_regfile_DataPath_Physical_RF_n4259,
         dp_id_stage_regfile_DataPath_Physical_RF_n4258,
         dp_id_stage_regfile_DataPath_Physical_RF_n4257,
         dp_id_stage_regfile_DataPath_Physical_RF_n4256,
         dp_id_stage_regfile_DataPath_Physical_RF_n4255,
         dp_id_stage_regfile_DataPath_Physical_RF_n4254,
         dp_id_stage_regfile_DataPath_Physical_RF_n4253,
         dp_id_stage_regfile_DataPath_Physical_RF_n4252,
         dp_id_stage_regfile_DataPath_Physical_RF_n4251,
         dp_id_stage_regfile_DataPath_Physical_RF_n4250,
         dp_id_stage_regfile_DataPath_Physical_RF_n4249,
         dp_id_stage_regfile_DataPath_Physical_RF_n4248,
         dp_id_stage_regfile_DataPath_Physical_RF_n4247,
         dp_id_stage_regfile_DataPath_Physical_RF_n4246,
         dp_id_stage_regfile_DataPath_Physical_RF_n4245,
         dp_id_stage_regfile_DataPath_Physical_RF_n4244,
         dp_id_stage_regfile_DataPath_Physical_RF_n4243,
         dp_id_stage_regfile_DataPath_Physical_RF_n4242,
         dp_id_stage_regfile_DataPath_Physical_RF_n4241,
         dp_id_stage_regfile_DataPath_Physical_RF_n4240,
         dp_id_stage_regfile_DataPath_Physical_RF_n4239,
         dp_id_stage_regfile_DataPath_Physical_RF_n4238,
         dp_id_stage_regfile_DataPath_Physical_RF_n4237,
         dp_id_stage_regfile_DataPath_Physical_RF_n4236,
         dp_id_stage_regfile_DataPath_Physical_RF_n4235,
         dp_id_stage_regfile_DataPath_Physical_RF_n4234,
         dp_id_stage_regfile_DataPath_Physical_RF_n4233,
         dp_id_stage_regfile_DataPath_Physical_RF_n4232,
         dp_id_stage_regfile_DataPath_Physical_RF_n4231,
         dp_id_stage_regfile_DataPath_Physical_RF_n4230,
         dp_id_stage_regfile_DataPath_Physical_RF_n4229,
         dp_id_stage_regfile_DataPath_Physical_RF_n4228,
         dp_id_stage_regfile_DataPath_Physical_RF_n4227,
         dp_id_stage_regfile_DataPath_Physical_RF_n4226,
         dp_id_stage_regfile_DataPath_Physical_RF_n4225,
         dp_id_stage_regfile_DataPath_Physical_RF_n4224,
         dp_id_stage_regfile_DataPath_Physical_RF_n4223,
         dp_id_stage_regfile_DataPath_Physical_RF_n4222,
         dp_id_stage_regfile_DataPath_Physical_RF_n4221,
         dp_id_stage_regfile_DataPath_Physical_RF_n4220,
         dp_id_stage_regfile_DataPath_Physical_RF_n4219,
         dp_id_stage_regfile_DataPath_Physical_RF_n4218,
         dp_id_stage_regfile_DataPath_Physical_RF_n4217,
         dp_id_stage_regfile_DataPath_Physical_RF_n4216,
         dp_id_stage_regfile_DataPath_Physical_RF_n4215,
         dp_id_stage_regfile_DataPath_Physical_RF_n4214,
         dp_id_stage_regfile_DataPath_Physical_RF_n4213,
         dp_id_stage_regfile_DataPath_Physical_RF_n4212,
         dp_id_stage_regfile_DataPath_Physical_RF_n4211,
         dp_id_stage_regfile_DataPath_Physical_RF_n4210,
         dp_id_stage_regfile_DataPath_Physical_RF_n4209,
         dp_id_stage_regfile_DataPath_Physical_RF_n4208,
         dp_id_stage_regfile_DataPath_Physical_RF_n4207,
         dp_id_stage_regfile_DataPath_Physical_RF_n4206,
         dp_id_stage_regfile_DataPath_Physical_RF_n4205,
         dp_id_stage_regfile_DataPath_Physical_RF_n4204,
         dp_id_stage_regfile_DataPath_Physical_RF_n4203,
         dp_id_stage_regfile_DataPath_Physical_RF_n4202,
         dp_id_stage_regfile_DataPath_Physical_RF_n4201,
         dp_id_stage_regfile_DataPath_Physical_RF_n4200,
         dp_id_stage_regfile_DataPath_Physical_RF_n4199,
         dp_id_stage_regfile_DataPath_Physical_RF_n4198,
         dp_id_stage_regfile_DataPath_Physical_RF_n4197,
         dp_id_stage_regfile_DataPath_Physical_RF_n4196,
         dp_id_stage_regfile_DataPath_Physical_RF_n4195,
         dp_id_stage_regfile_DataPath_Physical_RF_n4194,
         dp_id_stage_regfile_DataPath_Physical_RF_n4193,
         dp_id_stage_regfile_DataPath_Physical_RF_n4192,
         dp_id_stage_regfile_DataPath_Physical_RF_n4191,
         dp_id_stage_regfile_DataPath_Physical_RF_n4190,
         dp_id_stage_regfile_DataPath_Physical_RF_n4189,
         dp_id_stage_regfile_DataPath_Physical_RF_n4188,
         dp_id_stage_regfile_DataPath_Physical_RF_n4187,
         dp_id_stage_regfile_DataPath_Physical_RF_n4186,
         dp_id_stage_regfile_DataPath_Physical_RF_n4185,
         dp_id_stage_regfile_DataPath_Physical_RF_n4184,
         dp_id_stage_regfile_DataPath_Physical_RF_n4183,
         dp_id_stage_regfile_DataPath_Physical_RF_n4182,
         dp_id_stage_regfile_DataPath_Physical_RF_n4181,
         dp_id_stage_regfile_DataPath_Physical_RF_n4180,
         dp_id_stage_regfile_DataPath_Physical_RF_n4179,
         dp_id_stage_regfile_DataPath_Physical_RF_n4178,
         dp_id_stage_regfile_DataPath_Physical_RF_n4177,
         dp_id_stage_regfile_DataPath_Physical_RF_n4176,
         dp_id_stage_regfile_DataPath_Physical_RF_n4175,
         dp_id_stage_regfile_DataPath_Physical_RF_n4174,
         dp_id_stage_regfile_DataPath_Physical_RF_n4173,
         dp_id_stage_regfile_DataPath_Physical_RF_n4172,
         dp_id_stage_regfile_DataPath_Physical_RF_n4171,
         dp_id_stage_regfile_DataPath_Physical_RF_n4170,
         dp_id_stage_regfile_DataPath_Physical_RF_n4169,
         dp_id_stage_regfile_DataPath_Physical_RF_n4168,
         dp_id_stage_regfile_DataPath_Physical_RF_n4167,
         dp_id_stage_regfile_DataPath_Physical_RF_n4166,
         dp_id_stage_regfile_DataPath_Physical_RF_n4165,
         dp_id_stage_regfile_DataPath_Physical_RF_n4164,
         dp_id_stage_regfile_DataPath_Physical_RF_n4163,
         dp_id_stage_regfile_DataPath_Physical_RF_n4162,
         dp_id_stage_regfile_DataPath_Physical_RF_n4161,
         dp_id_stage_regfile_DataPath_Physical_RF_n4160,
         dp_id_stage_regfile_DataPath_Physical_RF_n4159,
         dp_id_stage_regfile_DataPath_Physical_RF_n4158,
         dp_id_stage_regfile_DataPath_Physical_RF_n4157,
         dp_id_stage_regfile_DataPath_Physical_RF_n4156,
         dp_id_stage_regfile_DataPath_Physical_RF_n4155,
         dp_id_stage_regfile_DataPath_Physical_RF_n4154,
         dp_id_stage_regfile_DataPath_Physical_RF_n4153,
         dp_id_stage_regfile_DataPath_Physical_RF_n4152,
         dp_id_stage_regfile_DataPath_Physical_RF_n4151,
         dp_id_stage_regfile_DataPath_Physical_RF_n4150,
         dp_id_stage_regfile_DataPath_Physical_RF_n4149,
         dp_id_stage_regfile_DataPath_Physical_RF_n4148,
         dp_id_stage_regfile_DataPath_Physical_RF_n4147,
         dp_id_stage_regfile_DataPath_Physical_RF_n4146,
         dp_id_stage_regfile_DataPath_Physical_RF_n4145,
         dp_id_stage_regfile_DataPath_Physical_RF_n4144,
         dp_id_stage_regfile_DataPath_Physical_RF_n4143,
         dp_id_stage_regfile_DataPath_Physical_RF_n4142,
         dp_id_stage_regfile_DataPath_Physical_RF_n4141,
         dp_id_stage_regfile_DataPath_Physical_RF_n4140,
         dp_id_stage_regfile_DataPath_Physical_RF_n4139,
         dp_id_stage_regfile_DataPath_Physical_RF_n4138,
         dp_id_stage_regfile_DataPath_Physical_RF_n4137,
         dp_id_stage_regfile_DataPath_Physical_RF_n4136,
         dp_id_stage_regfile_DataPath_Physical_RF_n4135,
         dp_id_stage_regfile_DataPath_Physical_RF_n4134,
         dp_id_stage_regfile_DataPath_Physical_RF_n4133,
         dp_id_stage_regfile_DataPath_Physical_RF_n4132,
         dp_id_stage_regfile_DataPath_Physical_RF_n4131,
         dp_id_stage_regfile_DataPath_Physical_RF_n4130,
         dp_id_stage_regfile_DataPath_Physical_RF_n4129,
         dp_id_stage_regfile_DataPath_Physical_RF_n4128,
         dp_id_stage_regfile_DataPath_Physical_RF_n4127,
         dp_id_stage_regfile_DataPath_Physical_RF_n4126,
         dp_id_stage_regfile_DataPath_Physical_RF_n4125,
         dp_id_stage_regfile_DataPath_Physical_RF_n4124,
         dp_id_stage_regfile_DataPath_Physical_RF_n4123,
         dp_id_stage_regfile_DataPath_Physical_RF_n4122,
         dp_id_stage_regfile_DataPath_Physical_RF_n4121,
         dp_id_stage_regfile_DataPath_Physical_RF_n4120,
         dp_id_stage_regfile_DataPath_Physical_RF_n4119,
         dp_id_stage_regfile_DataPath_Physical_RF_n4118,
         dp_id_stage_regfile_DataPath_Physical_RF_n4117,
         dp_id_stage_regfile_DataPath_Physical_RF_n4116,
         dp_id_stage_regfile_DataPath_Physical_RF_n4115,
         dp_id_stage_regfile_DataPath_Physical_RF_n4114,
         dp_id_stage_regfile_DataPath_Physical_RF_n4113,
         dp_id_stage_regfile_DataPath_Physical_RF_n4112,
         dp_id_stage_regfile_DataPath_Physical_RF_n4111,
         dp_id_stage_regfile_DataPath_Physical_RF_n4110,
         dp_id_stage_regfile_DataPath_Physical_RF_n4109,
         dp_id_stage_regfile_DataPath_Physical_RF_n4108,
         dp_id_stage_regfile_DataPath_Physical_RF_n4107,
         dp_id_stage_regfile_DataPath_Physical_RF_n4106,
         dp_id_stage_regfile_DataPath_Physical_RF_n4105,
         dp_id_stage_regfile_DataPath_Physical_RF_n4104,
         dp_id_stage_regfile_DataPath_Physical_RF_n4103,
         dp_id_stage_regfile_DataPath_Physical_RF_n4102,
         dp_id_stage_regfile_DataPath_Physical_RF_n4101,
         dp_id_stage_regfile_DataPath_Physical_RF_n4100,
         dp_id_stage_regfile_DataPath_Physical_RF_n4099,
         dp_id_stage_regfile_DataPath_Physical_RF_n4098,
         dp_id_stage_regfile_DataPath_Physical_RF_n4097,
         dp_id_stage_regfile_DataPath_Physical_RF_n4096,
         dp_id_stage_regfile_DataPath_Physical_RF_n4095,
         dp_id_stage_regfile_DataPath_Physical_RF_n4094,
         dp_id_stage_regfile_DataPath_Physical_RF_n4093,
         dp_id_stage_regfile_DataPath_Physical_RF_n4092,
         dp_id_stage_regfile_DataPath_Physical_RF_n4091,
         dp_id_stage_regfile_DataPath_Physical_RF_n4090,
         dp_id_stage_regfile_DataPath_Physical_RF_n4089,
         dp_id_stage_regfile_DataPath_Physical_RF_n4088,
         dp_id_stage_regfile_DataPath_Physical_RF_n4087,
         dp_id_stage_regfile_DataPath_Physical_RF_n4086,
         dp_id_stage_regfile_DataPath_Physical_RF_n4085,
         dp_id_stage_regfile_DataPath_Physical_RF_n4084,
         dp_id_stage_regfile_DataPath_Physical_RF_n4083,
         dp_id_stage_regfile_DataPath_Physical_RF_n4082,
         dp_id_stage_regfile_DataPath_Physical_RF_n4081,
         dp_id_stage_regfile_DataPath_Physical_RF_n4080,
         dp_id_stage_regfile_DataPath_Physical_RF_n4079,
         dp_id_stage_regfile_DataPath_Physical_RF_n4078,
         dp_id_stage_regfile_DataPath_Physical_RF_n4077,
         dp_id_stage_regfile_DataPath_Physical_RF_n4076,
         dp_id_stage_regfile_DataPath_Physical_RF_n4075,
         dp_id_stage_regfile_DataPath_Physical_RF_n4074,
         dp_id_stage_regfile_DataPath_Physical_RF_n4073,
         dp_id_stage_regfile_DataPath_Physical_RF_n4072,
         dp_id_stage_regfile_DataPath_Physical_RF_n4071,
         dp_id_stage_regfile_DataPath_Physical_RF_n4070,
         dp_id_stage_regfile_DataPath_Physical_RF_n4069,
         dp_id_stage_regfile_DataPath_Physical_RF_n4068,
         dp_id_stage_regfile_DataPath_Physical_RF_n4067,
         dp_id_stage_regfile_DataPath_Physical_RF_n4066,
         dp_id_stage_regfile_DataPath_Physical_RF_n4065,
         dp_id_stage_regfile_DataPath_Physical_RF_n4064,
         dp_id_stage_regfile_DataPath_Physical_RF_n4063,
         dp_id_stage_regfile_DataPath_Physical_RF_n4062,
         dp_id_stage_regfile_DataPath_Physical_RF_n4061,
         dp_id_stage_regfile_DataPath_Physical_RF_n4060,
         dp_id_stage_regfile_DataPath_Physical_RF_n4059,
         dp_id_stage_regfile_DataPath_Physical_RF_n4058,
         dp_id_stage_regfile_DataPath_Physical_RF_n4057,
         dp_id_stage_regfile_DataPath_Physical_RF_n4056,
         dp_id_stage_regfile_DataPath_Physical_RF_n4055,
         dp_id_stage_regfile_DataPath_Physical_RF_n4054,
         dp_id_stage_regfile_DataPath_Physical_RF_n4053,
         dp_id_stage_regfile_DataPath_Physical_RF_n4052,
         dp_id_stage_regfile_DataPath_Physical_RF_n4051,
         dp_id_stage_regfile_DataPath_Physical_RF_n4050,
         dp_id_stage_regfile_DataPath_Physical_RF_n4049,
         dp_id_stage_regfile_DataPath_Physical_RF_n4048,
         dp_id_stage_regfile_DataPath_Physical_RF_n4047,
         dp_id_stage_regfile_DataPath_Physical_RF_n4046,
         dp_id_stage_regfile_DataPath_Physical_RF_n4045,
         dp_id_stage_regfile_DataPath_Physical_RF_n4044,
         dp_id_stage_regfile_DataPath_Physical_RF_n4043,
         dp_id_stage_regfile_DataPath_Physical_RF_n4042,
         dp_id_stage_regfile_DataPath_Physical_RF_n4041,
         dp_id_stage_regfile_DataPath_Physical_RF_n4040,
         dp_id_stage_regfile_DataPath_Physical_RF_n4039,
         dp_id_stage_regfile_DataPath_Physical_RF_n4038,
         dp_id_stage_regfile_DataPath_Physical_RF_n4037,
         dp_id_stage_regfile_DataPath_Physical_RF_n4036,
         dp_id_stage_regfile_DataPath_Physical_RF_n4035,
         dp_id_stage_regfile_DataPath_Physical_RF_n4034,
         dp_id_stage_regfile_DataPath_Physical_RF_n4033,
         dp_id_stage_regfile_DataPath_Physical_RF_n4032,
         dp_id_stage_regfile_DataPath_Physical_RF_n4031,
         dp_id_stage_regfile_DataPath_Physical_RF_n4030,
         dp_id_stage_regfile_DataPath_Physical_RF_n4029,
         dp_id_stage_regfile_DataPath_Physical_RF_n4028,
         dp_id_stage_regfile_DataPath_Physical_RF_n4027,
         dp_id_stage_regfile_DataPath_Physical_RF_n4026,
         dp_id_stage_regfile_DataPath_Physical_RF_n4025,
         dp_id_stage_regfile_DataPath_Physical_RF_n4024,
         dp_id_stage_regfile_DataPath_Physical_RF_n4023,
         dp_id_stage_regfile_DataPath_Physical_RF_n4022,
         dp_id_stage_regfile_DataPath_Physical_RF_n4021,
         dp_id_stage_regfile_DataPath_Physical_RF_n4020,
         dp_id_stage_regfile_DataPath_Physical_RF_n4019,
         dp_id_stage_regfile_DataPath_Physical_RF_n4018,
         dp_id_stage_regfile_DataPath_Physical_RF_n4017,
         dp_id_stage_regfile_DataPath_Physical_RF_n4016,
         dp_id_stage_regfile_DataPath_Physical_RF_n4015,
         dp_id_stage_regfile_DataPath_Physical_RF_n4014,
         dp_id_stage_regfile_DataPath_Physical_RF_n4013,
         dp_id_stage_regfile_DataPath_Physical_RF_n4012,
         dp_id_stage_regfile_DataPath_Physical_RF_n4011,
         dp_id_stage_regfile_DataPath_Physical_RF_n4010,
         dp_id_stage_regfile_DataPath_Physical_RF_n4009,
         dp_id_stage_regfile_DataPath_Physical_RF_n4008,
         dp_id_stage_regfile_DataPath_Physical_RF_n4007,
         dp_id_stage_regfile_DataPath_Physical_RF_n4006,
         dp_id_stage_regfile_DataPath_Physical_RF_n4005,
         dp_id_stage_regfile_DataPath_Physical_RF_n4004,
         dp_id_stage_regfile_DataPath_Physical_RF_n4003,
         dp_id_stage_regfile_DataPath_Physical_RF_n4002,
         dp_id_stage_regfile_DataPath_Physical_RF_n4001,
         dp_id_stage_regfile_DataPath_Physical_RF_n4000,
         dp_id_stage_regfile_DataPath_Physical_RF_n3999,
         dp_id_stage_regfile_DataPath_Physical_RF_n3998,
         dp_id_stage_regfile_DataPath_Physical_RF_n3997,
         dp_id_stage_regfile_DataPath_Physical_RF_n3996,
         dp_id_stage_regfile_DataPath_Physical_RF_n3995,
         dp_id_stage_regfile_DataPath_Physical_RF_n3994,
         dp_id_stage_regfile_DataPath_Physical_RF_n3993,
         dp_id_stage_regfile_DataPath_Physical_RF_n3992,
         dp_id_stage_regfile_DataPath_Physical_RF_n3991,
         dp_id_stage_regfile_DataPath_Physical_RF_n3990,
         dp_id_stage_regfile_DataPath_Physical_RF_n3989,
         dp_id_stage_regfile_DataPath_Physical_RF_n3988,
         dp_id_stage_regfile_DataPath_Physical_RF_n3987,
         dp_id_stage_regfile_DataPath_Physical_RF_n3986,
         dp_id_stage_regfile_DataPath_Physical_RF_n3985,
         dp_id_stage_regfile_DataPath_Physical_RF_n3984,
         dp_id_stage_regfile_DataPath_Physical_RF_n3983,
         dp_id_stage_regfile_DataPath_Physical_RF_n3982,
         dp_id_stage_regfile_DataPath_Physical_RF_n3981,
         dp_id_stage_regfile_DataPath_Physical_RF_n3980,
         dp_id_stage_regfile_DataPath_Physical_RF_n3979,
         dp_id_stage_regfile_DataPath_Physical_RF_n3978,
         dp_id_stage_regfile_DataPath_Physical_RF_n3977,
         dp_id_stage_regfile_DataPath_Physical_RF_n3976,
         dp_id_stage_regfile_DataPath_Physical_RF_n3975,
         dp_id_stage_regfile_DataPath_Physical_RF_n3974,
         dp_id_stage_regfile_DataPath_Physical_RF_n3973,
         dp_id_stage_regfile_DataPath_Physical_RF_n3972,
         dp_id_stage_regfile_DataPath_Physical_RF_n3971,
         dp_id_stage_regfile_DataPath_Physical_RF_n3970,
         dp_id_stage_regfile_DataPath_Physical_RF_n3969,
         dp_id_stage_regfile_DataPath_Physical_RF_n3968,
         dp_id_stage_regfile_DataPath_Physical_RF_n3967,
         dp_id_stage_regfile_DataPath_Physical_RF_n3966,
         dp_id_stage_regfile_DataPath_Physical_RF_n3965,
         dp_id_stage_regfile_DataPath_Physical_RF_n3964,
         dp_id_stage_regfile_DataPath_Physical_RF_n3963,
         dp_id_stage_regfile_DataPath_Physical_RF_n3962,
         dp_id_stage_regfile_DataPath_Physical_RF_n3961,
         dp_id_stage_regfile_DataPath_Physical_RF_n3960,
         dp_id_stage_regfile_DataPath_Physical_RF_n3959,
         dp_id_stage_regfile_DataPath_Physical_RF_n3958,
         dp_id_stage_regfile_DataPath_Physical_RF_n3957,
         dp_id_stage_regfile_DataPath_Physical_RF_n3956,
         dp_id_stage_regfile_DataPath_Physical_RF_n3955,
         dp_id_stage_regfile_DataPath_Physical_RF_n3954,
         dp_id_stage_regfile_DataPath_Physical_RF_n3953,
         dp_id_stage_regfile_DataPath_Physical_RF_n3952,
         dp_id_stage_regfile_DataPath_Physical_RF_n3951,
         dp_id_stage_regfile_DataPath_Physical_RF_n3950,
         dp_id_stage_regfile_DataPath_Physical_RF_n3949,
         dp_id_stage_regfile_DataPath_Physical_RF_n3948,
         dp_id_stage_regfile_DataPath_Physical_RF_n3947,
         dp_id_stage_regfile_DataPath_Physical_RF_n3946,
         dp_id_stage_regfile_DataPath_Physical_RF_n3945,
         dp_id_stage_regfile_DataPath_Physical_RF_n3944,
         dp_id_stage_regfile_DataPath_Physical_RF_n3943,
         dp_id_stage_regfile_DataPath_Physical_RF_n3942,
         dp_id_stage_regfile_DataPath_Physical_RF_n3941,
         dp_id_stage_regfile_DataPath_Physical_RF_n3940,
         dp_id_stage_regfile_DataPath_Physical_RF_n3939,
         dp_id_stage_regfile_DataPath_Physical_RF_n3938,
         dp_id_stage_regfile_DataPath_Physical_RF_n3937,
         dp_id_stage_regfile_DataPath_Physical_RF_n3936,
         dp_id_stage_regfile_DataPath_Physical_RF_n3935,
         dp_id_stage_regfile_DataPath_Physical_RF_n3934,
         dp_id_stage_regfile_DataPath_Physical_RF_n3933,
         dp_id_stage_regfile_DataPath_Physical_RF_n3932,
         dp_id_stage_regfile_DataPath_Physical_RF_n3931,
         dp_id_stage_regfile_DataPath_Physical_RF_n3930,
         dp_id_stage_regfile_DataPath_Physical_RF_n3929,
         dp_id_stage_regfile_DataPath_Physical_RF_n3928,
         dp_id_stage_regfile_DataPath_Physical_RF_n3927,
         dp_id_stage_regfile_DataPath_Physical_RF_n3926,
         dp_id_stage_regfile_DataPath_Physical_RF_n3925,
         dp_id_stage_regfile_DataPath_Physical_RF_n3924,
         dp_id_stage_regfile_DataPath_Physical_RF_n3923,
         dp_id_stage_regfile_DataPath_Physical_RF_n3922,
         dp_id_stage_regfile_DataPath_Physical_RF_n3921,
         dp_id_stage_regfile_DataPath_Physical_RF_n3920,
         dp_id_stage_regfile_DataPath_Physical_RF_n3919,
         dp_id_stage_regfile_DataPath_Physical_RF_n3918,
         dp_id_stage_regfile_DataPath_Physical_RF_n3917,
         dp_id_stage_regfile_DataPath_Physical_RF_n3916,
         dp_id_stage_regfile_DataPath_Physical_RF_n3915,
         dp_id_stage_regfile_DataPath_Physical_RF_n3914,
         dp_id_stage_regfile_DataPath_Physical_RF_n3913,
         dp_id_stage_regfile_DataPath_Physical_RF_n3912,
         dp_id_stage_regfile_DataPath_Physical_RF_n3911,
         dp_id_stage_regfile_DataPath_Physical_RF_n3910,
         dp_id_stage_regfile_DataPath_Physical_RF_n3909,
         dp_id_stage_regfile_DataPath_Physical_RF_n3908,
         dp_id_stage_regfile_DataPath_Physical_RF_n3907,
         dp_id_stage_regfile_DataPath_Physical_RF_n3906,
         dp_id_stage_regfile_DataPath_Physical_RF_n3905,
         dp_id_stage_regfile_DataPath_Physical_RF_n3904,
         dp_id_stage_regfile_DataPath_Physical_RF_n3903,
         dp_id_stage_regfile_DataPath_Physical_RF_n3902,
         dp_id_stage_regfile_DataPath_Physical_RF_n3901,
         dp_id_stage_regfile_DataPath_Physical_RF_n3900,
         dp_id_stage_regfile_DataPath_Physical_RF_n3899,
         dp_id_stage_regfile_DataPath_Physical_RF_n3898,
         dp_id_stage_regfile_DataPath_Physical_RF_n3897,
         dp_id_stage_regfile_DataPath_Physical_RF_n3896,
         dp_id_stage_regfile_DataPath_Physical_RF_n3895,
         dp_id_stage_regfile_DataPath_Physical_RF_n3894,
         dp_id_stage_regfile_DataPath_Physical_RF_n3893,
         dp_id_stage_regfile_DataPath_Physical_RF_n3892,
         dp_id_stage_regfile_DataPath_Physical_RF_n3891,
         dp_id_stage_regfile_DataPath_Physical_RF_n3890,
         dp_id_stage_regfile_DataPath_Physical_RF_n3889,
         dp_id_stage_regfile_DataPath_Physical_RF_n3888,
         dp_id_stage_regfile_DataPath_Physical_RF_n3887,
         dp_id_stage_regfile_DataPath_Physical_RF_n3886,
         dp_id_stage_regfile_DataPath_Physical_RF_n3885,
         dp_id_stage_regfile_DataPath_Physical_RF_n3884,
         dp_id_stage_regfile_DataPath_Physical_RF_n3883,
         dp_id_stage_regfile_DataPath_Physical_RF_n3882,
         dp_id_stage_regfile_DataPath_Physical_RF_n3881,
         dp_id_stage_regfile_DataPath_Physical_RF_n3880,
         dp_id_stage_regfile_DataPath_Physical_RF_n3879,
         dp_id_stage_regfile_DataPath_Physical_RF_n3878,
         dp_id_stage_regfile_DataPath_Physical_RF_n3877,
         dp_id_stage_regfile_DataPath_Physical_RF_n3876,
         dp_id_stage_regfile_DataPath_Physical_RF_n3875,
         dp_id_stage_regfile_DataPath_Physical_RF_n3874,
         dp_id_stage_regfile_DataPath_Physical_RF_n3873,
         dp_id_stage_regfile_DataPath_Physical_RF_n3872,
         dp_id_stage_regfile_DataPath_Physical_RF_n3871,
         dp_id_stage_regfile_DataPath_Physical_RF_n3870,
         dp_id_stage_regfile_DataPath_Physical_RF_n3869,
         dp_id_stage_regfile_DataPath_Physical_RF_n3868,
         dp_id_stage_regfile_DataPath_Physical_RF_n3867,
         dp_id_stage_regfile_DataPath_Physical_RF_n3866,
         dp_id_stage_regfile_DataPath_Physical_RF_n3865,
         dp_id_stage_regfile_DataPath_Physical_RF_n3864,
         dp_id_stage_regfile_DataPath_Physical_RF_n3863,
         dp_id_stage_regfile_DataPath_Physical_RF_n3862,
         dp_id_stage_regfile_DataPath_Physical_RF_n3861,
         dp_id_stage_regfile_DataPath_Physical_RF_n3860,
         dp_id_stage_regfile_DataPath_Physical_RF_n3859,
         dp_id_stage_regfile_DataPath_Physical_RF_n3858,
         dp_id_stage_regfile_DataPath_Physical_RF_n3857,
         dp_id_stage_regfile_DataPath_Physical_RF_n3856,
         dp_id_stage_regfile_DataPath_Physical_RF_n3855,
         dp_id_stage_regfile_DataPath_Physical_RF_n3854,
         dp_id_stage_regfile_DataPath_Physical_RF_n3853,
         dp_id_stage_regfile_DataPath_Physical_RF_n3852,
         dp_id_stage_regfile_DataPath_Physical_RF_n3851,
         dp_id_stage_regfile_DataPath_Physical_RF_n3850,
         dp_id_stage_regfile_DataPath_Physical_RF_n3849,
         dp_id_stage_regfile_DataPath_Physical_RF_n3848,
         dp_id_stage_regfile_DataPath_Physical_RF_n3847,
         dp_id_stage_regfile_DataPath_Physical_RF_n3846,
         dp_id_stage_regfile_DataPath_Physical_RF_n3845,
         dp_id_stage_regfile_DataPath_Physical_RF_n3844,
         dp_id_stage_regfile_DataPath_Physical_RF_n3843,
         dp_id_stage_regfile_DataPath_Physical_RF_n3842,
         dp_id_stage_regfile_DataPath_Physical_RF_n3841,
         dp_id_stage_regfile_DataPath_Physical_RF_n3840,
         dp_id_stage_regfile_DataPath_Physical_RF_n3839,
         dp_id_stage_regfile_DataPath_Physical_RF_n3838,
         dp_id_stage_regfile_DataPath_Physical_RF_n3837,
         dp_id_stage_regfile_DataPath_Physical_RF_n3836,
         dp_id_stage_regfile_DataPath_Physical_RF_n3835,
         dp_id_stage_regfile_DataPath_Physical_RF_n3834,
         dp_id_stage_regfile_DataPath_Physical_RF_n3833,
         dp_id_stage_regfile_DataPath_Physical_RF_n3832,
         dp_id_stage_regfile_DataPath_Physical_RF_n3831,
         dp_id_stage_regfile_DataPath_Physical_RF_n3830,
         dp_id_stage_regfile_DataPath_Physical_RF_n3829,
         dp_id_stage_regfile_DataPath_Physical_RF_n3828,
         dp_id_stage_regfile_DataPath_Physical_RF_n3827,
         dp_id_stage_regfile_DataPath_Physical_RF_n3826,
         dp_id_stage_regfile_DataPath_Physical_RF_n3825,
         dp_id_stage_regfile_DataPath_Physical_RF_n3824,
         dp_id_stage_regfile_DataPath_Physical_RF_n3823,
         dp_id_stage_regfile_DataPath_Physical_RF_n3822,
         dp_id_stage_regfile_DataPath_Physical_RF_n3821,
         dp_id_stage_regfile_DataPath_Physical_RF_n3820,
         dp_id_stage_regfile_DataPath_Physical_RF_n3819,
         dp_id_stage_regfile_DataPath_Physical_RF_n3818,
         dp_id_stage_regfile_DataPath_Physical_RF_n3817,
         dp_id_stage_regfile_DataPath_Physical_RF_n3816,
         dp_id_stage_regfile_DataPath_Physical_RF_n3815,
         dp_id_stage_regfile_DataPath_Physical_RF_n3814,
         dp_id_stage_regfile_DataPath_Physical_RF_n3813,
         dp_id_stage_regfile_DataPath_Physical_RF_n3812,
         dp_id_stage_regfile_DataPath_Physical_RF_n3811,
         dp_id_stage_regfile_DataPath_Physical_RF_n3810,
         dp_id_stage_regfile_DataPath_Physical_RF_n3809,
         dp_id_stage_regfile_DataPath_Physical_RF_n3808,
         dp_id_stage_regfile_DataPath_Physical_RF_n3807,
         dp_id_stage_regfile_DataPath_Physical_RF_n3806,
         dp_id_stage_regfile_DataPath_Physical_RF_n3805,
         dp_id_stage_regfile_DataPath_Physical_RF_n3804,
         dp_id_stage_regfile_DataPath_Physical_RF_n3803,
         dp_id_stage_regfile_DataPath_Physical_RF_n3802,
         dp_id_stage_regfile_DataPath_Physical_RF_n3801,
         dp_id_stage_regfile_DataPath_Physical_RF_n3800,
         dp_id_stage_regfile_DataPath_Physical_RF_n3799,
         dp_id_stage_regfile_DataPath_Physical_RF_n3798,
         dp_id_stage_regfile_DataPath_Physical_RF_n3797,
         dp_id_stage_regfile_DataPath_Physical_RF_n3796,
         dp_id_stage_regfile_DataPath_Physical_RF_n3795,
         dp_id_stage_regfile_DataPath_Physical_RF_n3794,
         dp_id_stage_regfile_DataPath_Physical_RF_n3793,
         dp_id_stage_regfile_DataPath_Physical_RF_n3792,
         dp_id_stage_regfile_DataPath_Physical_RF_n3791,
         dp_id_stage_regfile_DataPath_Physical_RF_n3790,
         dp_id_stage_regfile_DataPath_Physical_RF_n3789,
         dp_id_stage_regfile_DataPath_Physical_RF_n3788,
         dp_id_stage_regfile_DataPath_Physical_RF_n3787,
         dp_id_stage_regfile_DataPath_Physical_RF_n3786,
         dp_id_stage_regfile_DataPath_Physical_RF_n3785,
         dp_id_stage_regfile_DataPath_Physical_RF_n3784,
         dp_id_stage_regfile_DataPath_Physical_RF_n3783,
         dp_id_stage_regfile_DataPath_Physical_RF_n3782,
         dp_id_stage_regfile_DataPath_Physical_RF_n3781,
         dp_id_stage_regfile_DataPath_Physical_RF_n3780,
         dp_id_stage_regfile_DataPath_Physical_RF_n3779,
         dp_id_stage_regfile_DataPath_Physical_RF_n3778,
         dp_id_stage_regfile_DataPath_Physical_RF_n3777,
         dp_id_stage_regfile_DataPath_Physical_RF_n3776,
         dp_id_stage_regfile_DataPath_Physical_RF_n3775,
         dp_id_stage_regfile_DataPath_Physical_RF_n3774,
         dp_id_stage_regfile_DataPath_Physical_RF_n3773,
         dp_id_stage_regfile_DataPath_Physical_RF_n3772,
         dp_id_stage_regfile_DataPath_Physical_RF_n3771,
         dp_id_stage_regfile_DataPath_Physical_RF_n3770,
         dp_id_stage_regfile_DataPath_Physical_RF_n3769,
         dp_id_stage_regfile_DataPath_Physical_RF_n3768,
         dp_id_stage_regfile_DataPath_Physical_RF_n3767,
         dp_id_stage_regfile_DataPath_Physical_RF_n3766,
         dp_id_stage_regfile_DataPath_Physical_RF_n3765,
         dp_id_stage_regfile_DataPath_Physical_RF_n3764,
         dp_id_stage_regfile_DataPath_Physical_RF_n3763,
         dp_id_stage_regfile_DataPath_Physical_RF_n3762,
         dp_id_stage_regfile_DataPath_Physical_RF_n3761,
         dp_id_stage_regfile_DataPath_Physical_RF_n3760,
         dp_id_stage_regfile_DataPath_Physical_RF_n3759,
         dp_id_stage_regfile_DataPath_Physical_RF_n3758,
         dp_id_stage_regfile_DataPath_Physical_RF_n3757,
         dp_id_stage_regfile_DataPath_Physical_RF_n3756,
         dp_id_stage_regfile_DataPath_Physical_RF_n3755,
         dp_id_stage_regfile_DataPath_Physical_RF_n3754,
         dp_id_stage_regfile_DataPath_Physical_RF_n3753,
         dp_id_stage_regfile_DataPath_Physical_RF_n3752,
         dp_id_stage_regfile_DataPath_Physical_RF_n3751,
         dp_id_stage_regfile_DataPath_Physical_RF_n3750,
         dp_id_stage_regfile_DataPath_Physical_RF_n3749,
         dp_id_stage_regfile_DataPath_Physical_RF_n3748,
         dp_id_stage_regfile_DataPath_Physical_RF_n3747,
         dp_id_stage_regfile_DataPath_Physical_RF_n3746,
         dp_id_stage_regfile_DataPath_Physical_RF_n3745,
         dp_id_stage_regfile_DataPath_Physical_RF_n3744,
         dp_id_stage_regfile_DataPath_Physical_RF_n3743,
         dp_id_stage_regfile_DataPath_Physical_RF_n3742,
         dp_id_stage_regfile_DataPath_Physical_RF_n3741,
         dp_id_stage_regfile_DataPath_Physical_RF_n3740,
         dp_id_stage_regfile_DataPath_Physical_RF_n3739,
         dp_id_stage_regfile_DataPath_Physical_RF_n3738,
         dp_id_stage_regfile_DataPath_Physical_RF_n3737,
         dp_id_stage_regfile_DataPath_Physical_RF_n3736,
         dp_id_stage_regfile_DataPath_Physical_RF_n3735,
         dp_id_stage_regfile_DataPath_Physical_RF_n3734,
         dp_id_stage_regfile_DataPath_Physical_RF_n3733,
         dp_id_stage_regfile_DataPath_Physical_RF_n3732,
         dp_id_stage_regfile_DataPath_Physical_RF_n3731,
         dp_id_stage_regfile_DataPath_Physical_RF_n3730,
         dp_id_stage_regfile_DataPath_Physical_RF_n3729,
         dp_id_stage_regfile_DataPath_Physical_RF_n3728,
         dp_id_stage_regfile_DataPath_Physical_RF_n3727,
         dp_id_stage_regfile_DataPath_Physical_RF_n3726,
         dp_id_stage_regfile_DataPath_Physical_RF_n3725,
         dp_id_stage_regfile_DataPath_Physical_RF_n3724,
         dp_id_stage_regfile_DataPath_Physical_RF_n3723,
         dp_id_stage_regfile_DataPath_Physical_RF_n3722,
         dp_id_stage_regfile_DataPath_Physical_RF_n3721,
         dp_id_stage_regfile_DataPath_Physical_RF_n3720,
         dp_id_stage_regfile_DataPath_Physical_RF_n3719,
         dp_id_stage_regfile_DataPath_Physical_RF_n3718,
         dp_id_stage_regfile_DataPath_Physical_RF_n3717,
         dp_id_stage_regfile_DataPath_Physical_RF_n3716,
         dp_id_stage_regfile_DataPath_Physical_RF_n3715,
         dp_id_stage_regfile_DataPath_Physical_RF_n3714,
         dp_id_stage_regfile_DataPath_Physical_RF_n3713,
         dp_id_stage_regfile_DataPath_Physical_RF_n3712,
         dp_id_stage_regfile_DataPath_Physical_RF_n3711,
         dp_id_stage_regfile_DataPath_Physical_RF_n3710,
         dp_id_stage_regfile_DataPath_Physical_RF_n3709,
         dp_id_stage_regfile_DataPath_Physical_RF_n3708,
         dp_id_stage_regfile_DataPath_Physical_RF_n3707,
         dp_id_stage_regfile_DataPath_Physical_RF_n3706,
         dp_id_stage_regfile_DataPath_Physical_RF_n3705,
         dp_id_stage_regfile_DataPath_Physical_RF_n3704,
         dp_id_stage_regfile_DataPath_Physical_RF_n3703,
         dp_id_stage_regfile_DataPath_Physical_RF_n3702,
         dp_id_stage_regfile_DataPath_Physical_RF_n3701,
         dp_id_stage_regfile_DataPath_Physical_RF_n3700,
         dp_id_stage_regfile_DataPath_Physical_RF_n3699,
         dp_id_stage_regfile_DataPath_Physical_RF_n3698,
         dp_id_stage_regfile_DataPath_Physical_RF_n3697,
         dp_id_stage_regfile_DataPath_Physical_RF_n3696,
         dp_id_stage_regfile_DataPath_Physical_RF_n3695,
         dp_id_stage_regfile_DataPath_Physical_RF_n3694,
         dp_id_stage_regfile_DataPath_Physical_RF_n3693,
         dp_id_stage_regfile_DataPath_Physical_RF_n1926,
         dp_id_stage_regfile_DataPath_Physical_RF_n1925,
         dp_id_stage_regfile_DataPath_Physical_RF_n1858,
         dp_id_stage_regfile_DataPath_Physical_RF_n1857,
         dp_id_stage_regfile_DataPath_Physical_RF_n1756,
         dp_id_stage_regfile_DataPath_Physical_RF_n1755,
         dp_id_stage_regfile_DataPath_Physical_RF_n1688,
         dp_id_stage_regfile_DataPath_Physical_RF_n1687,
         dp_id_stage_regfile_DataPath_Physical_RF_n1586,
         dp_id_stage_regfile_DataPath_Physical_RF_n1585,
         dp_id_stage_regfile_DataPath_Physical_RF_n1518,
         dp_id_stage_regfile_DataPath_Physical_RF_n1516,
         dp_id_stage_regfile_DataPath_Physical_RF_n1348,
         dp_id_stage_regfile_DataPath_Physical_RF_n1346,
         dp_id_stage_regfile_DataPath_Physical_RF_n1343,
         dp_id_stage_regfile_DataPath_Physical_RF_n1340,
         dp_id_stage_regfile_DataPath_Physical_RF_n1236,
         dp_id_stage_regfile_DataPath_Physical_RF_n1235,
         dp_id_stage_regfile_DataPath_Physical_RF_n1234,
         dp_id_stage_regfile_DataPath_Physical_RF_n1233,
         dp_id_stage_regfile_DataPath_Physical_RF_n1232,
         dp_id_stage_regfile_DataPath_Physical_RF_n1231,
         dp_id_stage_regfile_DataPath_Physical_RF_n1230,
         dp_id_stage_regfile_DataPath_Physical_RF_n1229,
         dp_id_stage_regfile_DataPath_Physical_RF_n1228,
         dp_id_stage_regfile_DataPath_Physical_RF_n1227,
         dp_id_stage_regfile_DataPath_Physical_RF_n1226,
         dp_id_stage_regfile_DataPath_Physical_RF_n1225,
         dp_id_stage_regfile_DataPath_Physical_RF_n1224,
         dp_id_stage_regfile_DataPath_Physical_RF_n1223,
         dp_id_stage_regfile_DataPath_Physical_RF_n1222,
         dp_id_stage_regfile_DataPath_Physical_RF_n1221,
         dp_id_stage_regfile_DataPath_Physical_RF_n1220,
         dp_id_stage_regfile_DataPath_Physical_RF_n1219,
         dp_id_stage_regfile_DataPath_Physical_RF_n1218,
         dp_id_stage_regfile_DataPath_Physical_RF_n1217,
         dp_id_stage_regfile_DataPath_Physical_RF_n1216,
         dp_id_stage_regfile_DataPath_Physical_RF_n1215,
         dp_id_stage_regfile_DataPath_Physical_RF_n1214,
         dp_id_stage_regfile_DataPath_Physical_RF_n1213,
         dp_id_stage_regfile_DataPath_Physical_RF_n1212,
         dp_id_stage_regfile_DataPath_Physical_RF_n1211,
         dp_id_stage_regfile_DataPath_Physical_RF_n1210,
         dp_id_stage_regfile_DataPath_Physical_RF_n1209,
         dp_id_stage_regfile_DataPath_Physical_RF_n1208,
         dp_id_stage_regfile_DataPath_Physical_RF_n1207,
         dp_id_stage_regfile_DataPath_Physical_RF_n1206,
         dp_id_stage_regfile_DataPath_Physical_RF_n1205,
         dp_id_stage_regfile_DataPath_Physical_RF_n1204,
         dp_id_stage_regfile_DataPath_Physical_RF_n1203,
         dp_id_stage_regfile_DataPath_Physical_RF_n1202,
         dp_id_stage_regfile_DataPath_Physical_RF_n1200,
         dp_id_stage_regfile_DataPath_Physical_RF_n1189,
         dp_id_stage_regfile_DataPath_Physical_RF_n1188,
         dp_id_stage_regfile_DataPath_Physical_RF_n1187,
         dp_id_stage_regfile_DataPath_Physical_RF_n1186,
         dp_id_stage_regfile_DataPath_Physical_RF_n1185,
         dp_id_stage_regfile_DataPath_Physical_RF_n1184,
         dp_id_stage_regfile_DataPath_Physical_RF_n1183,
         dp_id_stage_regfile_DataPath_Physical_RF_n1182,
         dp_id_stage_regfile_DataPath_Physical_RF_n1181,
         dp_id_stage_regfile_DataPath_Physical_RF_n1180,
         dp_id_stage_regfile_DataPath_Physical_RF_n1179,
         dp_id_stage_regfile_DataPath_Physical_RF_n1178,
         dp_id_stage_regfile_DataPath_Physical_RF_n1177,
         dp_id_stage_regfile_DataPath_Physical_RF_n1176,
         dp_id_stage_regfile_DataPath_Physical_RF_n1175,
         dp_id_stage_regfile_DataPath_Physical_RF_n1174,
         dp_id_stage_regfile_DataPath_Physical_RF_n1173,
         dp_id_stage_regfile_DataPath_Physical_RF_n1172,
         dp_id_stage_regfile_DataPath_Physical_RF_n1171,
         dp_id_stage_regfile_DataPath_Physical_RF_n1170,
         dp_id_stage_regfile_DataPath_Physical_RF_n1169,
         dp_id_stage_regfile_DataPath_Physical_RF_n1168,
         dp_id_stage_regfile_DataPath_Physical_RF_n1167,
         dp_id_stage_regfile_DataPath_Physical_RF_n1166,
         dp_id_stage_regfile_DataPath_Physical_RF_n1165,
         dp_id_stage_regfile_DataPath_Physical_RF_n1164,
         dp_id_stage_regfile_DataPath_Physical_RF_n1163,
         dp_id_stage_regfile_DataPath_Physical_RF_n1162,
         dp_id_stage_regfile_DataPath_Physical_RF_n1161,
         dp_id_stage_regfile_DataPath_Physical_RF_n1160,
         dp_id_stage_regfile_DataPath_Physical_RF_n1159,
         dp_id_stage_regfile_DataPath_Physical_RF_n1158,
         dp_id_stage_regfile_DataPath_Physical_RF_n1157,
         dp_id_stage_regfile_DataPath_Physical_RF_n1156,
         dp_id_stage_regfile_DataPath_Physical_RF_n1155,
         dp_id_stage_regfile_DataPath_Physical_RF_n1154,
         dp_id_stage_regfile_DataPath_Physical_RF_n1,
         dp_id_stage_regfile_DataPath_Physical_RF_n3692,
         dp_id_stage_regfile_DataPath_Physical_RF_n3691,
         dp_id_stage_regfile_DataPath_Physical_RF_n3690,
         dp_id_stage_regfile_DataPath_Physical_RF_n3689,
         dp_id_stage_regfile_DataPath_Physical_RF_n3688,
         dp_id_stage_regfile_DataPath_Physical_RF_n3687,
         dp_id_stage_regfile_DataPath_Physical_RF_n3686,
         dp_id_stage_regfile_DataPath_Physical_RF_n3685,
         dp_id_stage_regfile_DataPath_Physical_RF_n3684,
         dp_id_stage_regfile_DataPath_Physical_RF_n3683,
         dp_id_stage_regfile_DataPath_Physical_RF_n3682,
         dp_id_stage_regfile_DataPath_Physical_RF_n3681,
         dp_id_stage_regfile_DataPath_Physical_RF_n3680,
         dp_id_stage_regfile_DataPath_Physical_RF_n3679,
         dp_id_stage_regfile_DataPath_Physical_RF_n3678,
         dp_id_stage_regfile_DataPath_Physical_RF_n3677,
         dp_id_stage_regfile_DataPath_Physical_RF_n3676,
         dp_id_stage_regfile_DataPath_Physical_RF_n3675,
         dp_id_stage_regfile_DataPath_Physical_RF_n3674,
         dp_id_stage_regfile_DataPath_Physical_RF_n3673,
         dp_id_stage_regfile_DataPath_Physical_RF_n3672,
         dp_id_stage_regfile_DataPath_Physical_RF_n3671,
         dp_id_stage_regfile_DataPath_Physical_RF_n3670,
         dp_id_stage_regfile_DataPath_Physical_RF_n3669,
         dp_id_stage_regfile_DataPath_Physical_RF_n3668,
         dp_id_stage_regfile_DataPath_Physical_RF_n3667,
         dp_id_stage_regfile_DataPath_Physical_RF_n3666,
         dp_id_stage_regfile_DataPath_Physical_RF_n3665,
         dp_id_stage_regfile_DataPath_Physical_RF_n3664,
         dp_id_stage_regfile_DataPath_Physical_RF_n3663,
         dp_id_stage_regfile_DataPath_Physical_RF_n3662,
         dp_id_stage_regfile_DataPath_Physical_RF_n3661,
         dp_id_stage_regfile_DataPath_Physical_RF_n3660,
         dp_id_stage_regfile_DataPath_Physical_RF_n3659,
         dp_id_stage_regfile_DataPath_Physical_RF_n3658,
         dp_id_stage_regfile_DataPath_Physical_RF_n3657,
         dp_id_stage_regfile_DataPath_Physical_RF_n3656,
         dp_id_stage_regfile_DataPath_Physical_RF_n3655,
         dp_id_stage_regfile_DataPath_Physical_RF_n3654,
         dp_id_stage_regfile_DataPath_Physical_RF_n3653,
         dp_id_stage_regfile_DataPath_Physical_RF_n3652,
         dp_id_stage_regfile_DataPath_Physical_RF_n3651,
         dp_id_stage_regfile_DataPath_Physical_RF_n3650,
         dp_id_stage_regfile_DataPath_Physical_RF_n3649,
         dp_id_stage_regfile_DataPath_Physical_RF_n3648,
         dp_id_stage_regfile_DataPath_Physical_RF_n3647,
         dp_id_stage_regfile_DataPath_Physical_RF_n3646,
         dp_id_stage_regfile_DataPath_Physical_RF_n3645,
         dp_id_stage_regfile_DataPath_Physical_RF_n3644,
         dp_id_stage_regfile_DataPath_Physical_RF_n3643,
         dp_id_stage_regfile_DataPath_Physical_RF_n3642,
         dp_id_stage_regfile_DataPath_Physical_RF_n3641,
         dp_id_stage_regfile_DataPath_Physical_RF_n3640,
         dp_id_stage_regfile_DataPath_Physical_RF_n3639,
         dp_id_stage_regfile_DataPath_Physical_RF_n3638,
         dp_id_stage_regfile_DataPath_Physical_RF_n3637,
         dp_id_stage_regfile_DataPath_Physical_RF_n3636,
         dp_id_stage_regfile_DataPath_Physical_RF_n3635,
         dp_id_stage_regfile_DataPath_Physical_RF_n3634,
         dp_id_stage_regfile_DataPath_Physical_RF_n3633,
         dp_id_stage_regfile_DataPath_Physical_RF_n3632,
         dp_id_stage_regfile_DataPath_Physical_RF_n3631,
         dp_id_stage_regfile_DataPath_Physical_RF_n3630,
         dp_id_stage_regfile_DataPath_Physical_RF_n3629,
         dp_id_stage_regfile_DataPath_Physical_RF_n3628,
         dp_id_stage_regfile_DataPath_Physical_RF_n3627,
         dp_id_stage_regfile_DataPath_Physical_RF_n3626,
         dp_id_stage_regfile_DataPath_Physical_RF_n3625,
         dp_id_stage_regfile_DataPath_Physical_RF_n3624,
         dp_id_stage_regfile_DataPath_Physical_RF_n3623,
         dp_id_stage_regfile_DataPath_Physical_RF_n3622,
         dp_id_stage_regfile_DataPath_Physical_RF_n3621,
         dp_id_stage_regfile_DataPath_Physical_RF_n3620,
         dp_id_stage_regfile_DataPath_Physical_RF_n3619,
         dp_id_stage_regfile_DataPath_Physical_RF_n3618,
         dp_id_stage_regfile_DataPath_Physical_RF_n3617,
         dp_id_stage_regfile_DataPath_Physical_RF_n3616,
         dp_id_stage_regfile_DataPath_Physical_RF_n3615,
         dp_id_stage_regfile_DataPath_Physical_RF_n3614,
         dp_id_stage_regfile_DataPath_Physical_RF_n3613,
         dp_id_stage_regfile_DataPath_Physical_RF_n3612,
         dp_id_stage_regfile_DataPath_Physical_RF_n3611,
         dp_id_stage_regfile_DataPath_Physical_RF_n3610,
         dp_id_stage_regfile_DataPath_Physical_RF_n3609,
         dp_id_stage_regfile_DataPath_Physical_RF_n3608,
         dp_id_stage_regfile_DataPath_Physical_RF_n3607,
         dp_id_stage_regfile_DataPath_Physical_RF_n3606,
         dp_id_stage_regfile_DataPath_Physical_RF_n3605,
         dp_id_stage_regfile_DataPath_Physical_RF_n3604,
         dp_id_stage_regfile_DataPath_Physical_RF_n3603,
         dp_id_stage_regfile_DataPath_Physical_RF_n3602,
         dp_id_stage_regfile_DataPath_Physical_RF_n3601,
         dp_id_stage_regfile_DataPath_Physical_RF_n3600,
         dp_id_stage_regfile_DataPath_Physical_RF_n3599,
         dp_id_stage_regfile_DataPath_Physical_RF_n3598,
         dp_id_stage_regfile_DataPath_Physical_RF_n3597,
         dp_id_stage_regfile_DataPath_Physical_RF_n3596,
         dp_id_stage_regfile_DataPath_Physical_RF_n3595,
         dp_id_stage_regfile_DataPath_Physical_RF_n3594,
         dp_id_stage_regfile_DataPath_Physical_RF_n3593,
         dp_id_stage_regfile_DataPath_Physical_RF_n3592,
         dp_id_stage_regfile_DataPath_Physical_RF_n3591,
         dp_id_stage_regfile_DataPath_Physical_RF_n3590,
         dp_id_stage_regfile_DataPath_Physical_RF_n3589,
         dp_id_stage_regfile_DataPath_Physical_RF_n3588,
         dp_id_stage_regfile_DataPath_Physical_RF_n3587,
         dp_id_stage_regfile_DataPath_Physical_RF_n3586,
         dp_id_stage_regfile_DataPath_Physical_RF_n3585,
         dp_id_stage_regfile_DataPath_Physical_RF_n3584,
         dp_id_stage_regfile_DataPath_Physical_RF_n3583,
         dp_id_stage_regfile_DataPath_Physical_RF_n3582,
         dp_id_stage_regfile_DataPath_Physical_RF_n3581,
         dp_id_stage_regfile_DataPath_Physical_RF_n3580,
         dp_id_stage_regfile_DataPath_Physical_RF_n3579,
         dp_id_stage_regfile_DataPath_Physical_RF_n3578,
         dp_id_stage_regfile_DataPath_Physical_RF_n3577,
         dp_id_stage_regfile_DataPath_Physical_RF_n3576,
         dp_id_stage_regfile_DataPath_Physical_RF_n3575,
         dp_id_stage_regfile_DataPath_Physical_RF_n3574,
         dp_id_stage_regfile_DataPath_Physical_RF_n3573,
         dp_id_stage_regfile_DataPath_Physical_RF_n3572,
         dp_id_stage_regfile_DataPath_Physical_RF_n3571,
         dp_id_stage_regfile_DataPath_Physical_RF_n3570,
         dp_id_stage_regfile_DataPath_Physical_RF_n3569,
         dp_id_stage_regfile_DataPath_Physical_RF_n3568,
         dp_id_stage_regfile_DataPath_Physical_RF_n3567,
         dp_id_stage_regfile_DataPath_Physical_RF_n3566,
         dp_id_stage_regfile_DataPath_Physical_RF_n3565,
         dp_id_stage_regfile_DataPath_Physical_RF_n3564,
         dp_id_stage_regfile_DataPath_Physical_RF_n3563,
         dp_id_stage_regfile_DataPath_Physical_RF_n3562,
         dp_id_stage_regfile_DataPath_Physical_RF_n3561,
         dp_id_stage_regfile_DataPath_Physical_RF_n3560,
         dp_id_stage_regfile_DataPath_Physical_RF_n3559,
         dp_id_stage_regfile_DataPath_Physical_RF_n3558,
         dp_id_stage_regfile_DataPath_Physical_RF_n3557,
         dp_id_stage_regfile_DataPath_Physical_RF_n3556,
         dp_id_stage_regfile_DataPath_Physical_RF_n3555,
         dp_id_stage_regfile_DataPath_Physical_RF_n3554,
         dp_id_stage_regfile_DataPath_Physical_RF_n3553,
         dp_id_stage_regfile_DataPath_Physical_RF_n3552,
         dp_id_stage_regfile_DataPath_Physical_RF_n3551,
         dp_id_stage_regfile_DataPath_Physical_RF_n3550,
         dp_id_stage_regfile_DataPath_Physical_RF_n3549,
         dp_id_stage_regfile_DataPath_Physical_RF_n3548,
         dp_id_stage_regfile_DataPath_Physical_RF_n3547,
         dp_id_stage_regfile_DataPath_Physical_RF_n3546,
         dp_id_stage_regfile_DataPath_Physical_RF_n3545,
         dp_id_stage_regfile_DataPath_Physical_RF_n3544,
         dp_id_stage_regfile_DataPath_Physical_RF_n3543,
         dp_id_stage_regfile_DataPath_Physical_RF_n3542,
         dp_id_stage_regfile_DataPath_Physical_RF_n3541,
         dp_id_stage_regfile_DataPath_Physical_RF_n3540,
         dp_id_stage_regfile_DataPath_Physical_RF_n3539,
         dp_id_stage_regfile_DataPath_Physical_RF_n3538,
         dp_id_stage_regfile_DataPath_Physical_RF_n3537,
         dp_id_stage_regfile_DataPath_Physical_RF_n3536,
         dp_id_stage_regfile_DataPath_Physical_RF_n3535,
         dp_id_stage_regfile_DataPath_Physical_RF_n3534,
         dp_id_stage_regfile_DataPath_Physical_RF_n3533,
         dp_id_stage_regfile_DataPath_Physical_RF_n3532,
         dp_id_stage_regfile_DataPath_Physical_RF_n3531,
         dp_id_stage_regfile_DataPath_Physical_RF_n3530,
         dp_id_stage_regfile_DataPath_Physical_RF_n3529,
         dp_id_stage_regfile_DataPath_Physical_RF_n3528,
         dp_id_stage_regfile_DataPath_Physical_RF_n3527,
         dp_id_stage_regfile_DataPath_Physical_RF_n3526,
         dp_id_stage_regfile_DataPath_Physical_RF_n3525,
         dp_id_stage_regfile_DataPath_Physical_RF_n3524,
         dp_id_stage_regfile_DataPath_Physical_RF_n3523,
         dp_id_stage_regfile_DataPath_Physical_RF_n3522,
         dp_id_stage_regfile_DataPath_Physical_RF_n3521,
         dp_id_stage_regfile_DataPath_Physical_RF_n3520,
         dp_id_stage_regfile_DataPath_Physical_RF_n3519,
         dp_id_stage_regfile_DataPath_Physical_RF_n3518,
         dp_id_stage_regfile_DataPath_Physical_RF_n3517,
         dp_id_stage_regfile_DataPath_Physical_RF_n3516,
         dp_id_stage_regfile_DataPath_Physical_RF_n3515,
         dp_id_stage_regfile_DataPath_Physical_RF_n3514,
         dp_id_stage_regfile_DataPath_Physical_RF_n3513,
         dp_id_stage_regfile_DataPath_Physical_RF_n3512,
         dp_id_stage_regfile_DataPath_Physical_RF_n3511,
         dp_id_stage_regfile_DataPath_Physical_RF_n3510,
         dp_id_stage_regfile_DataPath_Physical_RF_n3509,
         dp_id_stage_regfile_DataPath_Physical_RF_n3508,
         dp_id_stage_regfile_DataPath_Physical_RF_n3507,
         dp_id_stage_regfile_DataPath_Physical_RF_n3506,
         dp_id_stage_regfile_DataPath_Physical_RF_n3505,
         dp_id_stage_regfile_DataPath_Physical_RF_n3504,
         dp_id_stage_regfile_DataPath_Physical_RF_n3503,
         dp_id_stage_regfile_DataPath_Physical_RF_n3502,
         dp_id_stage_regfile_DataPath_Physical_RF_n3501,
         dp_id_stage_regfile_DataPath_Physical_RF_n3500,
         dp_id_stage_regfile_DataPath_Physical_RF_n3499,
         dp_id_stage_regfile_DataPath_Physical_RF_n3498,
         dp_id_stage_regfile_DataPath_Physical_RF_n3497,
         dp_id_stage_regfile_DataPath_Physical_RF_n3496,
         dp_id_stage_regfile_DataPath_Physical_RF_n3495,
         dp_id_stage_regfile_DataPath_Physical_RF_n3494,
         dp_id_stage_regfile_DataPath_Physical_RF_n3493,
         dp_id_stage_regfile_DataPath_Physical_RF_n3492,
         dp_id_stage_regfile_DataPath_Physical_RF_n3491,
         dp_id_stage_regfile_DataPath_Physical_RF_n3490,
         dp_id_stage_regfile_DataPath_Physical_RF_n3489,
         dp_id_stage_regfile_DataPath_Physical_RF_n3488,
         dp_id_stage_regfile_DataPath_Physical_RF_n3487,
         dp_id_stage_regfile_DataPath_Physical_RF_n3486,
         dp_id_stage_regfile_DataPath_Physical_RF_n3485,
         dp_id_stage_regfile_DataPath_Physical_RF_n3484,
         dp_id_stage_regfile_DataPath_Physical_RF_n3483,
         dp_id_stage_regfile_DataPath_Physical_RF_n3482,
         dp_id_stage_regfile_DataPath_Physical_RF_n3481,
         dp_id_stage_regfile_DataPath_Physical_RF_n3480,
         dp_id_stage_regfile_DataPath_Physical_RF_n3479,
         dp_id_stage_regfile_DataPath_Physical_RF_n3478,
         dp_id_stage_regfile_DataPath_Physical_RF_n3477,
         dp_id_stage_regfile_DataPath_Physical_RF_n3476,
         dp_id_stage_regfile_DataPath_Physical_RF_n3475,
         dp_id_stage_regfile_DataPath_Physical_RF_n3474,
         dp_id_stage_regfile_DataPath_Physical_RF_n3473,
         dp_id_stage_regfile_DataPath_Physical_RF_n3472,
         dp_id_stage_regfile_DataPath_Physical_RF_n3471,
         dp_id_stage_regfile_DataPath_Physical_RF_n3470,
         dp_id_stage_regfile_DataPath_Physical_RF_n3469,
         dp_id_stage_regfile_DataPath_Physical_RF_n3468,
         dp_id_stage_regfile_DataPath_Physical_RF_n3467,
         dp_id_stage_regfile_DataPath_Physical_RF_n3466,
         dp_id_stage_regfile_DataPath_Physical_RF_n3465,
         dp_id_stage_regfile_DataPath_Physical_RF_n3464,
         dp_id_stage_regfile_DataPath_Physical_RF_n3463,
         dp_id_stage_regfile_DataPath_Physical_RF_n3462,
         dp_id_stage_regfile_DataPath_Physical_RF_n3461,
         dp_id_stage_regfile_DataPath_Physical_RF_n3460,
         dp_id_stage_regfile_DataPath_Physical_RF_n3459,
         dp_id_stage_regfile_DataPath_Physical_RF_n3458,
         dp_id_stage_regfile_DataPath_Physical_RF_n3457,
         dp_id_stage_regfile_DataPath_Physical_RF_n3456,
         dp_id_stage_regfile_DataPath_Physical_RF_n3455,
         dp_id_stage_regfile_DataPath_Physical_RF_n3454,
         dp_id_stage_regfile_DataPath_Physical_RF_n3453,
         dp_id_stage_regfile_DataPath_Physical_RF_n3452,
         dp_id_stage_regfile_DataPath_Physical_RF_n3451,
         dp_id_stage_regfile_DataPath_Physical_RF_n3450,
         dp_id_stage_regfile_DataPath_Physical_RF_n3449,
         dp_id_stage_regfile_DataPath_Physical_RF_n3448,
         dp_id_stage_regfile_DataPath_Physical_RF_n3447,
         dp_id_stage_regfile_DataPath_Physical_RF_n3446,
         dp_id_stage_regfile_DataPath_Physical_RF_n3445,
         dp_id_stage_regfile_DataPath_Physical_RF_n3444,
         dp_id_stage_regfile_DataPath_Physical_RF_n3443,
         dp_id_stage_regfile_DataPath_Physical_RF_n3442,
         dp_id_stage_regfile_DataPath_Physical_RF_n3441,
         dp_id_stage_regfile_DataPath_Physical_RF_n3440,
         dp_id_stage_regfile_DataPath_Physical_RF_n3439,
         dp_id_stage_regfile_DataPath_Physical_RF_n3438,
         dp_id_stage_regfile_DataPath_Physical_RF_n3437,
         dp_id_stage_regfile_DataPath_Physical_RF_n3436,
         dp_id_stage_regfile_DataPath_Physical_RF_n3435,
         dp_id_stage_regfile_DataPath_Physical_RF_n3434,
         dp_id_stage_regfile_DataPath_Physical_RF_n3433,
         dp_id_stage_regfile_DataPath_Physical_RF_n3432,
         dp_id_stage_regfile_DataPath_Physical_RF_n3431,
         dp_id_stage_regfile_DataPath_Physical_RF_n3430,
         dp_id_stage_regfile_DataPath_Physical_RF_n3429,
         dp_id_stage_regfile_DataPath_Physical_RF_n3428,
         dp_id_stage_regfile_DataPath_Physical_RF_n3427,
         dp_id_stage_regfile_DataPath_Physical_RF_n3426,
         dp_id_stage_regfile_DataPath_Physical_RF_n3425,
         dp_id_stage_regfile_DataPath_Physical_RF_n3424,
         dp_id_stage_regfile_DataPath_Physical_RF_n3423,
         dp_id_stage_regfile_DataPath_Physical_RF_n3422,
         dp_id_stage_regfile_DataPath_Physical_RF_n3421,
         dp_id_stage_regfile_DataPath_Physical_RF_n3420,
         dp_id_stage_regfile_DataPath_Physical_RF_n3419,
         dp_id_stage_regfile_DataPath_Physical_RF_n3418,
         dp_id_stage_regfile_DataPath_Physical_RF_n3417,
         dp_id_stage_regfile_DataPath_Physical_RF_n3416,
         dp_id_stage_regfile_DataPath_Physical_RF_n3415,
         dp_id_stage_regfile_DataPath_Physical_RF_n3414,
         dp_id_stage_regfile_DataPath_Physical_RF_n3413,
         dp_id_stage_regfile_DataPath_Physical_RF_n3412,
         dp_id_stage_regfile_DataPath_Physical_RF_n3411,
         dp_id_stage_regfile_DataPath_Physical_RF_n3410,
         dp_id_stage_regfile_DataPath_Physical_RF_n3409,
         dp_id_stage_regfile_DataPath_Physical_RF_n3408,
         dp_id_stage_regfile_DataPath_Physical_RF_n3407,
         dp_id_stage_regfile_DataPath_Physical_RF_n3406,
         dp_id_stage_regfile_DataPath_Physical_RF_n3405,
         dp_id_stage_regfile_DataPath_Physical_RF_n3404,
         dp_id_stage_regfile_DataPath_Physical_RF_n3403,
         dp_id_stage_regfile_DataPath_Physical_RF_n3402,
         dp_id_stage_regfile_DataPath_Physical_RF_n3401,
         dp_id_stage_regfile_DataPath_Physical_RF_n3400,
         dp_id_stage_regfile_DataPath_Physical_RF_n3399,
         dp_id_stage_regfile_DataPath_Physical_RF_n3398,
         dp_id_stage_regfile_DataPath_Physical_RF_n3397,
         dp_id_stage_regfile_DataPath_Physical_RF_n3396,
         dp_id_stage_regfile_DataPath_Physical_RF_n3395,
         dp_id_stage_regfile_DataPath_Physical_RF_n3394,
         dp_id_stage_regfile_DataPath_Physical_RF_n3393,
         dp_id_stage_regfile_DataPath_Physical_RF_n3392,
         dp_id_stage_regfile_DataPath_Physical_RF_n3391,
         dp_id_stage_regfile_DataPath_Physical_RF_n3390,
         dp_id_stage_regfile_DataPath_Physical_RF_n3389,
         dp_id_stage_regfile_DataPath_Physical_RF_n3388,
         dp_id_stage_regfile_DataPath_Physical_RF_n3387,
         dp_id_stage_regfile_DataPath_Physical_RF_n3386,
         dp_id_stage_regfile_DataPath_Physical_RF_n3385,
         dp_id_stage_regfile_DataPath_Physical_RF_n3384,
         dp_id_stage_regfile_DataPath_Physical_RF_n3383,
         dp_id_stage_regfile_DataPath_Physical_RF_n3382,
         dp_id_stage_regfile_DataPath_Physical_RF_n3381,
         dp_id_stage_regfile_DataPath_Physical_RF_n3380,
         dp_id_stage_regfile_DataPath_Physical_RF_n3379,
         dp_id_stage_regfile_DataPath_Physical_RF_n3378,
         dp_id_stage_regfile_DataPath_Physical_RF_n3377,
         dp_id_stage_regfile_DataPath_Physical_RF_n3376,
         dp_id_stage_regfile_DataPath_Physical_RF_n3375,
         dp_id_stage_regfile_DataPath_Physical_RF_n3374,
         dp_id_stage_regfile_DataPath_Physical_RF_n3373,
         dp_id_stage_regfile_DataPath_Physical_RF_n3372,
         dp_id_stage_regfile_DataPath_Physical_RF_n3371,
         dp_id_stage_regfile_DataPath_Physical_RF_n3370,
         dp_id_stage_regfile_DataPath_Physical_RF_n3369,
         dp_id_stage_regfile_DataPath_Physical_RF_n3368,
         dp_id_stage_regfile_DataPath_Physical_RF_n3367,
         dp_id_stage_regfile_DataPath_Physical_RF_n3366,
         dp_id_stage_regfile_DataPath_Physical_RF_n3365,
         dp_id_stage_regfile_DataPath_Physical_RF_n3364,
         dp_id_stage_regfile_DataPath_Physical_RF_n3363,
         dp_id_stage_regfile_DataPath_Physical_RF_n3362,
         dp_id_stage_regfile_DataPath_Physical_RF_n3361,
         dp_id_stage_regfile_DataPath_Physical_RF_n3360,
         dp_id_stage_regfile_DataPath_Physical_RF_n3359,
         dp_id_stage_regfile_DataPath_Physical_RF_n3358,
         dp_id_stage_regfile_DataPath_Physical_RF_n3357,
         dp_id_stage_regfile_DataPath_Physical_RF_n3356,
         dp_id_stage_regfile_DataPath_Physical_RF_n3355,
         dp_id_stage_regfile_DataPath_Physical_RF_n3354,
         dp_id_stage_regfile_DataPath_Physical_RF_n3353,
         dp_id_stage_regfile_DataPath_Physical_RF_n3352,
         dp_id_stage_regfile_DataPath_Physical_RF_n3351,
         dp_id_stage_regfile_DataPath_Physical_RF_n3350,
         dp_id_stage_regfile_DataPath_Physical_RF_n3349,
         dp_id_stage_regfile_DataPath_Physical_RF_n3348,
         dp_id_stage_regfile_DataPath_Physical_RF_n3347,
         dp_id_stage_regfile_DataPath_Physical_RF_n3346,
         dp_id_stage_regfile_DataPath_Physical_RF_n3345,
         dp_id_stage_regfile_DataPath_Physical_RF_n3344,
         dp_id_stage_regfile_DataPath_Physical_RF_n3343,
         dp_id_stage_regfile_DataPath_Physical_RF_n3342,
         dp_id_stage_regfile_DataPath_Physical_RF_n3341,
         dp_id_stage_regfile_DataPath_Physical_RF_n3340,
         dp_id_stage_regfile_DataPath_Physical_RF_n3339,
         dp_id_stage_regfile_DataPath_Physical_RF_n3338,
         dp_id_stage_regfile_DataPath_Physical_RF_n3337,
         dp_id_stage_regfile_DataPath_Physical_RF_n3336,
         dp_id_stage_regfile_DataPath_Physical_RF_n3335,
         dp_id_stage_regfile_DataPath_Physical_RF_n3334,
         dp_id_stage_regfile_DataPath_Physical_RF_n3333,
         dp_id_stage_regfile_DataPath_Physical_RF_n3332,
         dp_id_stage_regfile_DataPath_Physical_RF_n3331,
         dp_id_stage_regfile_DataPath_Physical_RF_n3330,
         dp_id_stage_regfile_DataPath_Physical_RF_n3329,
         dp_id_stage_regfile_DataPath_Physical_RF_n3328,
         dp_id_stage_regfile_DataPath_Physical_RF_n3327,
         dp_id_stage_regfile_DataPath_Physical_RF_n3326,
         dp_id_stage_regfile_DataPath_Physical_RF_n3325,
         dp_id_stage_regfile_DataPath_Physical_RF_n3324,
         dp_id_stage_regfile_DataPath_Physical_RF_n3323,
         dp_id_stage_regfile_DataPath_Physical_RF_n3322,
         dp_id_stage_regfile_DataPath_Physical_RF_n3321,
         dp_id_stage_regfile_DataPath_Physical_RF_n3320,
         dp_id_stage_regfile_DataPath_Physical_RF_n3319,
         dp_id_stage_regfile_DataPath_Physical_RF_n3318,
         dp_id_stage_regfile_DataPath_Physical_RF_n3317,
         dp_id_stage_regfile_DataPath_Physical_RF_n3316,
         dp_id_stage_regfile_DataPath_Physical_RF_n3315,
         dp_id_stage_regfile_DataPath_Physical_RF_n3314,
         dp_id_stage_regfile_DataPath_Physical_RF_n3313,
         dp_id_stage_regfile_DataPath_Physical_RF_n3312,
         dp_id_stage_regfile_DataPath_Physical_RF_n3311,
         dp_id_stage_regfile_DataPath_Physical_RF_n3310,
         dp_id_stage_regfile_DataPath_Physical_RF_n3309,
         dp_id_stage_regfile_DataPath_Physical_RF_n3308,
         dp_id_stage_regfile_DataPath_Physical_RF_n3307,
         dp_id_stage_regfile_DataPath_Physical_RF_n3306,
         dp_id_stage_regfile_DataPath_Physical_RF_n3305,
         dp_id_stage_regfile_DataPath_Physical_RF_n3304,
         dp_id_stage_regfile_DataPath_Physical_RF_n3303,
         dp_id_stage_regfile_DataPath_Physical_RF_n3302,
         dp_id_stage_regfile_DataPath_Physical_RF_n3301,
         dp_id_stage_regfile_DataPath_Physical_RF_n3300,
         dp_id_stage_regfile_DataPath_Physical_RF_n3299,
         dp_id_stage_regfile_DataPath_Physical_RF_n3298,
         dp_id_stage_regfile_DataPath_Physical_RF_n3297,
         dp_id_stage_regfile_DataPath_Physical_RF_n3296,
         dp_id_stage_regfile_DataPath_Physical_RF_n3295,
         dp_id_stage_regfile_DataPath_Physical_RF_n3294,
         dp_id_stage_regfile_DataPath_Physical_RF_n3293,
         dp_id_stage_regfile_DataPath_Physical_RF_n3292,
         dp_id_stage_regfile_DataPath_Physical_RF_n3291,
         dp_id_stage_regfile_DataPath_Physical_RF_n3290,
         dp_id_stage_regfile_DataPath_Physical_RF_n3289,
         dp_id_stage_regfile_DataPath_Physical_RF_n3288,
         dp_id_stage_regfile_DataPath_Physical_RF_n3287,
         dp_id_stage_regfile_DataPath_Physical_RF_n3286,
         dp_id_stage_regfile_DataPath_Physical_RF_n3285,
         dp_id_stage_regfile_DataPath_Physical_RF_n3284,
         dp_id_stage_regfile_DataPath_Physical_RF_n3283,
         dp_id_stage_regfile_DataPath_Physical_RF_n3282,
         dp_id_stage_regfile_DataPath_Physical_RF_n3281,
         dp_id_stage_regfile_DataPath_Physical_RF_n3280,
         dp_id_stage_regfile_DataPath_Physical_RF_n3279,
         dp_id_stage_regfile_DataPath_Physical_RF_n3278,
         dp_id_stage_regfile_DataPath_Physical_RF_n3277,
         dp_id_stage_regfile_DataPath_Physical_RF_n3276,
         dp_id_stage_regfile_DataPath_Physical_RF_n3275,
         dp_id_stage_regfile_DataPath_Physical_RF_n3274,
         dp_id_stage_regfile_DataPath_Physical_RF_n3273,
         dp_id_stage_regfile_DataPath_Physical_RF_n3272,
         dp_id_stage_regfile_DataPath_Physical_RF_n3271,
         dp_id_stage_regfile_DataPath_Physical_RF_n3270,
         dp_id_stage_regfile_DataPath_Physical_RF_n3269,
         dp_id_stage_regfile_DataPath_Physical_RF_n3268,
         dp_id_stage_regfile_DataPath_Physical_RF_n3267,
         dp_id_stage_regfile_DataPath_Physical_RF_n3266,
         dp_id_stage_regfile_DataPath_Physical_RF_n3265,
         dp_id_stage_regfile_DataPath_Physical_RF_n3264,
         dp_id_stage_regfile_DataPath_Physical_RF_n3263,
         dp_id_stage_regfile_DataPath_Physical_RF_n3262,
         dp_id_stage_regfile_DataPath_Physical_RF_n3261,
         dp_id_stage_regfile_DataPath_Physical_RF_n3260,
         dp_id_stage_regfile_DataPath_Physical_RF_n3259,
         dp_id_stage_regfile_DataPath_Physical_RF_n3258,
         dp_id_stage_regfile_DataPath_Physical_RF_n3257,
         dp_id_stage_regfile_DataPath_Physical_RF_n3256,
         dp_id_stage_regfile_DataPath_Physical_RF_n3255,
         dp_id_stage_regfile_DataPath_Physical_RF_n3254,
         dp_id_stage_regfile_DataPath_Physical_RF_n3253,
         dp_id_stage_regfile_DataPath_Physical_RF_n3252,
         dp_id_stage_regfile_DataPath_Physical_RF_n3251,
         dp_id_stage_regfile_DataPath_Physical_RF_n3250,
         dp_id_stage_regfile_DataPath_Physical_RF_n3249,
         dp_id_stage_regfile_DataPath_Physical_RF_n3248,
         dp_id_stage_regfile_DataPath_Physical_RF_n3247,
         dp_id_stage_regfile_DataPath_Physical_RF_n3246,
         dp_id_stage_regfile_DataPath_Physical_RF_n3245,
         dp_id_stage_regfile_DataPath_Physical_RF_n3244,
         dp_id_stage_regfile_DataPath_Physical_RF_n3243,
         dp_id_stage_regfile_DataPath_Physical_RF_n3242,
         dp_id_stage_regfile_DataPath_Physical_RF_n3241,
         dp_id_stage_regfile_DataPath_Physical_RF_n3240,
         dp_id_stage_regfile_DataPath_Physical_RF_n3239,
         dp_id_stage_regfile_DataPath_Physical_RF_n3238,
         dp_id_stage_regfile_DataPath_Physical_RF_n3237,
         dp_id_stage_regfile_DataPath_Physical_RF_n3236,
         dp_id_stage_regfile_DataPath_Physical_RF_n3235,
         dp_id_stage_regfile_DataPath_Physical_RF_n3234,
         dp_id_stage_regfile_DataPath_Physical_RF_n3233,
         dp_id_stage_regfile_DataPath_Physical_RF_n3232,
         dp_id_stage_regfile_DataPath_Physical_RF_n3231,
         dp_id_stage_regfile_DataPath_Physical_RF_n3230,
         dp_id_stage_regfile_DataPath_Physical_RF_n3229,
         dp_id_stage_regfile_DataPath_Physical_RF_n3228,
         dp_id_stage_regfile_DataPath_Physical_RF_n3227,
         dp_id_stage_regfile_DataPath_Physical_RF_n3226,
         dp_id_stage_regfile_DataPath_Physical_RF_n3225,
         dp_id_stage_regfile_DataPath_Physical_RF_n3224,
         dp_id_stage_regfile_DataPath_Physical_RF_n3223,
         dp_id_stage_regfile_DataPath_Physical_RF_n3222,
         dp_id_stage_regfile_DataPath_Physical_RF_n3221,
         dp_id_stage_regfile_DataPath_Physical_RF_n3220,
         dp_id_stage_regfile_DataPath_Physical_RF_n3219,
         dp_id_stage_regfile_DataPath_Physical_RF_n3218,
         dp_id_stage_regfile_DataPath_Physical_RF_n3217,
         dp_id_stage_regfile_DataPath_Physical_RF_n3216,
         dp_id_stage_regfile_DataPath_Physical_RF_n3215,
         dp_id_stage_regfile_DataPath_Physical_RF_n3214,
         dp_id_stage_regfile_DataPath_Physical_RF_n3213,
         dp_id_stage_regfile_DataPath_Physical_RF_n3212,
         dp_id_stage_regfile_DataPath_Physical_RF_n3211,
         dp_id_stage_regfile_DataPath_Physical_RF_n3210,
         dp_id_stage_regfile_DataPath_Physical_RF_n3209,
         dp_id_stage_regfile_DataPath_Physical_RF_n3208,
         dp_id_stage_regfile_DataPath_Physical_RF_n3207,
         dp_id_stage_regfile_DataPath_Physical_RF_n3206,
         dp_id_stage_regfile_DataPath_Physical_RF_n3205,
         dp_id_stage_regfile_DataPath_Physical_RF_n3204,
         dp_id_stage_regfile_DataPath_Physical_RF_n3203,
         dp_id_stage_regfile_DataPath_Physical_RF_n3202,
         dp_id_stage_regfile_DataPath_Physical_RF_n3201,
         dp_id_stage_regfile_DataPath_Physical_RF_n3200,
         dp_id_stage_regfile_DataPath_Physical_RF_n3199,
         dp_id_stage_regfile_DataPath_Physical_RF_n3198,
         dp_id_stage_regfile_DataPath_Physical_RF_n3197,
         dp_id_stage_regfile_DataPath_Physical_RF_n3196,
         dp_id_stage_regfile_DataPath_Physical_RF_n3195,
         dp_id_stage_regfile_DataPath_Physical_RF_n3194,
         dp_id_stage_regfile_DataPath_Physical_RF_n3193,
         dp_id_stage_regfile_DataPath_Physical_RF_n3192,
         dp_id_stage_regfile_DataPath_Physical_RF_n3191,
         dp_id_stage_regfile_DataPath_Physical_RF_n3190,
         dp_id_stage_regfile_DataPath_Physical_RF_n3189,
         dp_id_stage_regfile_DataPath_Physical_RF_n3188,
         dp_id_stage_regfile_DataPath_Physical_RF_n3187,
         dp_id_stage_regfile_DataPath_Physical_RF_n3186,
         dp_id_stage_regfile_DataPath_Physical_RF_n3185,
         dp_id_stage_regfile_DataPath_Physical_RF_n3184,
         dp_id_stage_regfile_DataPath_Physical_RF_n3183,
         dp_id_stage_regfile_DataPath_Physical_RF_n3182,
         dp_id_stage_regfile_DataPath_Physical_RF_n3181,
         dp_id_stage_regfile_DataPath_Physical_RF_n3180,
         dp_id_stage_regfile_DataPath_Physical_RF_n3179,
         dp_id_stage_regfile_DataPath_Physical_RF_n3178,
         dp_id_stage_regfile_DataPath_Physical_RF_n3177,
         dp_id_stage_regfile_DataPath_Physical_RF_n3176,
         dp_id_stage_regfile_DataPath_Physical_RF_n3175,
         dp_id_stage_regfile_DataPath_Physical_RF_n3174,
         dp_id_stage_regfile_DataPath_Physical_RF_n3173,
         dp_id_stage_regfile_DataPath_Physical_RF_n3172,
         dp_id_stage_regfile_DataPath_Physical_RF_n3171,
         dp_id_stage_regfile_DataPath_Physical_RF_n3170,
         dp_id_stage_regfile_DataPath_Physical_RF_n3169,
         dp_id_stage_regfile_DataPath_Physical_RF_n3168,
         dp_id_stage_regfile_DataPath_Physical_RF_n3167,
         dp_id_stage_regfile_DataPath_Physical_RF_n3166,
         dp_id_stage_regfile_DataPath_Physical_RF_n3165,
         dp_id_stage_regfile_DataPath_Physical_RF_n3164,
         dp_id_stage_regfile_DataPath_Physical_RF_n3163,
         dp_id_stage_regfile_DataPath_Physical_RF_n3162,
         dp_id_stage_regfile_DataPath_Physical_RF_n3161,
         dp_id_stage_regfile_DataPath_Physical_RF_n3160,
         dp_id_stage_regfile_DataPath_Physical_RF_n3159,
         dp_id_stage_regfile_DataPath_Physical_RF_n3158,
         dp_id_stage_regfile_DataPath_Physical_RF_n3157,
         dp_id_stage_regfile_DataPath_Physical_RF_n3156,
         dp_id_stage_regfile_DataPath_Physical_RF_n3155,
         dp_id_stage_regfile_DataPath_Physical_RF_n3154,
         dp_id_stage_regfile_DataPath_Physical_RF_n3153,
         dp_id_stage_regfile_DataPath_Physical_RF_n3152,
         dp_id_stage_regfile_DataPath_Physical_RF_n3151,
         dp_id_stage_regfile_DataPath_Physical_RF_n3150,
         dp_id_stage_regfile_DataPath_Physical_RF_n3149,
         dp_id_stage_regfile_DataPath_Physical_RF_n3148,
         dp_id_stage_regfile_DataPath_Physical_RF_n3147,
         dp_id_stage_regfile_DataPath_Physical_RF_n3146,
         dp_id_stage_regfile_DataPath_Physical_RF_n3145,
         dp_id_stage_regfile_DataPath_Physical_RF_n3144,
         dp_id_stage_regfile_DataPath_Physical_RF_n3143,
         dp_id_stage_regfile_DataPath_Physical_RF_n3142,
         dp_id_stage_regfile_DataPath_Physical_RF_n3141,
         dp_id_stage_regfile_DataPath_Physical_RF_n3140,
         dp_id_stage_regfile_DataPath_Physical_RF_n3139,
         dp_id_stage_regfile_DataPath_Physical_RF_n3138,
         dp_id_stage_regfile_DataPath_Physical_RF_n3137,
         dp_id_stage_regfile_DataPath_Physical_RF_n3136,
         dp_id_stage_regfile_DataPath_Physical_RF_n3135,
         dp_id_stage_regfile_DataPath_Physical_RF_n3134,
         dp_id_stage_regfile_DataPath_Physical_RF_n3133,
         dp_id_stage_regfile_DataPath_Physical_RF_n3132,
         dp_id_stage_regfile_DataPath_Physical_RF_n3131,
         dp_id_stage_regfile_DataPath_Physical_RF_n3130,
         dp_id_stage_regfile_DataPath_Physical_RF_n3129,
         dp_id_stage_regfile_DataPath_Physical_RF_n3128,
         dp_id_stage_regfile_DataPath_Physical_RF_n3127,
         dp_id_stage_regfile_DataPath_Physical_RF_n3126,
         dp_id_stage_regfile_DataPath_Physical_RF_n3125,
         dp_id_stage_regfile_DataPath_Physical_RF_n3124,
         dp_id_stage_regfile_DataPath_Physical_RF_n3123,
         dp_id_stage_regfile_DataPath_Physical_RF_n3122,
         dp_id_stage_regfile_DataPath_Physical_RF_n3121,
         dp_id_stage_regfile_DataPath_Physical_RF_n3120,
         dp_id_stage_regfile_DataPath_Physical_RF_n3119,
         dp_id_stage_regfile_DataPath_Physical_RF_n3118,
         dp_id_stage_regfile_DataPath_Physical_RF_n3117,
         dp_id_stage_regfile_DataPath_Physical_RF_n3116,
         dp_id_stage_regfile_DataPath_Physical_RF_n3115,
         dp_id_stage_regfile_DataPath_Physical_RF_n3114,
         dp_id_stage_regfile_DataPath_Physical_RF_n3113,
         dp_id_stage_regfile_DataPath_Physical_RF_n3112,
         dp_id_stage_regfile_DataPath_Physical_RF_n3111,
         dp_id_stage_regfile_DataPath_Physical_RF_n3110,
         dp_id_stage_regfile_DataPath_Physical_RF_n3109,
         dp_id_stage_regfile_DataPath_Physical_RF_n3108,
         dp_id_stage_regfile_DataPath_Physical_RF_n3107,
         dp_id_stage_regfile_DataPath_Physical_RF_n3106,
         dp_id_stage_regfile_DataPath_Physical_RF_n3105,
         dp_id_stage_regfile_DataPath_Physical_RF_n3104,
         dp_id_stage_regfile_DataPath_Physical_RF_n3103,
         dp_id_stage_regfile_DataPath_Physical_RF_n3102,
         dp_id_stage_regfile_DataPath_Physical_RF_n3101,
         dp_id_stage_regfile_DataPath_Physical_RF_n3100,
         dp_id_stage_regfile_DataPath_Physical_RF_n3099,
         dp_id_stage_regfile_DataPath_Physical_RF_n3098,
         dp_id_stage_regfile_DataPath_Physical_RF_n3097,
         dp_id_stage_regfile_DataPath_Physical_RF_n3096,
         dp_id_stage_regfile_DataPath_Physical_RF_n3095,
         dp_id_stage_regfile_DataPath_Physical_RF_n3094,
         dp_id_stage_regfile_DataPath_Physical_RF_n3093,
         dp_id_stage_regfile_DataPath_Physical_RF_n3092,
         dp_id_stage_regfile_DataPath_Physical_RF_n3091,
         dp_id_stage_regfile_DataPath_Physical_RF_n3090,
         dp_id_stage_regfile_DataPath_Physical_RF_n3089,
         dp_id_stage_regfile_DataPath_Physical_RF_n3088,
         dp_id_stage_regfile_DataPath_Physical_RF_n3087,
         dp_id_stage_regfile_DataPath_Physical_RF_n3086,
         dp_id_stage_regfile_DataPath_Physical_RF_n3085,
         dp_id_stage_regfile_DataPath_Physical_RF_n3084,
         dp_id_stage_regfile_DataPath_Physical_RF_n3083,
         dp_id_stage_regfile_DataPath_Physical_RF_n3082,
         dp_id_stage_regfile_DataPath_Physical_RF_n3081,
         dp_id_stage_regfile_DataPath_Physical_RF_n3080,
         dp_id_stage_regfile_DataPath_Physical_RF_n3079,
         dp_id_stage_regfile_DataPath_Physical_RF_n3078,
         dp_id_stage_regfile_DataPath_Physical_RF_n3077,
         dp_id_stage_regfile_DataPath_Physical_RF_n3076,
         dp_id_stage_regfile_DataPath_Physical_RF_n3075,
         dp_id_stage_regfile_DataPath_Physical_RF_n3074,
         dp_id_stage_regfile_DataPath_Physical_RF_n3073,
         dp_id_stage_regfile_DataPath_Physical_RF_n3072,
         dp_id_stage_regfile_DataPath_Physical_RF_n3071,
         dp_id_stage_regfile_DataPath_Physical_RF_n3070,
         dp_id_stage_regfile_DataPath_Physical_RF_n3069,
         dp_id_stage_regfile_DataPath_Physical_RF_n3068,
         dp_id_stage_regfile_DataPath_Physical_RF_n3067,
         dp_id_stage_regfile_DataPath_Physical_RF_n3066,
         dp_id_stage_regfile_DataPath_Physical_RF_n3065,
         dp_id_stage_regfile_DataPath_Physical_RF_n3064,
         dp_id_stage_regfile_DataPath_Physical_RF_n3063,
         dp_id_stage_regfile_DataPath_Physical_RF_n3062,
         dp_id_stage_regfile_DataPath_Physical_RF_n3061,
         dp_id_stage_regfile_DataPath_Physical_RF_n3060,
         dp_id_stage_regfile_DataPath_Physical_RF_n3059,
         dp_id_stage_regfile_DataPath_Physical_RF_n3058,
         dp_id_stage_regfile_DataPath_Physical_RF_n3057,
         dp_id_stage_regfile_DataPath_Physical_RF_n3056,
         dp_id_stage_regfile_DataPath_Physical_RF_n3055,
         dp_id_stage_regfile_DataPath_Physical_RF_n3054,
         dp_id_stage_regfile_DataPath_Physical_RF_n3053,
         dp_id_stage_regfile_DataPath_Physical_RF_n3052,
         dp_id_stage_regfile_DataPath_Physical_RF_n3051,
         dp_id_stage_regfile_DataPath_Physical_RF_n3050,
         dp_id_stage_regfile_DataPath_Physical_RF_n3049,
         dp_id_stage_regfile_DataPath_Physical_RF_n3048,
         dp_id_stage_regfile_DataPath_Physical_RF_n3047,
         dp_id_stage_regfile_DataPath_Physical_RF_n3046,
         dp_id_stage_regfile_DataPath_Physical_RF_n3045,
         dp_id_stage_regfile_DataPath_Physical_RF_n3044,
         dp_id_stage_regfile_DataPath_Physical_RF_n3043,
         dp_id_stage_regfile_DataPath_Physical_RF_n3042,
         dp_id_stage_regfile_DataPath_Physical_RF_n3041,
         dp_id_stage_regfile_DataPath_Physical_RF_n3040,
         dp_id_stage_regfile_DataPath_Physical_RF_n3039,
         dp_id_stage_regfile_DataPath_Physical_RF_n3038,
         dp_id_stage_regfile_DataPath_Physical_RF_n3037,
         dp_id_stage_regfile_DataPath_Physical_RF_n3036,
         dp_id_stage_regfile_DataPath_Physical_RF_n3035,
         dp_id_stage_regfile_DataPath_Physical_RF_n3034,
         dp_id_stage_regfile_DataPath_Physical_RF_n3033,
         dp_id_stage_regfile_DataPath_Physical_RF_n3032,
         dp_id_stage_regfile_DataPath_Physical_RF_n3031,
         dp_id_stage_regfile_DataPath_Physical_RF_n3030,
         dp_id_stage_regfile_DataPath_Physical_RF_n3029,
         dp_id_stage_regfile_DataPath_Physical_RF_n3028,
         dp_id_stage_regfile_DataPath_Physical_RF_n3027,
         dp_id_stage_regfile_DataPath_Physical_RF_n3026,
         dp_id_stage_regfile_DataPath_Physical_RF_n3025,
         dp_id_stage_regfile_DataPath_Physical_RF_n3024,
         dp_id_stage_regfile_DataPath_Physical_RF_n3023,
         dp_id_stage_regfile_DataPath_Physical_RF_n3022,
         dp_id_stage_regfile_DataPath_Physical_RF_n3021,
         dp_id_stage_regfile_DataPath_Physical_RF_n3020,
         dp_id_stage_regfile_DataPath_Physical_RF_n3019,
         dp_id_stage_regfile_DataPath_Physical_RF_n3018,
         dp_id_stage_regfile_DataPath_Physical_RF_n3017,
         dp_id_stage_regfile_DataPath_Physical_RF_n3016,
         dp_id_stage_regfile_DataPath_Physical_RF_n3015,
         dp_id_stage_regfile_DataPath_Physical_RF_n3014,
         dp_id_stage_regfile_DataPath_Physical_RF_n3013,
         dp_id_stage_regfile_DataPath_Physical_RF_n3012,
         dp_id_stage_regfile_DataPath_Physical_RF_n3011,
         dp_id_stage_regfile_DataPath_Physical_RF_n3010,
         dp_id_stage_regfile_DataPath_Physical_RF_n3009,
         dp_id_stage_regfile_DataPath_Physical_RF_n3008,
         dp_id_stage_regfile_DataPath_Physical_RF_n3007,
         dp_id_stage_regfile_DataPath_Physical_RF_n3006,
         dp_id_stage_regfile_DataPath_Physical_RF_n3005,
         dp_id_stage_regfile_DataPath_Physical_RF_n3004,
         dp_id_stage_regfile_DataPath_Physical_RF_n3003,
         dp_id_stage_regfile_DataPath_Physical_RF_n3002,
         dp_id_stage_regfile_DataPath_Physical_RF_n3001,
         dp_id_stage_regfile_DataPath_Physical_RF_n3000,
         dp_id_stage_regfile_DataPath_Physical_RF_n2999,
         dp_id_stage_regfile_DataPath_Physical_RF_n2998,
         dp_id_stage_regfile_DataPath_Physical_RF_n2997,
         dp_id_stage_regfile_DataPath_Physical_RF_n2996,
         dp_id_stage_regfile_DataPath_Physical_RF_n2995,
         dp_id_stage_regfile_DataPath_Physical_RF_n2994,
         dp_id_stage_regfile_DataPath_Physical_RF_n2993,
         dp_id_stage_regfile_DataPath_Physical_RF_n2992,
         dp_id_stage_regfile_DataPath_Physical_RF_n2991,
         dp_id_stage_regfile_DataPath_Physical_RF_n2990,
         dp_id_stage_regfile_DataPath_Physical_RF_n2989,
         dp_id_stage_regfile_DataPath_Physical_RF_n2988,
         dp_id_stage_regfile_DataPath_Physical_RF_n2987,
         dp_id_stage_regfile_DataPath_Physical_RF_n2986,
         dp_id_stage_regfile_DataPath_Physical_RF_n2985,
         dp_id_stage_regfile_DataPath_Physical_RF_n2984,
         dp_id_stage_regfile_DataPath_Physical_RF_n2983,
         dp_id_stage_regfile_DataPath_Physical_RF_n2982,
         dp_id_stage_regfile_DataPath_Physical_RF_n2981,
         dp_id_stage_regfile_DataPath_Physical_RF_n2980,
         dp_id_stage_regfile_DataPath_Physical_RF_n2979,
         dp_id_stage_regfile_DataPath_Physical_RF_n2978,
         dp_id_stage_regfile_DataPath_Physical_RF_n2977,
         dp_id_stage_regfile_DataPath_Physical_RF_n2976,
         dp_id_stage_regfile_DataPath_Physical_RF_n2975,
         dp_id_stage_regfile_DataPath_Physical_RF_n2974,
         dp_id_stage_regfile_DataPath_Physical_RF_n2973,
         dp_id_stage_regfile_DataPath_Physical_RF_n2972,
         dp_id_stage_regfile_DataPath_Physical_RF_n2971,
         dp_id_stage_regfile_DataPath_Physical_RF_n2970,
         dp_id_stage_regfile_DataPath_Physical_RF_n2969,
         dp_id_stage_regfile_DataPath_Physical_RF_n2968,
         dp_id_stage_regfile_DataPath_Physical_RF_n2967,
         dp_id_stage_regfile_DataPath_Physical_RF_n2966,
         dp_id_stage_regfile_DataPath_Physical_RF_n2965,
         dp_id_stage_regfile_DataPath_Physical_RF_n2964,
         dp_id_stage_regfile_DataPath_Physical_RF_n2963,
         dp_id_stage_regfile_DataPath_Physical_RF_n2962,
         dp_id_stage_regfile_DataPath_Physical_RF_n2961,
         dp_id_stage_regfile_DataPath_Physical_RF_n2960,
         dp_id_stage_regfile_DataPath_Physical_RF_n2959,
         dp_id_stage_regfile_DataPath_Physical_RF_n2958,
         dp_id_stage_regfile_DataPath_Physical_RF_n2957,
         dp_id_stage_regfile_DataPath_Physical_RF_n2956,
         dp_id_stage_regfile_DataPath_Physical_RF_n2955,
         dp_id_stage_regfile_DataPath_Physical_RF_n2954,
         dp_id_stage_regfile_DataPath_Physical_RF_n2953,
         dp_id_stage_regfile_DataPath_Physical_RF_n2952,
         dp_id_stage_regfile_DataPath_Physical_RF_n2951,
         dp_id_stage_regfile_DataPath_Physical_RF_n2950,
         dp_id_stage_regfile_DataPath_Physical_RF_n2949,
         dp_id_stage_regfile_DataPath_Physical_RF_n2948,
         dp_id_stage_regfile_DataPath_Physical_RF_n2947,
         dp_id_stage_regfile_DataPath_Physical_RF_n2946,
         dp_id_stage_regfile_DataPath_Physical_RF_n2945,
         dp_id_stage_regfile_DataPath_Physical_RF_n2944,
         dp_id_stage_regfile_DataPath_Physical_RF_n2943,
         dp_id_stage_regfile_DataPath_Physical_RF_n2942,
         dp_id_stage_regfile_DataPath_Physical_RF_n2941,
         dp_id_stage_regfile_DataPath_Physical_RF_n2940,
         dp_id_stage_regfile_DataPath_Physical_RF_n2939,
         dp_id_stage_regfile_DataPath_Physical_RF_n2938,
         dp_id_stage_regfile_DataPath_Physical_RF_n2937,
         dp_id_stage_regfile_DataPath_Physical_RF_n2936,
         dp_id_stage_regfile_DataPath_Physical_RF_n2935,
         dp_id_stage_regfile_DataPath_Physical_RF_n2934,
         dp_id_stage_regfile_DataPath_Physical_RF_n2933,
         dp_id_stage_regfile_DataPath_Physical_RF_n2932,
         dp_id_stage_regfile_DataPath_Physical_RF_n2931,
         dp_id_stage_regfile_DataPath_Physical_RF_n2930,
         dp_id_stage_regfile_DataPath_Physical_RF_n2929,
         dp_id_stage_regfile_DataPath_Physical_RF_n2928,
         dp_id_stage_regfile_DataPath_Physical_RF_n2927,
         dp_id_stage_regfile_DataPath_Physical_RF_n2926,
         dp_id_stage_regfile_DataPath_Physical_RF_n2925,
         dp_id_stage_regfile_DataPath_Physical_RF_n2924,
         dp_id_stage_regfile_DataPath_Physical_RF_n2923,
         dp_id_stage_regfile_DataPath_Physical_RF_n2922,
         dp_id_stage_regfile_DataPath_Physical_RF_n2921,
         dp_id_stage_regfile_DataPath_Physical_RF_n2920,
         dp_id_stage_regfile_DataPath_Physical_RF_n2919,
         dp_id_stage_regfile_DataPath_Physical_RF_n2918,
         dp_id_stage_regfile_DataPath_Physical_RF_n2917,
         dp_id_stage_regfile_DataPath_Physical_RF_n2916,
         dp_id_stage_regfile_DataPath_Physical_RF_n2915,
         dp_id_stage_regfile_DataPath_Physical_RF_n2914,
         dp_id_stage_regfile_DataPath_Physical_RF_n2913,
         dp_id_stage_regfile_DataPath_Physical_RF_n2912,
         dp_id_stage_regfile_DataPath_Physical_RF_n2911,
         dp_id_stage_regfile_DataPath_Physical_RF_n2910,
         dp_id_stage_regfile_DataPath_Physical_RF_n2909,
         dp_id_stage_regfile_DataPath_Physical_RF_n2908,
         dp_id_stage_regfile_DataPath_Physical_RF_n2907,
         dp_id_stage_regfile_DataPath_Physical_RF_n2906,
         dp_id_stage_regfile_DataPath_Physical_RF_n2905,
         dp_id_stage_regfile_DataPath_Physical_RF_n2904,
         dp_id_stage_regfile_DataPath_Physical_RF_n2903,
         dp_id_stage_regfile_DataPath_Physical_RF_n2902,
         dp_id_stage_regfile_DataPath_Physical_RF_n2901,
         dp_id_stage_regfile_DataPath_Physical_RF_n2900,
         dp_id_stage_regfile_DataPath_Physical_RF_n2899,
         dp_id_stage_regfile_DataPath_Physical_RF_n2898,
         dp_id_stage_regfile_DataPath_Physical_RF_n2897,
         dp_id_stage_regfile_DataPath_Physical_RF_n2896,
         dp_id_stage_regfile_DataPath_Physical_RF_n2895,
         dp_id_stage_regfile_DataPath_Physical_RF_n2894,
         dp_id_stage_regfile_DataPath_Physical_RF_n2893,
         dp_id_stage_regfile_DataPath_Physical_RF_n2892,
         dp_id_stage_regfile_DataPath_Physical_RF_n2891,
         dp_id_stage_regfile_DataPath_Physical_RF_n2890,
         dp_id_stage_regfile_DataPath_Physical_RF_n2889,
         dp_id_stage_regfile_DataPath_Physical_RF_n2888,
         dp_id_stage_regfile_DataPath_Physical_RF_n2887,
         dp_id_stage_regfile_DataPath_Physical_RF_n2886,
         dp_id_stage_regfile_DataPath_Physical_RF_n2885,
         dp_id_stage_regfile_DataPath_Physical_RF_n2884,
         dp_id_stage_regfile_DataPath_Physical_RF_n2883,
         dp_id_stage_regfile_DataPath_Physical_RF_n2882,
         dp_id_stage_regfile_DataPath_Physical_RF_n2881,
         dp_id_stage_regfile_DataPath_Physical_RF_n2880,
         dp_id_stage_regfile_DataPath_Physical_RF_n2879,
         dp_id_stage_regfile_DataPath_Physical_RF_n2878,
         dp_id_stage_regfile_DataPath_Physical_RF_n2877,
         dp_id_stage_regfile_DataPath_Physical_RF_n2876,
         dp_id_stage_regfile_DataPath_Physical_RF_n2875,
         dp_id_stage_regfile_DataPath_Physical_RF_n2874,
         dp_id_stage_regfile_DataPath_Physical_RF_n2873,
         dp_id_stage_regfile_DataPath_Physical_RF_n2872,
         dp_id_stage_regfile_DataPath_Physical_RF_n2871,
         dp_id_stage_regfile_DataPath_Physical_RF_n2870,
         dp_id_stage_regfile_DataPath_Physical_RF_n2869,
         dp_id_stage_regfile_DataPath_Physical_RF_n2868,
         dp_id_stage_regfile_DataPath_Physical_RF_n2867,
         dp_id_stage_regfile_DataPath_Physical_RF_n2866,
         dp_id_stage_regfile_DataPath_Physical_RF_n2865,
         dp_id_stage_regfile_DataPath_Physical_RF_n2864,
         dp_id_stage_regfile_DataPath_Physical_RF_n2863,
         dp_id_stage_regfile_DataPath_Physical_RF_n2862,
         dp_id_stage_regfile_DataPath_Physical_RF_n2861,
         dp_id_stage_regfile_DataPath_Physical_RF_n2860,
         dp_id_stage_regfile_DataPath_Physical_RF_n2859,
         dp_id_stage_regfile_DataPath_Physical_RF_n2858,
         dp_id_stage_regfile_DataPath_Physical_RF_n2857,
         dp_id_stage_regfile_DataPath_Physical_RF_n2856,
         dp_id_stage_regfile_DataPath_Physical_RF_n2855,
         dp_id_stage_regfile_DataPath_Physical_RF_n2854,
         dp_id_stage_regfile_DataPath_Physical_RF_n2853,
         dp_id_stage_regfile_DataPath_Physical_RF_n2852,
         dp_id_stage_regfile_DataPath_Physical_RF_n2851,
         dp_id_stage_regfile_DataPath_Physical_RF_n2850,
         dp_id_stage_regfile_DataPath_Physical_RF_n2849,
         dp_id_stage_regfile_DataPath_Physical_RF_n2848,
         dp_id_stage_regfile_DataPath_Physical_RF_n2847,
         dp_id_stage_regfile_DataPath_Physical_RF_n2846,
         dp_id_stage_regfile_DataPath_Physical_RF_n2845,
         dp_id_stage_regfile_DataPath_Physical_RF_n2844,
         dp_id_stage_regfile_DataPath_Physical_RF_n2843,
         dp_id_stage_regfile_DataPath_Physical_RF_n2842,
         dp_id_stage_regfile_DataPath_Physical_RF_n2841,
         dp_id_stage_regfile_DataPath_Physical_RF_n2840,
         dp_id_stage_regfile_DataPath_Physical_RF_n2839,
         dp_id_stage_regfile_DataPath_Physical_RF_n2838,
         dp_id_stage_regfile_DataPath_Physical_RF_n2837,
         dp_id_stage_regfile_DataPath_Physical_RF_n2836,
         dp_id_stage_regfile_DataPath_Physical_RF_n2835,
         dp_id_stage_regfile_DataPath_Physical_RF_n2834,
         dp_id_stage_regfile_DataPath_Physical_RF_n2833,
         dp_id_stage_regfile_DataPath_Physical_RF_n2832,
         dp_id_stage_regfile_DataPath_Physical_RF_n2831,
         dp_id_stage_regfile_DataPath_Physical_RF_n2830,
         dp_id_stage_regfile_DataPath_Physical_RF_n2829,
         dp_id_stage_regfile_DataPath_Physical_RF_n2828,
         dp_id_stage_regfile_DataPath_Physical_RF_n2827,
         dp_id_stage_regfile_DataPath_Physical_RF_n2826,
         dp_id_stage_regfile_DataPath_Physical_RF_n2825,
         dp_id_stage_regfile_DataPath_Physical_RF_n2824,
         dp_id_stage_regfile_DataPath_Physical_RF_n2823,
         dp_id_stage_regfile_DataPath_Physical_RF_n2822,
         dp_id_stage_regfile_DataPath_Physical_RF_n2821,
         dp_id_stage_regfile_DataPath_Physical_RF_n2820,
         dp_id_stage_regfile_DataPath_Physical_RF_n2819,
         dp_id_stage_regfile_DataPath_Physical_RF_n2818,
         dp_id_stage_regfile_DataPath_Physical_RF_n2817,
         dp_id_stage_regfile_DataPath_Physical_RF_n2816,
         dp_id_stage_regfile_DataPath_Physical_RF_n2815,
         dp_id_stage_regfile_DataPath_Physical_RF_n2814,
         dp_id_stage_regfile_DataPath_Physical_RF_n2813,
         dp_id_stage_regfile_DataPath_Physical_RF_n2812,
         dp_id_stage_regfile_DataPath_Physical_RF_n2811,
         dp_id_stage_regfile_DataPath_Physical_RF_n2810,
         dp_id_stage_regfile_DataPath_Physical_RF_n2809,
         dp_id_stage_regfile_DataPath_Physical_RF_n2808,
         dp_id_stage_regfile_DataPath_Physical_RF_n2807,
         dp_id_stage_regfile_DataPath_Physical_RF_n2806,
         dp_id_stage_regfile_DataPath_Physical_RF_n2805,
         dp_id_stage_regfile_DataPath_Physical_RF_n2804,
         dp_id_stage_regfile_DataPath_Physical_RF_n2803,
         dp_id_stage_regfile_DataPath_Physical_RF_n2802,
         dp_id_stage_regfile_DataPath_Physical_RF_n2801,
         dp_id_stage_regfile_DataPath_Physical_RF_n2800,
         dp_id_stage_regfile_DataPath_Physical_RF_n2799,
         dp_id_stage_regfile_DataPath_Physical_RF_n2798,
         dp_id_stage_regfile_DataPath_Physical_RF_n2797,
         dp_id_stage_regfile_DataPath_Physical_RF_n2796,
         dp_id_stage_regfile_DataPath_Physical_RF_n2795,
         dp_id_stage_regfile_DataPath_Physical_RF_n2794,
         dp_id_stage_regfile_DataPath_Physical_RF_n2793,
         dp_id_stage_regfile_DataPath_Physical_RF_n2792,
         dp_id_stage_regfile_DataPath_Physical_RF_n2791,
         dp_id_stage_regfile_DataPath_Physical_RF_n2790,
         dp_id_stage_regfile_DataPath_Physical_RF_n2789,
         dp_id_stage_regfile_DataPath_Physical_RF_n2788,
         dp_id_stage_regfile_DataPath_Physical_RF_n2787,
         dp_id_stage_regfile_DataPath_Physical_RF_n2786,
         dp_id_stage_regfile_DataPath_Physical_RF_n2785,
         dp_id_stage_regfile_DataPath_Physical_RF_n2784,
         dp_id_stage_regfile_DataPath_Physical_RF_n2783,
         dp_id_stage_regfile_DataPath_Physical_RF_n2782,
         dp_id_stage_regfile_DataPath_Physical_RF_n2781,
         dp_id_stage_regfile_DataPath_Physical_RF_n2780,
         dp_id_stage_regfile_DataPath_Physical_RF_n2779,
         dp_id_stage_regfile_DataPath_Physical_RF_n2778,
         dp_id_stage_regfile_DataPath_Physical_RF_n2777,
         dp_id_stage_regfile_DataPath_Physical_RF_n2776,
         dp_id_stage_regfile_DataPath_Physical_RF_n2775,
         dp_id_stage_regfile_DataPath_Physical_RF_n2774,
         dp_id_stage_regfile_DataPath_Physical_RF_n2773,
         dp_id_stage_regfile_DataPath_Physical_RF_n2772,
         dp_id_stage_regfile_DataPath_Physical_RF_n2771,
         dp_id_stage_regfile_DataPath_Physical_RF_n2770,
         dp_id_stage_regfile_DataPath_Physical_RF_n2769,
         dp_id_stage_regfile_DataPath_Physical_RF_n2768,
         dp_id_stage_regfile_DataPath_Physical_RF_n2767,
         dp_id_stage_regfile_DataPath_Physical_RF_n2766,
         dp_id_stage_regfile_DataPath_Physical_RF_n2765,
         dp_id_stage_regfile_DataPath_Physical_RF_n2764,
         dp_id_stage_regfile_DataPath_Physical_RF_n2763,
         dp_id_stage_regfile_DataPath_Physical_RF_n2762,
         dp_id_stage_regfile_DataPath_Physical_RF_n2761,
         dp_id_stage_regfile_DataPath_Physical_RF_n2760,
         dp_id_stage_regfile_DataPath_Physical_RF_n2759,
         dp_id_stage_regfile_DataPath_Physical_RF_n2758,
         dp_id_stage_regfile_DataPath_Physical_RF_n2757,
         dp_id_stage_regfile_DataPath_Physical_RF_n2756,
         dp_id_stage_regfile_DataPath_Physical_RF_n2755,
         dp_id_stage_regfile_DataPath_Physical_RF_n2754,
         dp_id_stage_regfile_DataPath_Physical_RF_n2753,
         dp_id_stage_regfile_DataPath_Physical_RF_n2752,
         dp_id_stage_regfile_DataPath_Physical_RF_n2751,
         dp_id_stage_regfile_DataPath_Physical_RF_n2750,
         dp_id_stage_regfile_DataPath_Physical_RF_n2749,
         dp_id_stage_regfile_DataPath_Physical_RF_n2748,
         dp_id_stage_regfile_DataPath_Physical_RF_n2747,
         dp_id_stage_regfile_DataPath_Physical_RF_n2746,
         dp_id_stage_regfile_DataPath_Physical_RF_n2745,
         dp_id_stage_regfile_DataPath_Physical_RF_n2744,
         dp_id_stage_regfile_DataPath_Physical_RF_n2743,
         dp_id_stage_regfile_DataPath_Physical_RF_n2742,
         dp_id_stage_regfile_DataPath_Physical_RF_n2741,
         dp_id_stage_regfile_DataPath_Physical_RF_n2740,
         dp_id_stage_regfile_DataPath_Physical_RF_n2739,
         dp_id_stage_regfile_DataPath_Physical_RF_n2738,
         dp_id_stage_regfile_DataPath_Physical_RF_n2737,
         dp_id_stage_regfile_DataPath_Physical_RF_n2736,
         dp_id_stage_regfile_DataPath_Physical_RF_n2735,
         dp_id_stage_regfile_DataPath_Physical_RF_n2734,
         dp_id_stage_regfile_DataPath_Physical_RF_n2733,
         dp_id_stage_regfile_DataPath_Physical_RF_n2732,
         dp_id_stage_regfile_DataPath_Physical_RF_n2731,
         dp_id_stage_regfile_DataPath_Physical_RF_n2730,
         dp_id_stage_regfile_DataPath_Physical_RF_n2729,
         dp_id_stage_regfile_DataPath_Physical_RF_n2728,
         dp_id_stage_regfile_DataPath_Physical_RF_n2727,
         dp_id_stage_regfile_DataPath_Physical_RF_n2726,
         dp_id_stage_regfile_DataPath_Physical_RF_n2725,
         dp_id_stage_regfile_DataPath_Physical_RF_n2724,
         dp_id_stage_regfile_DataPath_Physical_RF_n2723,
         dp_id_stage_regfile_DataPath_Physical_RF_n2722,
         dp_id_stage_regfile_DataPath_Physical_RF_n2721,
         dp_id_stage_regfile_DataPath_Physical_RF_n2720,
         dp_id_stage_regfile_DataPath_Physical_RF_n2719,
         dp_id_stage_regfile_DataPath_Physical_RF_n2718,
         dp_id_stage_regfile_DataPath_Physical_RF_n2717,
         dp_id_stage_regfile_DataPath_Physical_RF_n2716,
         dp_id_stage_regfile_DataPath_Physical_RF_n2715,
         dp_id_stage_regfile_DataPath_Physical_RF_n2714,
         dp_id_stage_regfile_DataPath_Physical_RF_n2713,
         dp_id_stage_regfile_DataPath_Physical_RF_n2712,
         dp_id_stage_regfile_DataPath_Physical_RF_n2711,
         dp_id_stage_regfile_DataPath_Physical_RF_n2710,
         dp_id_stage_regfile_DataPath_Physical_RF_n2709,
         dp_id_stage_regfile_DataPath_Physical_RF_n2708,
         dp_id_stage_regfile_DataPath_Physical_RF_n2707,
         dp_id_stage_regfile_DataPath_Physical_RF_n2706,
         dp_id_stage_regfile_DataPath_Physical_RF_n2705,
         dp_id_stage_regfile_DataPath_Physical_RF_n2704,
         dp_id_stage_regfile_DataPath_Physical_RF_n2703,
         dp_id_stage_regfile_DataPath_Physical_RF_n2702,
         dp_id_stage_regfile_DataPath_Physical_RF_n2701,
         dp_id_stage_regfile_DataPath_Physical_RF_n2700,
         dp_id_stage_regfile_DataPath_Physical_RF_n2699,
         dp_id_stage_regfile_DataPath_Physical_RF_n2698,
         dp_id_stage_regfile_DataPath_Physical_RF_n2697,
         dp_id_stage_regfile_DataPath_Physical_RF_n2696,
         dp_id_stage_regfile_DataPath_Physical_RF_n2695,
         dp_id_stage_regfile_DataPath_Physical_RF_n2694,
         dp_id_stage_regfile_DataPath_Physical_RF_n2693,
         dp_id_stage_regfile_DataPath_Physical_RF_n2692,
         dp_id_stage_regfile_DataPath_Physical_RF_n2691,
         dp_id_stage_regfile_DataPath_Physical_RF_n2690,
         dp_id_stage_regfile_DataPath_Physical_RF_n2689,
         dp_id_stage_regfile_DataPath_Physical_RF_n2688,
         dp_id_stage_regfile_DataPath_Physical_RF_n2687,
         dp_id_stage_regfile_DataPath_Physical_RF_n2686,
         dp_id_stage_regfile_DataPath_Physical_RF_n2685,
         dp_id_stage_regfile_DataPath_Physical_RF_n2684,
         dp_id_stage_regfile_DataPath_Physical_RF_n2683,
         dp_id_stage_regfile_DataPath_Physical_RF_n2682,
         dp_id_stage_regfile_DataPath_Physical_RF_n2681,
         dp_id_stage_regfile_DataPath_Physical_RF_n2680,
         dp_id_stage_regfile_DataPath_Physical_RF_n2679,
         dp_id_stage_regfile_DataPath_Physical_RF_n2678,
         dp_id_stage_regfile_DataPath_Physical_RF_n2677,
         dp_id_stage_regfile_DataPath_Physical_RF_n2676,
         dp_id_stage_regfile_DataPath_Physical_RF_n2675,
         dp_id_stage_regfile_DataPath_Physical_RF_n2674,
         dp_id_stage_regfile_DataPath_Physical_RF_n2673,
         dp_id_stage_regfile_DataPath_Physical_RF_n2672,
         dp_id_stage_regfile_DataPath_Physical_RF_n2671,
         dp_id_stage_regfile_DataPath_Physical_RF_n2670,
         dp_id_stage_regfile_DataPath_Physical_RF_n2669,
         dp_id_stage_regfile_DataPath_Physical_RF_n2668,
         dp_id_stage_regfile_DataPath_Physical_RF_n2667,
         dp_id_stage_regfile_DataPath_Physical_RF_n2666,
         dp_id_stage_regfile_DataPath_Physical_RF_n2665,
         dp_id_stage_regfile_DataPath_Physical_RF_n2664,
         dp_id_stage_regfile_DataPath_Physical_RF_n2663,
         dp_id_stage_regfile_DataPath_Physical_RF_n2662,
         dp_id_stage_regfile_DataPath_Physical_RF_n2661,
         dp_id_stage_regfile_DataPath_Physical_RF_n2660,
         dp_id_stage_regfile_DataPath_Physical_RF_n2659,
         dp_id_stage_regfile_DataPath_Physical_RF_n2658,
         dp_id_stage_regfile_DataPath_Physical_RF_n2657,
         dp_id_stage_regfile_DataPath_Physical_RF_n2656,
         dp_id_stage_regfile_DataPath_Physical_RF_n2655,
         dp_id_stage_regfile_DataPath_Physical_RF_n2654,
         dp_id_stage_regfile_DataPath_Physical_RF_n2653,
         dp_id_stage_regfile_DataPath_Physical_RF_n2652,
         dp_id_stage_regfile_DataPath_Physical_RF_n2651,
         dp_id_stage_regfile_DataPath_Physical_RF_n2650,
         dp_id_stage_regfile_DataPath_Physical_RF_n2649,
         dp_id_stage_regfile_DataPath_Physical_RF_n2648,
         dp_id_stage_regfile_DataPath_Physical_RF_n2647,
         dp_id_stage_regfile_DataPath_Physical_RF_n2646,
         dp_id_stage_regfile_DataPath_Physical_RF_n2645,
         dp_id_stage_regfile_DataPath_Physical_RF_n2644,
         dp_id_stage_regfile_DataPath_Physical_RF_n2643,
         dp_id_stage_regfile_DataPath_Physical_RF_n2642,
         dp_id_stage_regfile_DataPath_Physical_RF_n2641,
         dp_id_stage_regfile_DataPath_Physical_RF_n2640,
         dp_id_stage_regfile_DataPath_Physical_RF_n2639,
         dp_id_stage_regfile_DataPath_Physical_RF_n2638,
         dp_id_stage_regfile_DataPath_Physical_RF_n2637,
         dp_id_stage_regfile_DataPath_Physical_RF_n2636,
         dp_id_stage_regfile_DataPath_Physical_RF_n2635,
         dp_id_stage_regfile_DataPath_Physical_RF_n2634,
         dp_id_stage_regfile_DataPath_Physical_RF_n2633,
         dp_id_stage_regfile_DataPath_Physical_RF_n2632,
         dp_id_stage_regfile_DataPath_Physical_RF_n2631,
         dp_id_stage_regfile_DataPath_Physical_RF_n2630,
         dp_id_stage_regfile_DataPath_Physical_RF_n2629,
         dp_id_stage_regfile_DataPath_Physical_RF_n2628,
         dp_id_stage_regfile_DataPath_Physical_RF_n2627,
         dp_id_stage_regfile_DataPath_Physical_RF_n2626,
         dp_id_stage_regfile_DataPath_Physical_RF_n2625,
         dp_id_stage_regfile_DataPath_Physical_RF_n2624,
         dp_id_stage_regfile_DataPath_Physical_RF_n2623,
         dp_id_stage_regfile_DataPath_Physical_RF_n2622,
         dp_id_stage_regfile_DataPath_Physical_RF_n2621,
         dp_id_stage_regfile_DataPath_Physical_RF_n2620,
         dp_id_stage_regfile_DataPath_Physical_RF_n2619,
         dp_id_stage_regfile_DataPath_Physical_RF_n2618,
         dp_id_stage_regfile_DataPath_Physical_RF_n2617,
         dp_id_stage_regfile_DataPath_Physical_RF_n2616,
         dp_id_stage_regfile_DataPath_Physical_RF_n2615,
         dp_id_stage_regfile_DataPath_Physical_RF_n2614,
         dp_id_stage_regfile_DataPath_Physical_RF_n2613,
         dp_id_stage_regfile_DataPath_Physical_RF_n2612,
         dp_id_stage_regfile_DataPath_Physical_RF_n2611,
         dp_id_stage_regfile_DataPath_Physical_RF_n2610,
         dp_id_stage_regfile_DataPath_Physical_RF_n2609,
         dp_id_stage_regfile_DataPath_Physical_RF_n2608,
         dp_id_stage_regfile_DataPath_Physical_RF_n2607,
         dp_id_stage_regfile_DataPath_Physical_RF_n2606,
         dp_id_stage_regfile_DataPath_Physical_RF_n2605,
         dp_id_stage_regfile_DataPath_Physical_RF_n2604,
         dp_id_stage_regfile_DataPath_Physical_RF_n2603,
         dp_id_stage_regfile_DataPath_Physical_RF_n2602,
         dp_id_stage_regfile_DataPath_Physical_RF_n2601,
         dp_id_stage_regfile_DataPath_Physical_RF_n2600,
         dp_id_stage_regfile_DataPath_Physical_RF_n2599,
         dp_id_stage_regfile_DataPath_Physical_RF_n2598,
         dp_id_stage_regfile_DataPath_Physical_RF_n2597,
         dp_id_stage_regfile_DataPath_Physical_RF_n2596,
         dp_id_stage_regfile_DataPath_Physical_RF_n2595,
         dp_id_stage_regfile_DataPath_Physical_RF_n2594,
         dp_id_stage_regfile_DataPath_Physical_RF_n2593,
         dp_id_stage_regfile_DataPath_Physical_RF_n2592,
         dp_id_stage_regfile_DataPath_Physical_RF_n2591,
         dp_id_stage_regfile_DataPath_Physical_RF_n2590,
         dp_id_stage_regfile_DataPath_Physical_RF_n2589,
         dp_id_stage_regfile_DataPath_Physical_RF_n2588,
         dp_id_stage_regfile_DataPath_Physical_RF_n2587,
         dp_id_stage_regfile_DataPath_Physical_RF_n2586,
         dp_id_stage_regfile_DataPath_Physical_RF_n2585,
         dp_id_stage_regfile_DataPath_Physical_RF_n2584,
         dp_id_stage_regfile_DataPath_Physical_RF_n2583,
         dp_id_stage_regfile_DataPath_Physical_RF_n2582,
         dp_id_stage_regfile_DataPath_Physical_RF_n2581,
         dp_id_stage_regfile_DataPath_Physical_RF_n2580,
         dp_id_stage_regfile_DataPath_Physical_RF_n2579,
         dp_id_stage_regfile_DataPath_Physical_RF_n2578,
         dp_id_stage_regfile_DataPath_Physical_RF_n2577,
         dp_id_stage_regfile_DataPath_Physical_RF_n2576,
         dp_id_stage_regfile_DataPath_Physical_RF_n2575,
         dp_id_stage_regfile_DataPath_Physical_RF_n2574,
         dp_id_stage_regfile_DataPath_Physical_RF_n2573,
         dp_id_stage_regfile_DataPath_Physical_RF_n2572,
         dp_id_stage_regfile_DataPath_Physical_RF_n2571,
         dp_id_stage_regfile_DataPath_Physical_RF_n2570,
         dp_id_stage_regfile_DataPath_Physical_RF_n2569,
         dp_id_stage_regfile_DataPath_Physical_RF_n2568,
         dp_id_stage_regfile_DataPath_Physical_RF_n2567,
         dp_id_stage_regfile_DataPath_Physical_RF_n2566,
         dp_id_stage_regfile_DataPath_Physical_RF_n2565,
         dp_id_stage_regfile_DataPath_Physical_RF_n2564,
         dp_id_stage_regfile_DataPath_Physical_RF_n2563,
         dp_id_stage_regfile_DataPath_Physical_RF_n2562,
         dp_id_stage_regfile_DataPath_Physical_RF_n2561,
         dp_id_stage_regfile_DataPath_Physical_RF_n2560,
         dp_id_stage_regfile_DataPath_Physical_RF_n2559,
         dp_id_stage_regfile_DataPath_Physical_RF_n2558,
         dp_id_stage_regfile_DataPath_Physical_RF_n2557,
         dp_id_stage_regfile_DataPath_Physical_RF_n2556,
         dp_id_stage_regfile_DataPath_Physical_RF_n2555,
         dp_id_stage_regfile_DataPath_Physical_RF_n2554,
         dp_id_stage_regfile_DataPath_Physical_RF_n2553,
         dp_id_stage_regfile_DataPath_Physical_RF_n2552,
         dp_id_stage_regfile_DataPath_Physical_RF_n2551,
         dp_id_stage_regfile_DataPath_Physical_RF_n2550,
         dp_id_stage_regfile_DataPath_Physical_RF_n2549,
         dp_id_stage_regfile_DataPath_Physical_RF_n2548,
         dp_id_stage_regfile_DataPath_Physical_RF_n2547,
         dp_id_stage_regfile_DataPath_Physical_RF_n2546,
         dp_id_stage_regfile_DataPath_Physical_RF_n2545,
         dp_id_stage_regfile_DataPath_Physical_RF_n2544,
         dp_id_stage_regfile_DataPath_Physical_RF_n2543,
         dp_id_stage_regfile_DataPath_Physical_RF_n2542,
         dp_id_stage_regfile_DataPath_Physical_RF_n2541,
         dp_id_stage_regfile_DataPath_Physical_RF_n2540,
         dp_id_stage_regfile_DataPath_Physical_RF_n2539,
         dp_id_stage_regfile_DataPath_Physical_RF_n2538,
         dp_id_stage_regfile_DataPath_Physical_RF_n2537,
         dp_id_stage_regfile_DataPath_Physical_RF_n2536,
         dp_id_stage_regfile_DataPath_Physical_RF_n2535,
         dp_id_stage_regfile_DataPath_Physical_RF_n2534,
         dp_id_stage_regfile_DataPath_Physical_RF_n2533,
         dp_id_stage_regfile_DataPath_Physical_RF_n2532,
         dp_id_stage_regfile_DataPath_Physical_RF_n2531,
         dp_id_stage_regfile_DataPath_Physical_RF_n2530,
         dp_id_stage_regfile_DataPath_Physical_RF_n2529,
         dp_id_stage_regfile_DataPath_Physical_RF_n2528,
         dp_id_stage_regfile_DataPath_Physical_RF_n2527,
         dp_id_stage_regfile_DataPath_Physical_RF_n2526,
         dp_id_stage_regfile_DataPath_Physical_RF_n2525,
         dp_id_stage_regfile_DataPath_Physical_RF_n2524,
         dp_id_stage_regfile_DataPath_Physical_RF_n2523,
         dp_id_stage_regfile_DataPath_Physical_RF_n2522,
         dp_id_stage_regfile_DataPath_Physical_RF_n2521,
         dp_id_stage_regfile_DataPath_Physical_RF_n2520,
         dp_id_stage_regfile_DataPath_Physical_RF_n2519,
         dp_id_stage_regfile_DataPath_Physical_RF_n2518,
         dp_id_stage_regfile_DataPath_Physical_RF_n2517,
         dp_id_stage_regfile_DataPath_Physical_RF_n2516,
         dp_id_stage_regfile_DataPath_Physical_RF_n2515,
         dp_id_stage_regfile_DataPath_Physical_RF_n2514,
         dp_id_stage_regfile_DataPath_Physical_RF_n2513,
         dp_id_stage_regfile_DataPath_Physical_RF_n2512,
         dp_id_stage_regfile_DataPath_Physical_RF_n2511,
         dp_id_stage_regfile_DataPath_Physical_RF_n2510,
         dp_id_stage_regfile_DataPath_Physical_RF_n2509,
         dp_id_stage_regfile_DataPath_Physical_RF_n2508,
         dp_id_stage_regfile_DataPath_Physical_RF_n2507,
         dp_id_stage_regfile_DataPath_Physical_RF_n2506,
         dp_id_stage_regfile_DataPath_Physical_RF_n2505,
         dp_id_stage_regfile_DataPath_Physical_RF_n2504,
         dp_id_stage_regfile_DataPath_Physical_RF_n2503,
         dp_id_stage_regfile_DataPath_Physical_RF_n2502,
         dp_id_stage_regfile_DataPath_Physical_RF_n2501,
         dp_id_stage_regfile_DataPath_Physical_RF_n2500,
         dp_id_stage_regfile_DataPath_Physical_RF_n2499,
         dp_id_stage_regfile_DataPath_Physical_RF_n2498,
         dp_id_stage_regfile_DataPath_Physical_RF_n2497,
         dp_id_stage_regfile_DataPath_Physical_RF_n2496,
         dp_id_stage_regfile_DataPath_Physical_RF_n2495,
         dp_id_stage_regfile_DataPath_Physical_RF_n2494,
         dp_id_stage_regfile_DataPath_Physical_RF_n2493,
         dp_id_stage_regfile_DataPath_Physical_RF_n2492,
         dp_id_stage_regfile_DataPath_Physical_RF_n2491,
         dp_id_stage_regfile_DataPath_Physical_RF_n2490,
         dp_id_stage_regfile_DataPath_Physical_RF_n2489,
         dp_id_stage_regfile_DataPath_Physical_RF_n2488,
         dp_id_stage_regfile_DataPath_Physical_RF_n2487,
         dp_id_stage_regfile_DataPath_Physical_RF_n2486,
         dp_id_stage_regfile_DataPath_Physical_RF_n2485,
         dp_id_stage_regfile_DataPath_Physical_RF_n2484,
         dp_id_stage_regfile_DataPath_Physical_RF_n2483,
         dp_id_stage_regfile_DataPath_Physical_RF_n2482,
         dp_id_stage_regfile_DataPath_Physical_RF_n2481,
         dp_id_stage_regfile_DataPath_Physical_RF_n2480,
         dp_id_stage_regfile_DataPath_Physical_RF_n2479,
         dp_id_stage_regfile_DataPath_Physical_RF_n2478,
         dp_id_stage_regfile_DataPath_Physical_RF_n2477,
         dp_id_stage_regfile_DataPath_Physical_RF_n2476,
         dp_id_stage_regfile_DataPath_Physical_RF_n2475,
         dp_id_stage_regfile_DataPath_Physical_RF_n2474,
         dp_id_stage_regfile_DataPath_Physical_RF_n2473,
         dp_id_stage_regfile_DataPath_Physical_RF_n2472,
         dp_id_stage_regfile_DataPath_Physical_RF_n2471,
         dp_id_stage_regfile_DataPath_Physical_RF_n2470,
         dp_id_stage_regfile_DataPath_Physical_RF_n2469,
         dp_id_stage_regfile_DataPath_Physical_RF_n2468,
         dp_id_stage_regfile_DataPath_Physical_RF_n2467,
         dp_id_stage_regfile_DataPath_Physical_RF_n2466,
         dp_id_stage_regfile_DataPath_Physical_RF_n2465,
         dp_id_stage_regfile_DataPath_Physical_RF_n2464,
         dp_id_stage_regfile_DataPath_Physical_RF_n2463,
         dp_id_stage_regfile_DataPath_Physical_RF_n2462,
         dp_id_stage_regfile_DataPath_Physical_RF_n2461,
         dp_id_stage_regfile_DataPath_Physical_RF_n2460,
         dp_id_stage_regfile_DataPath_Physical_RF_n2459,
         dp_id_stage_regfile_DataPath_Physical_RF_n2458,
         dp_id_stage_regfile_DataPath_Physical_RF_n2457,
         dp_id_stage_regfile_DataPath_Physical_RF_n2456,
         dp_id_stage_regfile_DataPath_Physical_RF_n2455,
         dp_id_stage_regfile_DataPath_Physical_RF_n2454,
         dp_id_stage_regfile_DataPath_Physical_RF_n2453,
         dp_id_stage_regfile_DataPath_Physical_RF_n2452,
         dp_id_stage_regfile_DataPath_Physical_RF_n2451,
         dp_id_stage_regfile_DataPath_Physical_RF_n2450,
         dp_id_stage_regfile_DataPath_Physical_RF_n2449,
         dp_id_stage_regfile_DataPath_Physical_RF_n2448,
         dp_id_stage_regfile_DataPath_Physical_RF_n2447,
         dp_id_stage_regfile_DataPath_Physical_RF_n2446,
         dp_id_stage_regfile_DataPath_Physical_RF_n2445,
         dp_id_stage_regfile_DataPath_Physical_RF_n2444,
         dp_id_stage_regfile_DataPath_Physical_RF_n2443,
         dp_id_stage_regfile_DataPath_Physical_RF_n2442,
         dp_id_stage_regfile_DataPath_Physical_RF_n2441,
         dp_id_stage_regfile_DataPath_Physical_RF_n2440,
         dp_id_stage_regfile_DataPath_Physical_RF_n2439,
         dp_id_stage_regfile_DataPath_Physical_RF_n2438,
         dp_id_stage_regfile_DataPath_Physical_RF_n2437,
         dp_id_stage_regfile_DataPath_Physical_RF_n2436,
         dp_id_stage_regfile_DataPath_Physical_RF_n2435,
         dp_id_stage_regfile_DataPath_Physical_RF_n2434,
         dp_id_stage_regfile_DataPath_Physical_RF_n2433,
         dp_id_stage_regfile_DataPath_Physical_RF_n2432,
         dp_id_stage_regfile_DataPath_Physical_RF_n2431,
         dp_id_stage_regfile_DataPath_Physical_RF_n2430,
         dp_id_stage_regfile_DataPath_Physical_RF_n2429,
         dp_id_stage_regfile_DataPath_Physical_RF_n2428,
         dp_id_stage_regfile_DataPath_Physical_RF_n2427,
         dp_id_stage_regfile_DataPath_Physical_RF_n2426,
         dp_id_stage_regfile_DataPath_Physical_RF_n2425,
         dp_id_stage_regfile_DataPath_Physical_RF_n2424,
         dp_id_stage_regfile_DataPath_Physical_RF_n2423,
         dp_id_stage_regfile_DataPath_Physical_RF_n2422,
         dp_id_stage_regfile_DataPath_Physical_RF_n2421,
         dp_id_stage_regfile_DataPath_Physical_RF_n2420,
         dp_id_stage_regfile_DataPath_Physical_RF_n2419,
         dp_id_stage_regfile_DataPath_Physical_RF_n2418,
         dp_id_stage_regfile_DataPath_Physical_RF_n2417,
         dp_id_stage_regfile_DataPath_Physical_RF_n2416,
         dp_id_stage_regfile_DataPath_Physical_RF_n2415,
         dp_id_stage_regfile_DataPath_Physical_RF_n2414,
         dp_id_stage_regfile_DataPath_Physical_RF_n2413,
         dp_id_stage_regfile_DataPath_Physical_RF_n2412,
         dp_id_stage_regfile_DataPath_Physical_RF_n2411,
         dp_id_stage_regfile_DataPath_Physical_RF_n2410,
         dp_id_stage_regfile_DataPath_Physical_RF_n2409,
         dp_id_stage_regfile_DataPath_Physical_RF_n2408,
         dp_id_stage_regfile_DataPath_Physical_RF_n2407,
         dp_id_stage_regfile_DataPath_Physical_RF_n2406,
         dp_id_stage_regfile_DataPath_Physical_RF_n2405,
         dp_id_stage_regfile_DataPath_Physical_RF_n2404,
         dp_id_stage_regfile_DataPath_Physical_RF_n2403,
         dp_id_stage_regfile_DataPath_Physical_RF_n2402,
         dp_id_stage_regfile_DataPath_Physical_RF_n2401,
         dp_id_stage_regfile_DataPath_Physical_RF_n2400,
         dp_id_stage_regfile_DataPath_Physical_RF_n2399,
         dp_id_stage_regfile_DataPath_Physical_RF_n2398,
         dp_id_stage_regfile_DataPath_Physical_RF_n2397,
         dp_id_stage_regfile_DataPath_Physical_RF_n2396,
         dp_id_stage_regfile_DataPath_Physical_RF_n2395,
         dp_id_stage_regfile_DataPath_Physical_RF_n2394,
         dp_id_stage_regfile_DataPath_Physical_RF_n2393,
         dp_id_stage_regfile_DataPath_Physical_RF_n2392,
         dp_id_stage_regfile_DataPath_Physical_RF_n2391,
         dp_id_stage_regfile_DataPath_Physical_RF_n2390,
         dp_id_stage_regfile_DataPath_Physical_RF_n2389,
         dp_id_stage_regfile_DataPath_Physical_RF_n2388,
         dp_id_stage_regfile_DataPath_Physical_RF_n2387,
         dp_id_stage_regfile_DataPath_Physical_RF_n2386,
         dp_id_stage_regfile_DataPath_Physical_RF_n2385,
         dp_id_stage_regfile_DataPath_Physical_RF_n2384,
         dp_id_stage_regfile_DataPath_Physical_RF_n2383,
         dp_id_stage_regfile_DataPath_Physical_RF_n2382,
         dp_id_stage_regfile_DataPath_Physical_RF_n2381,
         dp_id_stage_regfile_DataPath_Physical_RF_n2380,
         dp_id_stage_regfile_DataPath_Physical_RF_n2379,
         dp_id_stage_regfile_DataPath_Physical_RF_n2378,
         dp_id_stage_regfile_DataPath_Physical_RF_n2377,
         dp_id_stage_regfile_DataPath_Physical_RF_n2376,
         dp_id_stage_regfile_DataPath_Physical_RF_n2375,
         dp_id_stage_regfile_DataPath_Physical_RF_n2374,
         dp_id_stage_regfile_DataPath_Physical_RF_n2373,
         dp_id_stage_regfile_DataPath_Physical_RF_n2372,
         dp_id_stage_regfile_DataPath_Physical_RF_n2371,
         dp_id_stage_regfile_DataPath_Physical_RF_n2370,
         dp_id_stage_regfile_DataPath_Physical_RF_n2369,
         dp_id_stage_regfile_DataPath_Physical_RF_n2368,
         dp_id_stage_regfile_DataPath_Physical_RF_n2367,
         dp_id_stage_regfile_DataPath_Physical_RF_n2366,
         dp_id_stage_regfile_DataPath_Physical_RF_n2365,
         dp_id_stage_regfile_DataPath_Physical_RF_n2364,
         dp_id_stage_regfile_DataPath_Physical_RF_n2363,
         dp_id_stage_regfile_DataPath_Physical_RF_n2362,
         dp_id_stage_regfile_DataPath_Physical_RF_n2361,
         dp_id_stage_regfile_DataPath_Physical_RF_n2360,
         dp_id_stage_regfile_DataPath_Physical_RF_n2359,
         dp_id_stage_regfile_DataPath_Physical_RF_n2358,
         dp_id_stage_regfile_DataPath_Physical_RF_n2357,
         dp_id_stage_regfile_DataPath_Physical_RF_n2356,
         dp_id_stage_regfile_DataPath_Physical_RF_n2355,
         dp_id_stage_regfile_DataPath_Physical_RF_n2354,
         dp_id_stage_regfile_DataPath_Physical_RF_n2353,
         dp_id_stage_regfile_DataPath_Physical_RF_n2352,
         dp_id_stage_regfile_DataPath_Physical_RF_n2351,
         dp_id_stage_regfile_DataPath_Physical_RF_n2350,
         dp_id_stage_regfile_DataPath_Physical_RF_n2349,
         dp_id_stage_regfile_DataPath_Physical_RF_n2348,
         dp_id_stage_regfile_DataPath_Physical_RF_n2347,
         dp_id_stage_regfile_DataPath_Physical_RF_n2346,
         dp_id_stage_regfile_DataPath_Physical_RF_n2345,
         dp_id_stage_regfile_DataPath_Physical_RF_n2344,
         dp_id_stage_regfile_DataPath_Physical_RF_n2343,
         dp_id_stage_regfile_DataPath_Physical_RF_n2342,
         dp_id_stage_regfile_DataPath_Physical_RF_n2341,
         dp_id_stage_regfile_DataPath_Physical_RF_n2340,
         dp_id_stage_regfile_DataPath_Physical_RF_n2339,
         dp_id_stage_regfile_DataPath_Physical_RF_n2338,
         dp_id_stage_regfile_DataPath_Physical_RF_n2337,
         dp_id_stage_regfile_DataPath_Physical_RF_n2336,
         dp_id_stage_regfile_DataPath_Physical_RF_n2335,
         dp_id_stage_regfile_DataPath_Physical_RF_n2334,
         dp_id_stage_regfile_DataPath_Physical_RF_n2333,
         dp_id_stage_regfile_DataPath_Physical_RF_n2332,
         dp_id_stage_regfile_DataPath_Physical_RF_n2331,
         dp_id_stage_regfile_DataPath_Physical_RF_n2330,
         dp_id_stage_regfile_DataPath_Physical_RF_n2329,
         dp_id_stage_regfile_DataPath_Physical_RF_n2328,
         dp_id_stage_regfile_DataPath_Physical_RF_n2327,
         dp_id_stage_regfile_DataPath_Physical_RF_n2326,
         dp_id_stage_regfile_DataPath_Physical_RF_n2325,
         dp_id_stage_regfile_DataPath_Physical_RF_n2324,
         dp_id_stage_regfile_DataPath_Physical_RF_n2323,
         dp_id_stage_regfile_DataPath_Physical_RF_n2322,
         dp_id_stage_regfile_DataPath_Physical_RF_n2321,
         dp_id_stage_regfile_DataPath_Physical_RF_n2320,
         dp_id_stage_regfile_DataPath_Physical_RF_n2319,
         dp_id_stage_regfile_DataPath_Physical_RF_n2318,
         dp_id_stage_regfile_DataPath_Physical_RF_n2317,
         dp_id_stage_regfile_DataPath_Physical_RF_n2316,
         dp_id_stage_regfile_DataPath_Physical_RF_n2315,
         dp_id_stage_regfile_DataPath_Physical_RF_n2314,
         dp_id_stage_regfile_DataPath_Physical_RF_n2313,
         dp_id_stage_regfile_DataPath_Physical_RF_n2312,
         dp_id_stage_regfile_DataPath_Physical_RF_n2311,
         dp_id_stage_regfile_DataPath_Physical_RF_n2310,
         dp_id_stage_regfile_DataPath_Physical_RF_n2309,
         dp_id_stage_regfile_DataPath_Physical_RF_n2308,
         dp_id_stage_regfile_DataPath_Physical_RF_n2307,
         dp_id_stage_regfile_DataPath_Physical_RF_n2306,
         dp_id_stage_regfile_DataPath_Physical_RF_n2305,
         dp_id_stage_regfile_DataPath_Physical_RF_n2304,
         dp_id_stage_regfile_DataPath_Physical_RF_n2303,
         dp_id_stage_regfile_DataPath_Physical_RF_n2302,
         dp_id_stage_regfile_DataPath_Physical_RF_n2301,
         dp_id_stage_regfile_DataPath_Physical_RF_n2300,
         dp_id_stage_regfile_DataPath_Physical_RF_n2299,
         dp_id_stage_regfile_DataPath_Physical_RF_n2298,
         dp_id_stage_regfile_DataPath_Physical_RF_n2297,
         dp_id_stage_regfile_DataPath_Physical_RF_n2296,
         dp_id_stage_regfile_DataPath_Physical_RF_n2295,
         dp_id_stage_regfile_DataPath_Physical_RF_n2294,
         dp_id_stage_regfile_DataPath_Physical_RF_n2293,
         dp_id_stage_regfile_DataPath_Physical_RF_n2292,
         dp_id_stage_regfile_DataPath_Physical_RF_n2291,
         dp_id_stage_regfile_DataPath_Physical_RF_n2290,
         dp_id_stage_regfile_DataPath_Physical_RF_n2289,
         dp_id_stage_regfile_DataPath_Physical_RF_n2288,
         dp_id_stage_regfile_DataPath_Physical_RF_n2287,
         dp_id_stage_regfile_DataPath_Physical_RF_n2286,
         dp_id_stage_regfile_DataPath_Physical_RF_n2285,
         dp_id_stage_regfile_DataPath_Physical_RF_n2284,
         dp_id_stage_regfile_DataPath_Physical_RF_n2283,
         dp_id_stage_regfile_DataPath_Physical_RF_n2282,
         dp_id_stage_regfile_DataPath_Physical_RF_n2281,
         dp_id_stage_regfile_DataPath_Physical_RF_n2280,
         dp_id_stage_regfile_DataPath_Physical_RF_n2279,
         dp_id_stage_regfile_DataPath_Physical_RF_n2278,
         dp_id_stage_regfile_DataPath_Physical_RF_n2277,
         dp_id_stage_regfile_DataPath_Physical_RF_n2276,
         dp_id_stage_regfile_DataPath_Physical_RF_n2275,
         dp_id_stage_regfile_DataPath_Physical_RF_n2274,
         dp_id_stage_regfile_DataPath_Physical_RF_n2273,
         dp_id_stage_regfile_DataPath_Physical_RF_n2272,
         dp_id_stage_regfile_DataPath_Physical_RF_n2271,
         dp_id_stage_regfile_DataPath_Physical_RF_n2270,
         dp_id_stage_regfile_DataPath_Physical_RF_n2269,
         dp_id_stage_regfile_DataPath_Physical_RF_n2268,
         dp_id_stage_regfile_DataPath_Physical_RF_n2267,
         dp_id_stage_regfile_DataPath_Physical_RF_n2266,
         dp_id_stage_regfile_DataPath_Physical_RF_n2265,
         dp_id_stage_regfile_DataPath_Physical_RF_n2264,
         dp_id_stage_regfile_DataPath_Physical_RF_n2263,
         dp_id_stage_regfile_DataPath_Physical_RF_n2262,
         dp_id_stage_regfile_DataPath_Physical_RF_n2261,
         dp_id_stage_regfile_DataPath_Physical_RF_n2260,
         dp_id_stage_regfile_DataPath_Physical_RF_n2259,
         dp_id_stage_regfile_DataPath_Physical_RF_n2258,
         dp_id_stage_regfile_DataPath_Physical_RF_n2257,
         dp_id_stage_regfile_DataPath_Physical_RF_n2256,
         dp_id_stage_regfile_DataPath_Physical_RF_n2255,
         dp_id_stage_regfile_DataPath_Physical_RF_n2254,
         dp_id_stage_regfile_DataPath_Physical_RF_n2253,
         dp_id_stage_regfile_DataPath_Physical_RF_n2252,
         dp_id_stage_regfile_DataPath_Physical_RF_n2251,
         dp_id_stage_regfile_DataPath_Physical_RF_n2250,
         dp_id_stage_regfile_DataPath_Physical_RF_n2249,
         dp_id_stage_regfile_DataPath_Physical_RF_n2248,
         dp_id_stage_regfile_DataPath_Physical_RF_n2247,
         dp_id_stage_regfile_DataPath_Physical_RF_n2246,
         dp_id_stage_regfile_DataPath_Physical_RF_n2245,
         dp_id_stage_regfile_DataPath_Physical_RF_n2244,
         dp_id_stage_regfile_DataPath_Physical_RF_n2243,
         dp_id_stage_regfile_DataPath_Physical_RF_n2242,
         dp_id_stage_regfile_DataPath_Physical_RF_n2241,
         dp_id_stage_regfile_DataPath_Physical_RF_n2240,
         dp_id_stage_regfile_DataPath_Physical_RF_n2239,
         dp_id_stage_regfile_DataPath_Physical_RF_n2238,
         dp_id_stage_regfile_DataPath_Physical_RF_n2237,
         dp_id_stage_regfile_DataPath_Physical_RF_n2236,
         dp_id_stage_regfile_DataPath_Physical_RF_n2235,
         dp_id_stage_regfile_DataPath_Physical_RF_n2234,
         dp_id_stage_regfile_DataPath_Physical_RF_n2233,
         dp_id_stage_regfile_DataPath_Physical_RF_n2232,
         dp_id_stage_regfile_DataPath_Physical_RF_n2231,
         dp_id_stage_regfile_DataPath_Physical_RF_n2230,
         dp_id_stage_regfile_DataPath_Physical_RF_n2229,
         dp_id_stage_regfile_DataPath_Physical_RF_n2228,
         dp_id_stage_regfile_DataPath_Physical_RF_n2227,
         dp_id_stage_regfile_DataPath_Physical_RF_n2226,
         dp_id_stage_regfile_DataPath_Physical_RF_n2225,
         dp_id_stage_regfile_DataPath_Physical_RF_n2224,
         dp_id_stage_regfile_DataPath_Physical_RF_n2223,
         dp_id_stage_regfile_DataPath_Physical_RF_n2222,
         dp_id_stage_regfile_DataPath_Physical_RF_n2221,
         dp_id_stage_regfile_DataPath_Physical_RF_n2220,
         dp_id_stage_regfile_DataPath_Physical_RF_n2219,
         dp_id_stage_regfile_DataPath_Physical_RF_n2218,
         dp_id_stage_regfile_DataPath_Physical_RF_n2217,
         dp_id_stage_regfile_DataPath_Physical_RF_n2216,
         dp_id_stage_regfile_DataPath_Physical_RF_n2215,
         dp_id_stage_regfile_DataPath_Physical_RF_n2214,
         dp_id_stage_regfile_DataPath_Physical_RF_n2213,
         dp_id_stage_regfile_DataPath_Physical_RF_n2212,
         dp_id_stage_regfile_DataPath_Physical_RF_n2211,
         dp_id_stage_regfile_DataPath_Physical_RF_n2210,
         dp_id_stage_regfile_DataPath_Physical_RF_n2209,
         dp_id_stage_regfile_DataPath_Physical_RF_n2208,
         dp_id_stage_regfile_DataPath_Physical_RF_n2207,
         dp_id_stage_regfile_DataPath_Physical_RF_n2206,
         dp_id_stage_regfile_DataPath_Physical_RF_n2205,
         dp_id_stage_regfile_DataPath_Physical_RF_n2204,
         dp_id_stage_regfile_DataPath_Physical_RF_n2203,
         dp_id_stage_regfile_DataPath_Physical_RF_n2202,
         dp_id_stage_regfile_DataPath_Physical_RF_n2201,
         dp_id_stage_regfile_DataPath_Physical_RF_n2200,
         dp_id_stage_regfile_DataPath_Physical_RF_n2199,
         dp_id_stage_regfile_DataPath_Physical_RF_n2198,
         dp_id_stage_regfile_DataPath_Physical_RF_n2197,
         dp_id_stage_regfile_DataPath_Physical_RF_n2196,
         dp_id_stage_regfile_DataPath_Physical_RF_n2195,
         dp_id_stage_regfile_DataPath_Physical_RF_n2194,
         dp_id_stage_regfile_DataPath_Physical_RF_n2193,
         dp_id_stage_regfile_DataPath_Physical_RF_n2192,
         dp_id_stage_regfile_DataPath_Physical_RF_n2191,
         dp_id_stage_regfile_DataPath_Physical_RF_n2190,
         dp_id_stage_regfile_DataPath_Physical_RF_n2189,
         dp_id_stage_regfile_DataPath_Physical_RF_n2188,
         dp_id_stage_regfile_DataPath_Physical_RF_n2187,
         dp_id_stage_regfile_DataPath_Physical_RF_n2186,
         dp_id_stage_regfile_DataPath_Physical_RF_n2185,
         dp_id_stage_regfile_DataPath_Physical_RF_n2184,
         dp_id_stage_regfile_DataPath_Physical_RF_n2183,
         dp_id_stage_regfile_DataPath_Physical_RF_n2182,
         dp_id_stage_regfile_DataPath_Physical_RF_n2181,
         dp_id_stage_regfile_DataPath_Physical_RF_n2180,
         dp_id_stage_regfile_DataPath_Physical_RF_n2179,
         dp_id_stage_regfile_DataPath_Physical_RF_n2178,
         dp_id_stage_regfile_DataPath_Physical_RF_n2177,
         dp_id_stage_regfile_DataPath_Physical_RF_n2176,
         dp_id_stage_regfile_DataPath_Physical_RF_n2175,
         dp_id_stage_regfile_DataPath_Physical_RF_n2174,
         dp_id_stage_regfile_DataPath_Physical_RF_n2173,
         dp_id_stage_regfile_DataPath_Physical_RF_n2172,
         dp_id_stage_regfile_DataPath_Physical_RF_n2171,
         dp_id_stage_regfile_DataPath_Physical_RF_n2170,
         dp_id_stage_regfile_DataPath_Physical_RF_n2169,
         dp_id_stage_regfile_DataPath_Physical_RF_n2168,
         dp_id_stage_regfile_DataPath_Physical_RF_n2167,
         dp_id_stage_regfile_DataPath_Physical_RF_n2166,
         dp_id_stage_regfile_DataPath_Physical_RF_n2165,
         dp_id_stage_regfile_DataPath_Physical_RF_n2164,
         dp_id_stage_regfile_DataPath_Physical_RF_n2163,
         dp_id_stage_regfile_DataPath_Physical_RF_n2162,
         dp_id_stage_regfile_DataPath_Physical_RF_n2161,
         dp_id_stage_regfile_DataPath_Physical_RF_n2160,
         dp_id_stage_regfile_DataPath_Physical_RF_n2159,
         dp_id_stage_regfile_DataPath_Physical_RF_n2158,
         dp_id_stage_regfile_DataPath_Physical_RF_n2157,
         dp_id_stage_regfile_DataPath_Physical_RF_n2156,
         dp_id_stage_regfile_DataPath_Physical_RF_n2155,
         dp_id_stage_regfile_DataPath_Physical_RF_n2154,
         dp_id_stage_regfile_DataPath_Physical_RF_n2153,
         dp_id_stage_regfile_DataPath_Physical_RF_n2152,
         dp_id_stage_regfile_DataPath_Physical_RF_n2151,
         dp_id_stage_regfile_DataPath_Physical_RF_n2150,
         dp_id_stage_regfile_DataPath_Physical_RF_n2149,
         dp_id_stage_regfile_DataPath_Physical_RF_n2148,
         dp_id_stage_regfile_DataPath_Physical_RF_n2147,
         dp_id_stage_regfile_DataPath_Physical_RF_n2146,
         dp_id_stage_regfile_DataPath_Physical_RF_n2145,
         dp_id_stage_regfile_DataPath_Physical_RF_n2144,
         dp_id_stage_regfile_DataPath_Physical_RF_n2143,
         dp_id_stage_regfile_DataPath_Physical_RF_n2142,
         dp_id_stage_regfile_DataPath_Physical_RF_n2141,
         dp_id_stage_regfile_DataPath_Physical_RF_n2140,
         dp_id_stage_regfile_DataPath_Physical_RF_n2139,
         dp_id_stage_regfile_DataPath_Physical_RF_n2138,
         dp_id_stage_regfile_DataPath_Physical_RF_n2137,
         dp_id_stage_regfile_DataPath_Physical_RF_n2136,
         dp_id_stage_regfile_DataPath_Physical_RF_n2135,
         dp_id_stage_regfile_DataPath_Physical_RF_n2134,
         dp_id_stage_regfile_DataPath_Physical_RF_n2133,
         dp_id_stage_regfile_DataPath_Physical_RF_n2132,
         dp_id_stage_regfile_DataPath_Physical_RF_n2131,
         dp_id_stage_regfile_DataPath_Physical_RF_n2130,
         dp_id_stage_regfile_DataPath_Physical_RF_n2129,
         dp_id_stage_regfile_DataPath_Physical_RF_n2128,
         dp_id_stage_regfile_DataPath_Physical_RF_n2127,
         dp_id_stage_regfile_DataPath_Physical_RF_n2126,
         dp_id_stage_regfile_DataPath_Physical_RF_n2125,
         dp_id_stage_regfile_DataPath_Physical_RF_n2124,
         dp_id_stage_regfile_DataPath_Physical_RF_n2123,
         dp_id_stage_regfile_DataPath_Physical_RF_n2122,
         dp_id_stage_regfile_DataPath_Physical_RF_n2121,
         dp_id_stage_regfile_DataPath_Physical_RF_n2120,
         dp_id_stage_regfile_DataPath_Physical_RF_n2119,
         dp_id_stage_regfile_DataPath_Physical_RF_n2118,
         dp_id_stage_regfile_DataPath_Physical_RF_n2117,
         dp_id_stage_regfile_DataPath_Physical_RF_n2116,
         dp_id_stage_regfile_DataPath_Physical_RF_n2115,
         dp_id_stage_regfile_DataPath_Physical_RF_n2114,
         dp_id_stage_regfile_DataPath_Physical_RF_n2113,
         dp_id_stage_regfile_DataPath_Physical_RF_n2112,
         dp_id_stage_regfile_DataPath_Physical_RF_n2111,
         dp_id_stage_regfile_DataPath_Physical_RF_n2110,
         dp_id_stage_regfile_DataPath_Physical_RF_n2109,
         dp_id_stage_regfile_DataPath_Physical_RF_n2108,
         dp_id_stage_regfile_DataPath_Physical_RF_n2107,
         dp_id_stage_regfile_DataPath_Physical_RF_n2106,
         dp_id_stage_regfile_DataPath_Physical_RF_n2105,
         dp_id_stage_regfile_DataPath_Physical_RF_n2104,
         dp_id_stage_regfile_DataPath_Physical_RF_n2103,
         dp_id_stage_regfile_DataPath_Physical_RF_n2102,
         dp_id_stage_regfile_DataPath_Physical_RF_n2101,
         dp_id_stage_regfile_DataPath_Physical_RF_n2100,
         dp_id_stage_regfile_DataPath_Physical_RF_n2099,
         dp_id_stage_regfile_DataPath_Physical_RF_n2098,
         dp_id_stage_regfile_DataPath_Physical_RF_n2097,
         dp_id_stage_regfile_DataPath_Physical_RF_n2096,
         dp_id_stage_regfile_DataPath_Physical_RF_n2095,
         dp_id_stage_regfile_DataPath_Physical_RF_n2094,
         dp_id_stage_regfile_DataPath_Physical_RF_n2093,
         dp_id_stage_regfile_DataPath_Physical_RF_n2092,
         dp_id_stage_regfile_DataPath_Physical_RF_n2091,
         dp_id_stage_regfile_DataPath_Physical_RF_n2090,
         dp_id_stage_regfile_DataPath_Physical_RF_n2089,
         dp_id_stage_regfile_DataPath_Physical_RF_n2088,
         dp_id_stage_regfile_DataPath_Physical_RF_n2087,
         dp_id_stage_regfile_DataPath_Physical_RF_n2086,
         dp_id_stage_regfile_DataPath_Physical_RF_n2085,
         dp_id_stage_regfile_DataPath_Physical_RF_n2084,
         dp_id_stage_regfile_DataPath_Physical_RF_n2083,
         dp_id_stage_regfile_DataPath_Physical_RF_n2082,
         dp_id_stage_regfile_DataPath_Physical_RF_n2081,
         dp_id_stage_regfile_DataPath_Physical_RF_n2080,
         dp_id_stage_regfile_DataPath_Physical_RF_n2079,
         dp_id_stage_regfile_DataPath_Physical_RF_n2078,
         dp_id_stage_regfile_DataPath_Physical_RF_n2077,
         dp_id_stage_regfile_DataPath_Physical_RF_n2076,
         dp_id_stage_regfile_DataPath_Physical_RF_n2075,
         dp_id_stage_regfile_DataPath_Physical_RF_n2074,
         dp_id_stage_regfile_DataPath_Physical_RF_n2073,
         dp_id_stage_regfile_DataPath_Physical_RF_n2072,
         dp_id_stage_regfile_DataPath_Physical_RF_n2071,
         dp_id_stage_regfile_DataPath_Physical_RF_n2070,
         dp_id_stage_regfile_DataPath_Physical_RF_n2069,
         dp_id_stage_regfile_DataPath_Physical_RF_n2068,
         dp_id_stage_regfile_DataPath_Physical_RF_n2067,
         dp_id_stage_regfile_DataPath_Physical_RF_n2066,
         dp_id_stage_regfile_DataPath_Physical_RF_n2065,
         dp_id_stage_regfile_DataPath_Physical_RF_n2064,
         dp_id_stage_regfile_DataPath_Physical_RF_n2063,
         dp_id_stage_regfile_DataPath_Physical_RF_n2062,
         dp_id_stage_regfile_DataPath_Physical_RF_n2061,
         dp_id_stage_regfile_DataPath_Physical_RF_n2060,
         dp_id_stage_regfile_DataPath_Physical_RF_n2059,
         dp_id_stage_regfile_DataPath_Physical_RF_n2058,
         dp_id_stage_regfile_DataPath_Physical_RF_n2057,
         dp_id_stage_regfile_DataPath_Physical_RF_n2056,
         dp_id_stage_regfile_DataPath_Physical_RF_n2055,
         dp_id_stage_regfile_DataPath_Physical_RF_n2054,
         dp_id_stage_regfile_DataPath_Physical_RF_n2053,
         dp_id_stage_regfile_DataPath_Physical_RF_n2052,
         dp_id_stage_regfile_DataPath_Physical_RF_n2051,
         dp_id_stage_regfile_DataPath_Physical_RF_n2050,
         dp_id_stage_regfile_DataPath_Physical_RF_n2049,
         dp_id_stage_regfile_DataPath_Physical_RF_n2048,
         dp_id_stage_regfile_DataPath_Physical_RF_n2047,
         dp_id_stage_regfile_DataPath_Physical_RF_n2046,
         dp_id_stage_regfile_DataPath_Physical_RF_n2045,
         dp_id_stage_regfile_DataPath_Physical_RF_n2044,
         dp_id_stage_regfile_DataPath_Physical_RF_n2043,
         dp_id_stage_regfile_DataPath_Physical_RF_n2042,
         dp_id_stage_regfile_DataPath_Physical_RF_n2041,
         dp_id_stage_regfile_DataPath_Physical_RF_n2040,
         dp_id_stage_regfile_DataPath_Physical_RF_n2039,
         dp_id_stage_regfile_DataPath_Physical_RF_n2038,
         dp_id_stage_regfile_DataPath_Physical_RF_n2037,
         dp_id_stage_regfile_DataPath_Physical_RF_n2036,
         dp_id_stage_regfile_DataPath_Physical_RF_n2035,
         dp_id_stage_regfile_DataPath_Physical_RF_n2034,
         dp_id_stage_regfile_DataPath_Physical_RF_n2033,
         dp_id_stage_regfile_DataPath_Physical_RF_n2032,
         dp_id_stage_regfile_DataPath_Physical_RF_n2031,
         dp_id_stage_regfile_DataPath_Physical_RF_n2030,
         dp_id_stage_regfile_DataPath_Physical_RF_n2029,
         dp_id_stage_regfile_DataPath_Physical_RF_n2028,
         dp_id_stage_regfile_DataPath_Physical_RF_n2027,
         dp_id_stage_regfile_DataPath_Physical_RF_n2026,
         dp_id_stage_regfile_DataPath_Physical_RF_n2025,
         dp_id_stage_regfile_DataPath_Physical_RF_n2024,
         dp_id_stage_regfile_DataPath_Physical_RF_n2023,
         dp_id_stage_regfile_DataPath_Physical_RF_n2022,
         dp_id_stage_regfile_DataPath_Physical_RF_n2021,
         dp_id_stage_regfile_DataPath_Physical_RF_n2020,
         dp_id_stage_regfile_DataPath_Physical_RF_n2019,
         dp_id_stage_regfile_DataPath_Physical_RF_n2018,
         dp_id_stage_regfile_DataPath_Physical_RF_n2017,
         dp_id_stage_regfile_DataPath_Physical_RF_n2016,
         dp_id_stage_regfile_DataPath_Physical_RF_n2015,
         dp_id_stage_regfile_DataPath_Physical_RF_n2014,
         dp_id_stage_regfile_DataPath_Physical_RF_n2013,
         dp_id_stage_regfile_DataPath_Physical_RF_n2012,
         dp_id_stage_regfile_DataPath_Physical_RF_n2011,
         dp_id_stage_regfile_DataPath_Physical_RF_n2010,
         dp_id_stage_regfile_DataPath_Physical_RF_n2009,
         dp_id_stage_regfile_DataPath_Physical_RF_n2008,
         dp_id_stage_regfile_DataPath_Physical_RF_n2007,
         dp_id_stage_regfile_DataPath_Physical_RF_n2006,
         dp_id_stage_regfile_DataPath_Physical_RF_n2005,
         dp_id_stage_regfile_DataPath_Physical_RF_n2004,
         dp_id_stage_regfile_DataPath_Physical_RF_n2003,
         dp_id_stage_regfile_DataPath_Physical_RF_n2002,
         dp_id_stage_regfile_DataPath_Physical_RF_n2001,
         dp_id_stage_regfile_DataPath_Physical_RF_n2000,
         dp_id_stage_regfile_DataPath_Physical_RF_n1999,
         dp_id_stage_regfile_DataPath_Physical_RF_n1998,
         dp_id_stage_regfile_DataPath_Physical_RF_n1997,
         dp_id_stage_regfile_DataPath_Physical_RF_n1996,
         dp_id_stage_regfile_DataPath_Physical_RF_n1995,
         dp_id_stage_regfile_DataPath_Physical_RF_n1994,
         dp_id_stage_regfile_DataPath_Physical_RF_n1993,
         dp_id_stage_regfile_DataPath_Physical_RF_n1992,
         dp_id_stage_regfile_DataPath_Physical_RF_n1991,
         dp_id_stage_regfile_DataPath_Physical_RF_n1990,
         dp_id_stage_regfile_DataPath_Physical_RF_n1989,
         dp_id_stage_regfile_DataPath_Physical_RF_n1988,
         dp_id_stage_regfile_DataPath_Physical_RF_n1987,
         dp_id_stage_regfile_DataPath_Physical_RF_n1986,
         dp_id_stage_regfile_DataPath_Physical_RF_n1985,
         dp_id_stage_regfile_DataPath_Physical_RF_n1984,
         dp_id_stage_regfile_DataPath_Physical_RF_n1983,
         dp_id_stage_regfile_DataPath_Physical_RF_n1982,
         dp_id_stage_regfile_DataPath_Physical_RF_n1981,
         dp_id_stage_regfile_DataPath_Physical_RF_n1980,
         dp_id_stage_regfile_DataPath_Physical_RF_n1979,
         dp_id_stage_regfile_DataPath_Physical_RF_n1978,
         dp_id_stage_regfile_DataPath_Physical_RF_n1977,
         dp_id_stage_regfile_DataPath_Physical_RF_n1976,
         dp_id_stage_regfile_DataPath_Physical_RF_n1975,
         dp_id_stage_regfile_DataPath_Physical_RF_n1974,
         dp_id_stage_regfile_DataPath_Physical_RF_n1973,
         dp_id_stage_regfile_DataPath_Physical_RF_n1972,
         dp_id_stage_regfile_DataPath_Physical_RF_n1971,
         dp_id_stage_regfile_DataPath_Physical_RF_n1970,
         dp_id_stage_regfile_DataPath_Physical_RF_n1969,
         dp_id_stage_regfile_DataPath_Physical_RF_n1968,
         dp_id_stage_regfile_DataPath_Physical_RF_n1967,
         dp_id_stage_regfile_DataPath_Physical_RF_n1966,
         dp_id_stage_regfile_DataPath_Physical_RF_n1965,
         dp_id_stage_regfile_DataPath_Physical_RF_n1964,
         dp_id_stage_regfile_DataPath_Physical_RF_n1963,
         dp_id_stage_regfile_DataPath_Physical_RF_n1962,
         dp_id_stage_regfile_DataPath_Physical_RF_n1961,
         dp_id_stage_regfile_DataPath_Physical_RF_n1960,
         dp_id_stage_regfile_DataPath_Physical_RF_n1959,
         dp_id_stage_regfile_DataPath_Physical_RF_n1958,
         dp_id_stage_regfile_DataPath_Physical_RF_n1957,
         dp_id_stage_regfile_DataPath_Physical_RF_n1956,
         dp_id_stage_regfile_DataPath_Physical_RF_n1955,
         dp_id_stage_regfile_DataPath_Physical_RF_n1954,
         dp_id_stage_regfile_DataPath_Physical_RF_n1953,
         dp_id_stage_regfile_DataPath_Physical_RF_n1952,
         dp_id_stage_regfile_DataPath_Physical_RF_n1951,
         dp_id_stage_regfile_DataPath_Physical_RF_n1950,
         dp_id_stage_regfile_DataPath_Physical_RF_n1949,
         dp_id_stage_regfile_DataPath_Physical_RF_n1948,
         dp_id_stage_regfile_DataPath_Physical_RF_n1947,
         dp_id_stage_regfile_DataPath_Physical_RF_n1946,
         dp_id_stage_regfile_DataPath_Physical_RF_n1945,
         dp_id_stage_regfile_DataPath_Physical_RF_n1944,
         dp_id_stage_regfile_DataPath_Physical_RF_n1943,
         dp_id_stage_regfile_DataPath_Physical_RF_n1942,
         dp_id_stage_regfile_DataPath_Physical_RF_n1941,
         dp_id_stage_regfile_DataPath_Physical_RF_n1940,
         dp_id_stage_regfile_DataPath_Physical_RF_n1939,
         dp_id_stage_regfile_DataPath_Physical_RF_n1938,
         dp_id_stage_regfile_DataPath_Physical_RF_n1937,
         dp_id_stage_regfile_DataPath_Physical_RF_n1936,
         dp_id_stage_regfile_DataPath_Physical_RF_n1935,
         dp_id_stage_regfile_DataPath_Physical_RF_n1934,
         dp_id_stage_regfile_DataPath_Physical_RF_n1933,
         dp_id_stage_regfile_DataPath_Physical_RF_n1932,
         dp_id_stage_regfile_DataPath_Physical_RF_n1931,
         dp_id_stage_regfile_DataPath_Physical_RF_n1930,
         dp_id_stage_regfile_DataPath_Physical_RF_n1929,
         dp_id_stage_regfile_DataPath_Physical_RF_n1928,
         dp_id_stage_regfile_DataPath_Physical_RF_n1927,
         dp_id_stage_regfile_DataPath_Physical_RF_n1924,
         dp_id_stage_regfile_DataPath_Physical_RF_n1923,
         dp_id_stage_regfile_DataPath_Physical_RF_n1922,
         dp_id_stage_regfile_DataPath_Physical_RF_n1921,
         dp_id_stage_regfile_DataPath_Physical_RF_n1920,
         dp_id_stage_regfile_DataPath_Physical_RF_n1919,
         dp_id_stage_regfile_DataPath_Physical_RF_n1918,
         dp_id_stage_regfile_DataPath_Physical_RF_n1917,
         dp_id_stage_regfile_DataPath_Physical_RF_n1916,
         dp_id_stage_regfile_DataPath_Physical_RF_n1915,
         dp_id_stage_regfile_DataPath_Physical_RF_n1914,
         dp_id_stage_regfile_DataPath_Physical_RF_n1913,
         dp_id_stage_regfile_DataPath_Physical_RF_n1912,
         dp_id_stage_regfile_DataPath_Physical_RF_n1911,
         dp_id_stage_regfile_DataPath_Physical_RF_n1910,
         dp_id_stage_regfile_DataPath_Physical_RF_n1909,
         dp_id_stage_regfile_DataPath_Physical_RF_n1908,
         dp_id_stage_regfile_DataPath_Physical_RF_n1907,
         dp_id_stage_regfile_DataPath_Physical_RF_n1906,
         dp_id_stage_regfile_DataPath_Physical_RF_n1905,
         dp_id_stage_regfile_DataPath_Physical_RF_n1904,
         dp_id_stage_regfile_DataPath_Physical_RF_n1903,
         dp_id_stage_regfile_DataPath_Physical_RF_n1902,
         dp_id_stage_regfile_DataPath_Physical_RF_n1901,
         dp_id_stage_regfile_DataPath_Physical_RF_n1900,
         dp_id_stage_regfile_DataPath_Physical_RF_n1899,
         dp_id_stage_regfile_DataPath_Physical_RF_n1898,
         dp_id_stage_regfile_DataPath_Physical_RF_n1897,
         dp_id_stage_regfile_DataPath_Physical_RF_n1896,
         dp_id_stage_regfile_DataPath_Physical_RF_n1895,
         dp_id_stage_regfile_DataPath_Physical_RF_n1894,
         dp_id_stage_regfile_DataPath_Physical_RF_n1893,
         dp_id_stage_regfile_DataPath_Physical_RF_n1892,
         dp_id_stage_regfile_DataPath_Physical_RF_n1891,
         dp_id_stage_regfile_DataPath_Physical_RF_n1890,
         dp_id_stage_regfile_DataPath_Physical_RF_n1889,
         dp_id_stage_regfile_DataPath_Physical_RF_n1888,
         dp_id_stage_regfile_DataPath_Physical_RF_n1887,
         dp_id_stage_regfile_DataPath_Physical_RF_n1886,
         dp_id_stage_regfile_DataPath_Physical_RF_n1885,
         dp_id_stage_regfile_DataPath_Physical_RF_n1884,
         dp_id_stage_regfile_DataPath_Physical_RF_n1883,
         dp_id_stage_regfile_DataPath_Physical_RF_n1882,
         dp_id_stage_regfile_DataPath_Physical_RF_n1881,
         dp_id_stage_regfile_DataPath_Physical_RF_n1880,
         dp_id_stage_regfile_DataPath_Physical_RF_n1879,
         dp_id_stage_regfile_DataPath_Physical_RF_n1878,
         dp_id_stage_regfile_DataPath_Physical_RF_n1877,
         dp_id_stage_regfile_DataPath_Physical_RF_n1876,
         dp_id_stage_regfile_DataPath_Physical_RF_n1875,
         dp_id_stage_regfile_DataPath_Physical_RF_n1874,
         dp_id_stage_regfile_DataPath_Physical_RF_n1873,
         dp_id_stage_regfile_DataPath_Physical_RF_n1872,
         dp_id_stage_regfile_DataPath_Physical_RF_n1871,
         dp_id_stage_regfile_DataPath_Physical_RF_n1870,
         dp_id_stage_regfile_DataPath_Physical_RF_n1869,
         dp_id_stage_regfile_DataPath_Physical_RF_n1868,
         dp_id_stage_regfile_DataPath_Physical_RF_n1867,
         dp_id_stage_regfile_DataPath_Physical_RF_n1866,
         dp_id_stage_regfile_DataPath_Physical_RF_n1865,
         dp_id_stage_regfile_DataPath_Physical_RF_n1864,
         dp_id_stage_regfile_DataPath_Physical_RF_n1863,
         dp_id_stage_regfile_DataPath_Physical_RF_n1862,
         dp_id_stage_regfile_DataPath_Physical_RF_n1861,
         dp_id_stage_regfile_DataPath_Physical_RF_n1860,
         dp_id_stage_regfile_DataPath_Physical_RF_n1859,
         dp_id_stage_regfile_DataPath_Physical_RF_n1856,
         dp_id_stage_regfile_DataPath_Physical_RF_n1855,
         dp_id_stage_regfile_DataPath_Physical_RF_n1854,
         dp_id_stage_regfile_DataPath_Physical_RF_n1853,
         dp_id_stage_regfile_DataPath_Physical_RF_n1852,
         dp_id_stage_regfile_DataPath_Physical_RF_n1851,
         dp_id_stage_regfile_DataPath_Physical_RF_n1850,
         dp_id_stage_regfile_DataPath_Physical_RF_n1849,
         dp_id_stage_regfile_DataPath_Physical_RF_n1848,
         dp_id_stage_regfile_DataPath_Physical_RF_n1847,
         dp_id_stage_regfile_DataPath_Physical_RF_n1846,
         dp_id_stage_regfile_DataPath_Physical_RF_n1845,
         dp_id_stage_regfile_DataPath_Physical_RF_n1844,
         dp_id_stage_regfile_DataPath_Physical_RF_n1843,
         dp_id_stage_regfile_DataPath_Physical_RF_n1842,
         dp_id_stage_regfile_DataPath_Physical_RF_n1841,
         dp_id_stage_regfile_DataPath_Physical_RF_n1840,
         dp_id_stage_regfile_DataPath_Physical_RF_n1839,
         dp_id_stage_regfile_DataPath_Physical_RF_n1838,
         dp_id_stage_regfile_DataPath_Physical_RF_n1837,
         dp_id_stage_regfile_DataPath_Physical_RF_n1836,
         dp_id_stage_regfile_DataPath_Physical_RF_n1835,
         dp_id_stage_regfile_DataPath_Physical_RF_n1834,
         dp_id_stage_regfile_DataPath_Physical_RF_n1833,
         dp_id_stage_regfile_DataPath_Physical_RF_n1832,
         dp_id_stage_regfile_DataPath_Physical_RF_n1831,
         dp_id_stage_regfile_DataPath_Physical_RF_n1830,
         dp_id_stage_regfile_DataPath_Physical_RF_n1829,
         dp_id_stage_regfile_DataPath_Physical_RF_n1828,
         dp_id_stage_regfile_DataPath_Physical_RF_n1827,
         dp_id_stage_regfile_DataPath_Physical_RF_n1826,
         dp_id_stage_regfile_DataPath_Physical_RF_n1825,
         dp_id_stage_regfile_DataPath_Physical_RF_n1824,
         dp_id_stage_regfile_DataPath_Physical_RF_n1823,
         dp_id_stage_regfile_DataPath_Physical_RF_n1822,
         dp_id_stage_regfile_DataPath_Physical_RF_n1821,
         dp_id_stage_regfile_DataPath_Physical_RF_n1820,
         dp_id_stage_regfile_DataPath_Physical_RF_n1819,
         dp_id_stage_regfile_DataPath_Physical_RF_n1818,
         dp_id_stage_regfile_DataPath_Physical_RF_n1817,
         dp_id_stage_regfile_DataPath_Physical_RF_n1816,
         dp_id_stage_regfile_DataPath_Physical_RF_n1815,
         dp_id_stage_regfile_DataPath_Physical_RF_n1814,
         dp_id_stage_regfile_DataPath_Physical_RF_n1813,
         dp_id_stage_regfile_DataPath_Physical_RF_n1812,
         dp_id_stage_regfile_DataPath_Physical_RF_n1811,
         dp_id_stage_regfile_DataPath_Physical_RF_n1810,
         dp_id_stage_regfile_DataPath_Physical_RF_n1809,
         dp_id_stage_regfile_DataPath_Physical_RF_n1808,
         dp_id_stage_regfile_DataPath_Physical_RF_n1807,
         dp_id_stage_regfile_DataPath_Physical_RF_n1806,
         dp_id_stage_regfile_DataPath_Physical_RF_n1805,
         dp_id_stage_regfile_DataPath_Physical_RF_n1804,
         dp_id_stage_regfile_DataPath_Physical_RF_n1803,
         dp_id_stage_regfile_DataPath_Physical_RF_n1802,
         dp_id_stage_regfile_DataPath_Physical_RF_n1801,
         dp_id_stage_regfile_DataPath_Physical_RF_n1800,
         dp_id_stage_regfile_DataPath_Physical_RF_n1799,
         dp_id_stage_regfile_DataPath_Physical_RF_n1798,
         dp_id_stage_regfile_DataPath_Physical_RF_n1797,
         dp_id_stage_regfile_DataPath_Physical_RF_n1796,
         dp_id_stage_regfile_DataPath_Physical_RF_n1795,
         dp_id_stage_regfile_DataPath_Physical_RF_n1794,
         dp_id_stage_regfile_DataPath_Physical_RF_n1793,
         dp_id_stage_regfile_DataPath_Physical_RF_n1792,
         dp_id_stage_regfile_DataPath_Physical_RF_n1791,
         dp_id_stage_regfile_DataPath_Physical_RF_n1790,
         dp_id_stage_regfile_DataPath_Physical_RF_n1789,
         dp_id_stage_regfile_DataPath_Physical_RF_n1788,
         dp_id_stage_regfile_DataPath_Physical_RF_n1787,
         dp_id_stage_regfile_DataPath_Physical_RF_n1786,
         dp_id_stage_regfile_DataPath_Physical_RF_n1785,
         dp_id_stage_regfile_DataPath_Physical_RF_n1784,
         dp_id_stage_regfile_DataPath_Physical_RF_n1783,
         dp_id_stage_regfile_DataPath_Physical_RF_n1782,
         dp_id_stage_regfile_DataPath_Physical_RF_n1781,
         dp_id_stage_regfile_DataPath_Physical_RF_n1780,
         dp_id_stage_regfile_DataPath_Physical_RF_n1779,
         dp_id_stage_regfile_DataPath_Physical_RF_n1778,
         dp_id_stage_regfile_DataPath_Physical_RF_n1777,
         dp_id_stage_regfile_DataPath_Physical_RF_n1776,
         dp_id_stage_regfile_DataPath_Physical_RF_n1775,
         dp_id_stage_regfile_DataPath_Physical_RF_n1774,
         dp_id_stage_regfile_DataPath_Physical_RF_n1773,
         dp_id_stage_regfile_DataPath_Physical_RF_n1772,
         dp_id_stage_regfile_DataPath_Physical_RF_n1771,
         dp_id_stage_regfile_DataPath_Physical_RF_n1770,
         dp_id_stage_regfile_DataPath_Physical_RF_n1769,
         dp_id_stage_regfile_DataPath_Physical_RF_n1768,
         dp_id_stage_regfile_DataPath_Physical_RF_n1767,
         dp_id_stage_regfile_DataPath_Physical_RF_n1766,
         dp_id_stage_regfile_DataPath_Physical_RF_n1765,
         dp_id_stage_regfile_DataPath_Physical_RF_n1764,
         dp_id_stage_regfile_DataPath_Physical_RF_n1763,
         dp_id_stage_regfile_DataPath_Physical_RF_n1762,
         dp_id_stage_regfile_DataPath_Physical_RF_n1761,
         dp_id_stage_regfile_DataPath_Physical_RF_n1760,
         dp_id_stage_regfile_DataPath_Physical_RF_n1759,
         dp_id_stage_regfile_DataPath_Physical_RF_n1758,
         dp_id_stage_regfile_DataPath_Physical_RF_n1757,
         dp_id_stage_regfile_DataPath_Physical_RF_n1754,
         dp_id_stage_regfile_DataPath_Physical_RF_n1753,
         dp_id_stage_regfile_DataPath_Physical_RF_n1752,
         dp_id_stage_regfile_DataPath_Physical_RF_n1751,
         dp_id_stage_regfile_DataPath_Physical_RF_n1750,
         dp_id_stage_regfile_DataPath_Physical_RF_n1749,
         dp_id_stage_regfile_DataPath_Physical_RF_n1748,
         dp_id_stage_regfile_DataPath_Physical_RF_n1747,
         dp_id_stage_regfile_DataPath_Physical_RF_n1746,
         dp_id_stage_regfile_DataPath_Physical_RF_n1745,
         dp_id_stage_regfile_DataPath_Physical_RF_n1744,
         dp_id_stage_regfile_DataPath_Physical_RF_n1743,
         dp_id_stage_regfile_DataPath_Physical_RF_n1742,
         dp_id_stage_regfile_DataPath_Physical_RF_n1741,
         dp_id_stage_regfile_DataPath_Physical_RF_n1740,
         dp_id_stage_regfile_DataPath_Physical_RF_n1739,
         dp_id_stage_regfile_DataPath_Physical_RF_n1738,
         dp_id_stage_regfile_DataPath_Physical_RF_n1737,
         dp_id_stage_regfile_DataPath_Physical_RF_n1736,
         dp_id_stage_regfile_DataPath_Physical_RF_n1735,
         dp_id_stage_regfile_DataPath_Physical_RF_n1734,
         dp_id_stage_regfile_DataPath_Physical_RF_n1733,
         dp_id_stage_regfile_DataPath_Physical_RF_n1732,
         dp_id_stage_regfile_DataPath_Physical_RF_n1731,
         dp_id_stage_regfile_DataPath_Physical_RF_n1730,
         dp_id_stage_regfile_DataPath_Physical_RF_n1729,
         dp_id_stage_regfile_DataPath_Physical_RF_n1728,
         dp_id_stage_regfile_DataPath_Physical_RF_n1727,
         dp_id_stage_regfile_DataPath_Physical_RF_n1726,
         dp_id_stage_regfile_DataPath_Physical_RF_n1725,
         dp_id_stage_regfile_DataPath_Physical_RF_n1724,
         dp_id_stage_regfile_DataPath_Physical_RF_n1723,
         dp_id_stage_regfile_DataPath_Physical_RF_n1722,
         dp_id_stage_regfile_DataPath_Physical_RF_n1721,
         dp_id_stage_regfile_DataPath_Physical_RF_n1720,
         dp_id_stage_regfile_DataPath_Physical_RF_n1719,
         dp_id_stage_regfile_DataPath_Physical_RF_n1718,
         dp_id_stage_regfile_DataPath_Physical_RF_n1717,
         dp_id_stage_regfile_DataPath_Physical_RF_n1716,
         dp_id_stage_regfile_DataPath_Physical_RF_n1715,
         dp_id_stage_regfile_DataPath_Physical_RF_n1714,
         dp_id_stage_regfile_DataPath_Physical_RF_n1713,
         dp_id_stage_regfile_DataPath_Physical_RF_n1712,
         dp_id_stage_regfile_DataPath_Physical_RF_n1711,
         dp_id_stage_regfile_DataPath_Physical_RF_n1710,
         dp_id_stage_regfile_DataPath_Physical_RF_n1709,
         dp_id_stage_regfile_DataPath_Physical_RF_n1708,
         dp_id_stage_regfile_DataPath_Physical_RF_n1707,
         dp_id_stage_regfile_DataPath_Physical_RF_n1706,
         dp_id_stage_regfile_DataPath_Physical_RF_n1705,
         dp_id_stage_regfile_DataPath_Physical_RF_n1704,
         dp_id_stage_regfile_DataPath_Physical_RF_n1703,
         dp_id_stage_regfile_DataPath_Physical_RF_n1702,
         dp_id_stage_regfile_DataPath_Physical_RF_n1701,
         dp_id_stage_regfile_DataPath_Physical_RF_n1700,
         dp_id_stage_regfile_DataPath_Physical_RF_n1699,
         dp_id_stage_regfile_DataPath_Physical_RF_n1698,
         dp_id_stage_regfile_DataPath_Physical_RF_n1697,
         dp_id_stage_regfile_DataPath_Physical_RF_n1696,
         dp_id_stage_regfile_DataPath_Physical_RF_n1695,
         dp_id_stage_regfile_DataPath_Physical_RF_n1694,
         dp_id_stage_regfile_DataPath_Physical_RF_n1693,
         dp_id_stage_regfile_DataPath_Physical_RF_n1692,
         dp_id_stage_regfile_DataPath_Physical_RF_n1691,
         dp_id_stage_regfile_DataPath_Physical_RF_n1690,
         dp_id_stage_regfile_DataPath_Physical_RF_n1689,
         dp_id_stage_regfile_DataPath_Physical_RF_n1686,
         dp_id_stage_regfile_DataPath_Physical_RF_n1685,
         dp_id_stage_regfile_DataPath_Physical_RF_n1684,
         dp_id_stage_regfile_DataPath_Physical_RF_n1683,
         dp_id_stage_regfile_DataPath_Physical_RF_n1682,
         dp_id_stage_regfile_DataPath_Physical_RF_n1681,
         dp_id_stage_regfile_DataPath_Physical_RF_n1680,
         dp_id_stage_regfile_DataPath_Physical_RF_n1679,
         dp_id_stage_regfile_DataPath_Physical_RF_n1678,
         dp_id_stage_regfile_DataPath_Physical_RF_n1677,
         dp_id_stage_regfile_DataPath_Physical_RF_n1676,
         dp_id_stage_regfile_DataPath_Physical_RF_n1675,
         dp_id_stage_regfile_DataPath_Physical_RF_n1674,
         dp_id_stage_regfile_DataPath_Physical_RF_n1673,
         dp_id_stage_regfile_DataPath_Physical_RF_n1672,
         dp_id_stage_regfile_DataPath_Physical_RF_n1671,
         dp_id_stage_regfile_DataPath_Physical_RF_n1670,
         dp_id_stage_regfile_DataPath_Physical_RF_n1669,
         dp_id_stage_regfile_DataPath_Physical_RF_n1668,
         dp_id_stage_regfile_DataPath_Physical_RF_n1667,
         dp_id_stage_regfile_DataPath_Physical_RF_n1666,
         dp_id_stage_regfile_DataPath_Physical_RF_n1665,
         dp_id_stage_regfile_DataPath_Physical_RF_n1664,
         dp_id_stage_regfile_DataPath_Physical_RF_n1663,
         dp_id_stage_regfile_DataPath_Physical_RF_n1662,
         dp_id_stage_regfile_DataPath_Physical_RF_n1661,
         dp_id_stage_regfile_DataPath_Physical_RF_n1660,
         dp_id_stage_regfile_DataPath_Physical_RF_n1659,
         dp_id_stage_regfile_DataPath_Physical_RF_n1658,
         dp_id_stage_regfile_DataPath_Physical_RF_n1657,
         dp_id_stage_regfile_DataPath_Physical_RF_n1656,
         dp_id_stage_regfile_DataPath_Physical_RF_n1655,
         dp_id_stage_regfile_DataPath_Physical_RF_n1654,
         dp_id_stage_regfile_DataPath_Physical_RF_n1653,
         dp_id_stage_regfile_DataPath_Physical_RF_n1652,
         dp_id_stage_regfile_DataPath_Physical_RF_n1651,
         dp_id_stage_regfile_DataPath_Physical_RF_n1650,
         dp_id_stage_regfile_DataPath_Physical_RF_n1649,
         dp_id_stage_regfile_DataPath_Physical_RF_n1648,
         dp_id_stage_regfile_DataPath_Physical_RF_n1647,
         dp_id_stage_regfile_DataPath_Physical_RF_n1646,
         dp_id_stage_regfile_DataPath_Physical_RF_n1645,
         dp_id_stage_regfile_DataPath_Physical_RF_n1644,
         dp_id_stage_regfile_DataPath_Physical_RF_n1643,
         dp_id_stage_regfile_DataPath_Physical_RF_n1642,
         dp_id_stage_regfile_DataPath_Physical_RF_n1641,
         dp_id_stage_regfile_DataPath_Physical_RF_n1640,
         dp_id_stage_regfile_DataPath_Physical_RF_n1639,
         dp_id_stage_regfile_DataPath_Physical_RF_n1638,
         dp_id_stage_regfile_DataPath_Physical_RF_n1637,
         dp_id_stage_regfile_DataPath_Physical_RF_n1636,
         dp_id_stage_regfile_DataPath_Physical_RF_n1635,
         dp_id_stage_regfile_DataPath_Physical_RF_n1634,
         dp_id_stage_regfile_DataPath_Physical_RF_n1633,
         dp_id_stage_regfile_DataPath_Physical_RF_n1632,
         dp_id_stage_regfile_DataPath_Physical_RF_n1631,
         dp_id_stage_regfile_DataPath_Physical_RF_n1630,
         dp_id_stage_regfile_DataPath_Physical_RF_n1629,
         dp_id_stage_regfile_DataPath_Physical_RF_n1628,
         dp_id_stage_regfile_DataPath_Physical_RF_n1627,
         dp_id_stage_regfile_DataPath_Physical_RF_n1626,
         dp_id_stage_regfile_DataPath_Physical_RF_n1625,
         dp_id_stage_regfile_DataPath_Physical_RF_n1624,
         dp_id_stage_regfile_DataPath_Physical_RF_n1623,
         dp_id_stage_regfile_DataPath_Physical_RF_n1622,
         dp_id_stage_regfile_DataPath_Physical_RF_n1621,
         dp_id_stage_regfile_DataPath_Physical_RF_n1620,
         dp_id_stage_regfile_DataPath_Physical_RF_n1619,
         dp_id_stage_regfile_DataPath_Physical_RF_n1618,
         dp_id_stage_regfile_DataPath_Physical_RF_n1617,
         dp_id_stage_regfile_DataPath_Physical_RF_n1616,
         dp_id_stage_regfile_DataPath_Physical_RF_n1615,
         dp_id_stage_regfile_DataPath_Physical_RF_n1614,
         dp_id_stage_regfile_DataPath_Physical_RF_n1613,
         dp_id_stage_regfile_DataPath_Physical_RF_n1612,
         dp_id_stage_regfile_DataPath_Physical_RF_n1611,
         dp_id_stage_regfile_DataPath_Physical_RF_n1610,
         dp_id_stage_regfile_DataPath_Physical_RF_n1609,
         dp_id_stage_regfile_DataPath_Physical_RF_n1608,
         dp_id_stage_regfile_DataPath_Physical_RF_n1607,
         dp_id_stage_regfile_DataPath_Physical_RF_n1606,
         dp_id_stage_regfile_DataPath_Physical_RF_n1605,
         dp_id_stage_regfile_DataPath_Physical_RF_n1604,
         dp_id_stage_regfile_DataPath_Physical_RF_n1603,
         dp_id_stage_regfile_DataPath_Physical_RF_n1602,
         dp_id_stage_regfile_DataPath_Physical_RF_n1601,
         dp_id_stage_regfile_DataPath_Physical_RF_n1600,
         dp_id_stage_regfile_DataPath_Physical_RF_n1599,
         dp_id_stage_regfile_DataPath_Physical_RF_n1598,
         dp_id_stage_regfile_DataPath_Physical_RF_n1597,
         dp_id_stage_regfile_DataPath_Physical_RF_n1596,
         dp_id_stage_regfile_DataPath_Physical_RF_n1595,
         dp_id_stage_regfile_DataPath_Physical_RF_n1594,
         dp_id_stage_regfile_DataPath_Physical_RF_n1593,
         dp_id_stage_regfile_DataPath_Physical_RF_n1592,
         dp_id_stage_regfile_DataPath_Physical_RF_n1591,
         dp_id_stage_regfile_DataPath_Physical_RF_n1590,
         dp_id_stage_regfile_DataPath_Physical_RF_n1589,
         dp_id_stage_regfile_DataPath_Physical_RF_n1588,
         dp_id_stage_regfile_DataPath_Physical_RF_n1587,
         dp_id_stage_regfile_DataPath_Physical_RF_n1584,
         dp_id_stage_regfile_DataPath_Physical_RF_n1583,
         dp_id_stage_regfile_DataPath_Physical_RF_n1582,
         dp_id_stage_regfile_DataPath_Physical_RF_n1581,
         dp_id_stage_regfile_DataPath_Physical_RF_n1580,
         dp_id_stage_regfile_DataPath_Physical_RF_n1579,
         dp_id_stage_regfile_DataPath_Physical_RF_n1578,
         dp_id_stage_regfile_DataPath_Physical_RF_n1577,
         dp_id_stage_regfile_DataPath_Physical_RF_n1576,
         dp_id_stage_regfile_DataPath_Physical_RF_n1575,
         dp_id_stage_regfile_DataPath_Physical_RF_n1574,
         dp_id_stage_regfile_DataPath_Physical_RF_n1573,
         dp_id_stage_regfile_DataPath_Physical_RF_n1572,
         dp_id_stage_regfile_DataPath_Physical_RF_n1571,
         dp_id_stage_regfile_DataPath_Physical_RF_n1570,
         dp_id_stage_regfile_DataPath_Physical_RF_n1569,
         dp_id_stage_regfile_DataPath_Physical_RF_n1568,
         dp_id_stage_regfile_DataPath_Physical_RF_n1567,
         dp_id_stage_regfile_DataPath_Physical_RF_n1566,
         dp_id_stage_regfile_DataPath_Physical_RF_n1565,
         dp_id_stage_regfile_DataPath_Physical_RF_n1564,
         dp_id_stage_regfile_DataPath_Physical_RF_n1563,
         dp_id_stage_regfile_DataPath_Physical_RF_n1562,
         dp_id_stage_regfile_DataPath_Physical_RF_n1561,
         dp_id_stage_regfile_DataPath_Physical_RF_n1560,
         dp_id_stage_regfile_DataPath_Physical_RF_n1559,
         dp_id_stage_regfile_DataPath_Physical_RF_n1558,
         dp_id_stage_regfile_DataPath_Physical_RF_n1557,
         dp_id_stage_regfile_DataPath_Physical_RF_n1556,
         dp_id_stage_regfile_DataPath_Physical_RF_n1555,
         dp_id_stage_regfile_DataPath_Physical_RF_n1554,
         dp_id_stage_regfile_DataPath_Physical_RF_n1553,
         dp_id_stage_regfile_DataPath_Physical_RF_n1552,
         dp_id_stage_regfile_DataPath_Physical_RF_n1551,
         dp_id_stage_regfile_DataPath_Physical_RF_n1550,
         dp_id_stage_regfile_DataPath_Physical_RF_n1549,
         dp_id_stage_regfile_DataPath_Physical_RF_n1548,
         dp_id_stage_regfile_DataPath_Physical_RF_n1547,
         dp_id_stage_regfile_DataPath_Physical_RF_n1546,
         dp_id_stage_regfile_DataPath_Physical_RF_n1545,
         dp_id_stage_regfile_DataPath_Physical_RF_n1544,
         dp_id_stage_regfile_DataPath_Physical_RF_n1543,
         dp_id_stage_regfile_DataPath_Physical_RF_n1542,
         dp_id_stage_regfile_DataPath_Physical_RF_n1541,
         dp_id_stage_regfile_DataPath_Physical_RF_n1540,
         dp_id_stage_regfile_DataPath_Physical_RF_n1539,
         dp_id_stage_regfile_DataPath_Physical_RF_n1538,
         dp_id_stage_regfile_DataPath_Physical_RF_n1537,
         dp_id_stage_regfile_DataPath_Physical_RF_n1536,
         dp_id_stage_regfile_DataPath_Physical_RF_n1535,
         dp_id_stage_regfile_DataPath_Physical_RF_n1534,
         dp_id_stage_regfile_DataPath_Physical_RF_n1533,
         dp_id_stage_regfile_DataPath_Physical_RF_n1532,
         dp_id_stage_regfile_DataPath_Physical_RF_n1531,
         dp_id_stage_regfile_DataPath_Physical_RF_n1530,
         dp_id_stage_regfile_DataPath_Physical_RF_n1529,
         dp_id_stage_regfile_DataPath_Physical_RF_n1528,
         dp_id_stage_regfile_DataPath_Physical_RF_n1527,
         dp_id_stage_regfile_DataPath_Physical_RF_n1526,
         dp_id_stage_regfile_DataPath_Physical_RF_n1525,
         dp_id_stage_regfile_DataPath_Physical_RF_n1524,
         dp_id_stage_regfile_DataPath_Physical_RF_n1523,
         dp_id_stage_regfile_DataPath_Physical_RF_n1522,
         dp_id_stage_regfile_DataPath_Physical_RF_n1521,
         dp_id_stage_regfile_DataPath_Physical_RF_n1520,
         dp_id_stage_regfile_DataPath_Physical_RF_n1519,
         dp_id_stage_regfile_DataPath_Physical_RF_n1517,
         dp_id_stage_regfile_DataPath_Physical_RF_n1515,
         dp_id_stage_regfile_DataPath_Physical_RF_n1514,
         dp_id_stage_regfile_DataPath_Physical_RF_n1513,
         dp_id_stage_regfile_DataPath_Physical_RF_n1512,
         dp_id_stage_regfile_DataPath_Physical_RF_n1511,
         dp_id_stage_regfile_DataPath_Physical_RF_n1510,
         dp_id_stage_regfile_DataPath_Physical_RF_n1509,
         dp_id_stage_regfile_DataPath_Physical_RF_n1508,
         dp_id_stage_regfile_DataPath_Physical_RF_n1507,
         dp_id_stage_regfile_DataPath_Physical_RF_n1506,
         dp_id_stage_regfile_DataPath_Physical_RF_n1505,
         dp_id_stage_regfile_DataPath_Physical_RF_n1504,
         dp_id_stage_regfile_DataPath_Physical_RF_n1503,
         dp_id_stage_regfile_DataPath_Physical_RF_n1502,
         dp_id_stage_regfile_DataPath_Physical_RF_n1501,
         dp_id_stage_regfile_DataPath_Physical_RF_n1500,
         dp_id_stage_regfile_DataPath_Physical_RF_n1499,
         dp_id_stage_regfile_DataPath_Physical_RF_n1498,
         dp_id_stage_regfile_DataPath_Physical_RF_n1497,
         dp_id_stage_regfile_DataPath_Physical_RF_n1496,
         dp_id_stage_regfile_DataPath_Physical_RF_n1495,
         dp_id_stage_regfile_DataPath_Physical_RF_n1494,
         dp_id_stage_regfile_DataPath_Physical_RF_n1493,
         dp_id_stage_regfile_DataPath_Physical_RF_n1492,
         dp_id_stage_regfile_DataPath_Physical_RF_n1491,
         dp_id_stage_regfile_DataPath_Physical_RF_n1490,
         dp_id_stage_regfile_DataPath_Physical_RF_n1489,
         dp_id_stage_regfile_DataPath_Physical_RF_n1488,
         dp_id_stage_regfile_DataPath_Physical_RF_n1487,
         dp_id_stage_regfile_DataPath_Physical_RF_n1486,
         dp_id_stage_regfile_DataPath_Physical_RF_n1485,
         dp_id_stage_regfile_DataPath_Physical_RF_n1484,
         dp_id_stage_regfile_DataPath_Physical_RF_n1483,
         dp_id_stage_regfile_DataPath_Physical_RF_n1482,
         dp_id_stage_regfile_DataPath_Physical_RF_n1481,
         dp_id_stage_regfile_DataPath_Physical_RF_n1480,
         dp_id_stage_regfile_DataPath_Physical_RF_n1479,
         dp_id_stage_regfile_DataPath_Physical_RF_n1478,
         dp_id_stage_regfile_DataPath_Physical_RF_n1477,
         dp_id_stage_regfile_DataPath_Physical_RF_n1476,
         dp_id_stage_regfile_DataPath_Physical_RF_n1475,
         dp_id_stage_regfile_DataPath_Physical_RF_n1474,
         dp_id_stage_regfile_DataPath_Physical_RF_n1473,
         dp_id_stage_regfile_DataPath_Physical_RF_n1472,
         dp_id_stage_regfile_DataPath_Physical_RF_n1471,
         dp_id_stage_regfile_DataPath_Physical_RF_n1470,
         dp_id_stage_regfile_DataPath_Physical_RF_n1469,
         dp_id_stage_regfile_DataPath_Physical_RF_n1468,
         dp_id_stage_regfile_DataPath_Physical_RF_n1467,
         dp_id_stage_regfile_DataPath_Physical_RF_n1466,
         dp_id_stage_regfile_DataPath_Physical_RF_n1465,
         dp_id_stage_regfile_DataPath_Physical_RF_n1464,
         dp_id_stage_regfile_DataPath_Physical_RF_n1463,
         dp_id_stage_regfile_DataPath_Physical_RF_n1462,
         dp_id_stage_regfile_DataPath_Physical_RF_n1461,
         dp_id_stage_regfile_DataPath_Physical_RF_n1460,
         dp_id_stage_regfile_DataPath_Physical_RF_n1459,
         dp_id_stage_regfile_DataPath_Physical_RF_n1458,
         dp_id_stage_regfile_DataPath_Physical_RF_n1457,
         dp_id_stage_regfile_DataPath_Physical_RF_n1456,
         dp_id_stage_regfile_DataPath_Physical_RF_n1455,
         dp_id_stage_regfile_DataPath_Physical_RF_n1454,
         dp_id_stage_regfile_DataPath_Physical_RF_n1453,
         dp_id_stage_regfile_DataPath_Physical_RF_n1452,
         dp_id_stage_regfile_DataPath_Physical_RF_n1451,
         dp_id_stage_regfile_DataPath_Physical_RF_n1450,
         dp_id_stage_regfile_DataPath_Physical_RF_n1449,
         dp_id_stage_regfile_DataPath_Physical_RF_n1448,
         dp_id_stage_regfile_DataPath_Physical_RF_n1447,
         dp_id_stage_regfile_DataPath_Physical_RF_n1446,
         dp_id_stage_regfile_DataPath_Physical_RF_n1445,
         dp_id_stage_regfile_DataPath_Physical_RF_n1444,
         dp_id_stage_regfile_DataPath_Physical_RF_n1443,
         dp_id_stage_regfile_DataPath_Physical_RF_n1442,
         dp_id_stage_regfile_DataPath_Physical_RF_n1441,
         dp_id_stage_regfile_DataPath_Physical_RF_n1440,
         dp_id_stage_regfile_DataPath_Physical_RF_n1439,
         dp_id_stage_regfile_DataPath_Physical_RF_n1438,
         dp_id_stage_regfile_DataPath_Physical_RF_n1437,
         dp_id_stage_regfile_DataPath_Physical_RF_n1436,
         dp_id_stage_regfile_DataPath_Physical_RF_n1435,
         dp_id_stage_regfile_DataPath_Physical_RF_n1434,
         dp_id_stage_regfile_DataPath_Physical_RF_n1433,
         dp_id_stage_regfile_DataPath_Physical_RF_n1432,
         dp_id_stage_regfile_DataPath_Physical_RF_n1431,
         dp_id_stage_regfile_DataPath_Physical_RF_n1430,
         dp_id_stage_regfile_DataPath_Physical_RF_n1429,
         dp_id_stage_regfile_DataPath_Physical_RF_n1428,
         dp_id_stage_regfile_DataPath_Physical_RF_n1427,
         dp_id_stage_regfile_DataPath_Physical_RF_n1426,
         dp_id_stage_regfile_DataPath_Physical_RF_n1425,
         dp_id_stage_regfile_DataPath_Physical_RF_n1424,
         dp_id_stage_regfile_DataPath_Physical_RF_n1423,
         dp_id_stage_regfile_DataPath_Physical_RF_n1422,
         dp_id_stage_regfile_DataPath_Physical_RF_n1421,
         dp_id_stage_regfile_DataPath_Physical_RF_n1420,
         dp_id_stage_regfile_DataPath_Physical_RF_n1419,
         dp_id_stage_regfile_DataPath_Physical_RF_n1418,
         dp_id_stage_regfile_DataPath_Physical_RF_n1417,
         dp_id_stage_regfile_DataPath_Physical_RF_n1416,
         dp_id_stage_regfile_DataPath_Physical_RF_n1415,
         dp_id_stage_regfile_DataPath_Physical_RF_n1414,
         dp_id_stage_regfile_DataPath_Physical_RF_n1413,
         dp_id_stage_regfile_DataPath_Physical_RF_n1412,
         dp_id_stage_regfile_DataPath_Physical_RF_n1411,
         dp_id_stage_regfile_DataPath_Physical_RF_n1410,
         dp_id_stage_regfile_DataPath_Physical_RF_n1409,
         dp_id_stage_regfile_DataPath_Physical_RF_n1408,
         dp_id_stage_regfile_DataPath_Physical_RF_n1407,
         dp_id_stage_regfile_DataPath_Physical_RF_n1406,
         dp_id_stage_regfile_DataPath_Physical_RF_n1405,
         dp_id_stage_regfile_DataPath_Physical_RF_n1404,
         dp_id_stage_regfile_DataPath_Physical_RF_n1403,
         dp_id_stage_regfile_DataPath_Physical_RF_n1402,
         dp_id_stage_regfile_DataPath_Physical_RF_n1401,
         dp_id_stage_regfile_DataPath_Physical_RF_n1400,
         dp_id_stage_regfile_DataPath_Physical_RF_n1399,
         dp_id_stage_regfile_DataPath_Physical_RF_n1398,
         dp_id_stage_regfile_DataPath_Physical_RF_n1397,
         dp_id_stage_regfile_DataPath_Physical_RF_n1396,
         dp_id_stage_regfile_DataPath_Physical_RF_n1395,
         dp_id_stage_regfile_DataPath_Physical_RF_n1394,
         dp_id_stage_regfile_DataPath_Physical_RF_n1393,
         dp_id_stage_regfile_DataPath_Physical_RF_n1392,
         dp_id_stage_regfile_DataPath_Physical_RF_n1391,
         dp_id_stage_regfile_DataPath_Physical_RF_n1390,
         dp_id_stage_regfile_DataPath_Physical_RF_n1389,
         dp_id_stage_regfile_DataPath_Physical_RF_n1388,
         dp_id_stage_regfile_DataPath_Physical_RF_n1387,
         dp_id_stage_regfile_DataPath_Physical_RF_n1386,
         dp_id_stage_regfile_DataPath_Physical_RF_n1385,
         dp_id_stage_regfile_DataPath_Physical_RF_n1384,
         dp_id_stage_regfile_DataPath_Physical_RF_n1383,
         dp_id_stage_regfile_DataPath_Physical_RF_n1382,
         dp_id_stage_regfile_DataPath_Physical_RF_n1381,
         dp_id_stage_regfile_DataPath_Physical_RF_n1380,
         dp_id_stage_regfile_DataPath_Physical_RF_n1379,
         dp_id_stage_regfile_DataPath_Physical_RF_n1378,
         dp_id_stage_regfile_DataPath_Physical_RF_n1377,
         dp_id_stage_regfile_DataPath_Physical_RF_n1376,
         dp_id_stage_regfile_DataPath_Physical_RF_n1375,
         dp_id_stage_regfile_DataPath_Physical_RF_n1374,
         dp_id_stage_regfile_DataPath_Physical_RF_n1373,
         dp_id_stage_regfile_DataPath_Physical_RF_n1372,
         dp_id_stage_regfile_DataPath_Physical_RF_n1371,
         dp_id_stage_regfile_DataPath_Physical_RF_n1370,
         dp_id_stage_regfile_DataPath_Physical_RF_n1369,
         dp_id_stage_regfile_DataPath_Physical_RF_n1368,
         dp_id_stage_regfile_DataPath_Physical_RF_n1367,
         dp_id_stage_regfile_DataPath_Physical_RF_n1366,
         dp_id_stage_regfile_DataPath_Physical_RF_n1365,
         dp_id_stage_regfile_DataPath_Physical_RF_n1364,
         dp_id_stage_regfile_DataPath_Physical_RF_n1363,
         dp_id_stage_regfile_DataPath_Physical_RF_n1362,
         dp_id_stage_regfile_DataPath_Physical_RF_n1361,
         dp_id_stage_regfile_DataPath_Physical_RF_n1360,
         dp_id_stage_regfile_DataPath_Physical_RF_n1359,
         dp_id_stage_regfile_DataPath_Physical_RF_n1358,
         dp_id_stage_regfile_DataPath_Physical_RF_n1357,
         dp_id_stage_regfile_DataPath_Physical_RF_n1356,
         dp_id_stage_regfile_DataPath_Physical_RF_n1355,
         dp_id_stage_regfile_DataPath_Physical_RF_n1354,
         dp_id_stage_regfile_DataPath_Physical_RF_n1353,
         dp_id_stage_regfile_DataPath_Physical_RF_n1352,
         dp_id_stage_regfile_DataPath_Physical_RF_n1351,
         dp_id_stage_regfile_DataPath_Physical_RF_n1350,
         dp_id_stage_regfile_DataPath_Physical_RF_n1349,
         dp_id_stage_regfile_DataPath_Physical_RF_n1347,
         dp_id_stage_regfile_DataPath_Physical_RF_n1345,
         dp_id_stage_regfile_DataPath_Physical_RF_n1344,
         dp_id_stage_regfile_DataPath_Physical_RF_n1342,
         dp_id_stage_regfile_DataPath_Physical_RF_n1341,
         dp_id_stage_regfile_DataPath_Physical_RF_n1339,
         dp_id_stage_regfile_DataPath_Physical_RF_n1338,
         dp_id_stage_regfile_DataPath_Physical_RF_n1337,
         dp_id_stage_regfile_DataPath_Physical_RF_n1336,
         dp_id_stage_regfile_DataPath_Physical_RF_n1335,
         dp_id_stage_regfile_DataPath_Physical_RF_n1334,
         dp_id_stage_regfile_DataPath_Physical_RF_n1333,
         dp_id_stage_regfile_DataPath_Physical_RF_n1332,
         dp_id_stage_regfile_DataPath_Physical_RF_n1331,
         dp_id_stage_regfile_DataPath_Physical_RF_n1330,
         dp_id_stage_regfile_DataPath_Physical_RF_n1329,
         dp_id_stage_regfile_DataPath_Physical_RF_n1328,
         dp_id_stage_regfile_DataPath_Physical_RF_n1327,
         dp_id_stage_regfile_DataPath_Physical_RF_n1326,
         dp_id_stage_regfile_DataPath_Physical_RF_n1325,
         dp_id_stage_regfile_DataPath_Physical_RF_n1324,
         dp_id_stage_regfile_DataPath_Physical_RF_n1323,
         dp_id_stage_regfile_DataPath_Physical_RF_n1322,
         dp_id_stage_regfile_DataPath_Physical_RF_n1321,
         dp_id_stage_regfile_DataPath_Physical_RF_n1320,
         dp_id_stage_regfile_DataPath_Physical_RF_n1319,
         dp_id_stage_regfile_DataPath_Physical_RF_n1318,
         dp_id_stage_regfile_DataPath_Physical_RF_n1317,
         dp_id_stage_regfile_DataPath_Physical_RF_n1316,
         dp_id_stage_regfile_DataPath_Physical_RF_n1315,
         dp_id_stage_regfile_DataPath_Physical_RF_n1314,
         dp_id_stage_regfile_DataPath_Physical_RF_n1313,
         dp_id_stage_regfile_DataPath_Physical_RF_n1312,
         dp_id_stage_regfile_DataPath_Physical_RF_n1311,
         dp_id_stage_regfile_DataPath_Physical_RF_n1310,
         dp_id_stage_regfile_DataPath_Physical_RF_n1309,
         dp_id_stage_regfile_DataPath_Physical_RF_n1308,
         dp_id_stage_regfile_DataPath_Physical_RF_n1307,
         dp_id_stage_regfile_DataPath_Physical_RF_n1306,
         dp_id_stage_regfile_DataPath_Physical_RF_n1305,
         dp_id_stage_regfile_DataPath_Physical_RF_n1304,
         dp_id_stage_regfile_DataPath_Physical_RF_n1303,
         dp_id_stage_regfile_DataPath_Physical_RF_n1302,
         dp_id_stage_regfile_DataPath_Physical_RF_n1301,
         dp_id_stage_regfile_DataPath_Physical_RF_n1300,
         dp_id_stage_regfile_DataPath_Physical_RF_n1299,
         dp_id_stage_regfile_DataPath_Physical_RF_n1298,
         dp_id_stage_regfile_DataPath_Physical_RF_n1297,
         dp_id_stage_regfile_DataPath_Physical_RF_n1296,
         dp_id_stage_regfile_DataPath_Physical_RF_n1295,
         dp_id_stage_regfile_DataPath_Physical_RF_n1294,
         dp_id_stage_regfile_DataPath_Physical_RF_n1293,
         dp_id_stage_regfile_DataPath_Physical_RF_n1292,
         dp_id_stage_regfile_DataPath_Physical_RF_n1291,
         dp_id_stage_regfile_DataPath_Physical_RF_n1290,
         dp_id_stage_regfile_DataPath_Physical_RF_n1289,
         dp_id_stage_regfile_DataPath_Physical_RF_n1288,
         dp_id_stage_regfile_DataPath_Physical_RF_n1287,
         dp_id_stage_regfile_DataPath_Physical_RF_n1286,
         dp_id_stage_regfile_DataPath_Physical_RF_n1285,
         dp_id_stage_regfile_DataPath_Physical_RF_n1284,
         dp_id_stage_regfile_DataPath_Physical_RF_n1283,
         dp_id_stage_regfile_DataPath_Physical_RF_n1282,
         dp_id_stage_regfile_DataPath_Physical_RF_n1281,
         dp_id_stage_regfile_DataPath_Physical_RF_n1280,
         dp_id_stage_regfile_DataPath_Physical_RF_n1279,
         dp_id_stage_regfile_DataPath_Physical_RF_n1278,
         dp_id_stage_regfile_DataPath_Physical_RF_n1277,
         dp_id_stage_regfile_DataPath_Physical_RF_n1276,
         dp_id_stage_regfile_DataPath_Physical_RF_n1275,
         dp_id_stage_regfile_DataPath_Physical_RF_n1274,
         dp_id_stage_regfile_DataPath_Physical_RF_n1273,
         dp_id_stage_regfile_DataPath_Physical_RF_n1272,
         dp_id_stage_regfile_DataPath_Physical_RF_n1271,
         dp_id_stage_regfile_DataPath_Physical_RF_n1270,
         dp_id_stage_regfile_DataPath_Physical_RF_n1269,
         dp_id_stage_regfile_DataPath_Physical_RF_n1268,
         dp_id_stage_regfile_DataPath_Physical_RF_n1267,
         dp_id_stage_regfile_DataPath_Physical_RF_n1266,
         dp_id_stage_regfile_DataPath_Physical_RF_n1265,
         dp_id_stage_regfile_DataPath_Physical_RF_n1264,
         dp_id_stage_regfile_DataPath_Physical_RF_n1263,
         dp_id_stage_regfile_DataPath_Physical_RF_n1262,
         dp_id_stage_regfile_DataPath_Physical_RF_n1261,
         dp_id_stage_regfile_DataPath_Physical_RF_n1260,
         dp_id_stage_regfile_DataPath_Physical_RF_n1259,
         dp_id_stage_regfile_DataPath_Physical_RF_n1258,
         dp_id_stage_regfile_DataPath_Physical_RF_n1257,
         dp_id_stage_regfile_DataPath_Physical_RF_n1256,
         dp_id_stage_regfile_DataPath_Physical_RF_n1255,
         dp_id_stage_regfile_DataPath_Physical_RF_n1254,
         dp_id_stage_regfile_DataPath_Physical_RF_n1253,
         dp_id_stage_regfile_DataPath_Physical_RF_n1252,
         dp_id_stage_regfile_DataPath_Physical_RF_n1251,
         dp_id_stage_regfile_DataPath_Physical_RF_n1250,
         dp_id_stage_regfile_DataPath_Physical_RF_n1249,
         dp_id_stage_regfile_DataPath_Physical_RF_n1248,
         dp_id_stage_regfile_DataPath_Physical_RF_n1247,
         dp_id_stage_regfile_DataPath_Physical_RF_n1246,
         dp_id_stage_regfile_DataPath_Physical_RF_n1245,
         dp_id_stage_regfile_DataPath_Physical_RF_n1244,
         dp_id_stage_regfile_DataPath_Physical_RF_n1243,
         dp_id_stage_regfile_DataPath_Physical_RF_n1242,
         dp_id_stage_regfile_DataPath_Physical_RF_n1241,
         dp_id_stage_regfile_DataPath_Physical_RF_n1240,
         dp_id_stage_regfile_DataPath_Physical_RF_n1239,
         dp_id_stage_regfile_DataPath_Physical_RF_n1238,
         dp_id_stage_regfile_DataPath_Physical_RF_n1237,
         dp_id_stage_regfile_DataPath_Physical_RF_n1201,
         dp_id_stage_regfile_DataPath_Physical_RF_n1199,
         dp_id_stage_regfile_DataPath_Physical_RF_n1198,
         dp_id_stage_regfile_DataPath_Physical_RF_n1197,
         dp_id_stage_regfile_DataPath_Physical_RF_n1196,
         dp_id_stage_regfile_DataPath_Physical_RF_n1195,
         dp_id_stage_regfile_DataPath_Physical_RF_n1194,
         dp_id_stage_regfile_DataPath_Physical_RF_n1193,
         dp_id_stage_regfile_DataPath_Physical_RF_n1192,
         dp_id_stage_regfile_DataPath_Physical_RF_n1191,
         dp_id_stage_regfile_DataPath_Physical_RF_n1190,
         dp_id_stage_regfile_DataPath_Physical_RF_n1153,
         dp_id_stage_regfile_DataPath_Physical_RF_n1152,
         dp_id_stage_regfile_DataPath_Physical_RF_n1151,
         dp_id_stage_regfile_DataPath_Physical_RF_n1150,
         dp_id_stage_regfile_DataPath_Physical_RF_n1149,
         dp_id_stage_regfile_DataPath_Physical_RF_n1148,
         dp_id_stage_regfile_DataPath_Physical_RF_n1147,
         dp_id_stage_regfile_DataPath_Physical_RF_n1146,
         dp_id_stage_regfile_DataPath_Physical_RF_n1145,
         dp_id_stage_regfile_DataPath_Physical_RF_n1144,
         dp_id_stage_regfile_DataPath_Physical_RF_n1143,
         dp_id_stage_regfile_DataPath_Physical_RF_n1142,
         dp_id_stage_regfile_DataPath_Physical_RF_n1141,
         dp_id_stage_regfile_DataPath_Physical_RF_n1140,
         dp_id_stage_regfile_DataPath_Physical_RF_n1139,
         dp_id_stage_regfile_DataPath_Physical_RF_n1138,
         dp_id_stage_regfile_DataPath_Physical_RF_n1137,
         dp_id_stage_regfile_DataPath_Physical_RF_n1136,
         dp_id_stage_regfile_DataPath_Physical_RF_n1135,
         dp_id_stage_regfile_DataPath_Physical_RF_n1134,
         dp_id_stage_regfile_DataPath_Physical_RF_n1133,
         dp_id_stage_regfile_DataPath_Physical_RF_n1132,
         dp_id_stage_regfile_DataPath_Physical_RF_n1131,
         dp_id_stage_regfile_DataPath_Physical_RF_n1130,
         dp_id_stage_regfile_DataPath_Physical_RF_n1129,
         dp_id_stage_regfile_DataPath_Physical_RF_n1128,
         dp_id_stage_regfile_DataPath_Physical_RF_n1127,
         dp_id_stage_regfile_DataPath_Physical_RF_n1126,
         dp_id_stage_regfile_DataPath_Physical_RF_n1125,
         dp_id_stage_regfile_DataPath_Physical_RF_n1124,
         dp_id_stage_regfile_DataPath_Physical_RF_n1123,
         dp_id_stage_regfile_DataPath_Physical_RF_n1122,
         dp_id_stage_regfile_DataPath_Physical_RF_n1121,
         dp_id_stage_regfile_DataPath_Physical_RF_n1120,
         dp_id_stage_regfile_DataPath_Physical_RF_n1119,
         dp_id_stage_regfile_DataPath_Physical_RF_n1118,
         dp_id_stage_regfile_DataPath_Physical_RF_n1117,
         dp_id_stage_regfile_DataPath_Physical_RF_n1116,
         dp_id_stage_regfile_DataPath_Physical_RF_n1115,
         dp_id_stage_regfile_DataPath_Physical_RF_n1114,
         dp_id_stage_regfile_DataPath_Physical_RF_n1113,
         dp_id_stage_regfile_DataPath_Physical_RF_n1112,
         dp_id_stage_regfile_DataPath_Physical_RF_n1111,
         dp_id_stage_regfile_DataPath_Physical_RF_n1110,
         dp_id_stage_regfile_DataPath_Physical_RF_n1109,
         dp_id_stage_regfile_DataPath_Physical_RF_n1108,
         dp_id_stage_regfile_DataPath_Physical_RF_n1107,
         dp_id_stage_regfile_DataPath_Physical_RF_n1106,
         dp_id_stage_regfile_DataPath_Physical_RF_n1105,
         dp_id_stage_regfile_DataPath_Physical_RF_n1104,
         dp_id_stage_regfile_DataPath_Physical_RF_n1103,
         dp_id_stage_regfile_DataPath_Physical_RF_n1102,
         dp_id_stage_regfile_DataPath_Physical_RF_n1101,
         dp_id_stage_regfile_DataPath_Physical_RF_n1100,
         dp_id_stage_regfile_DataPath_Physical_RF_n1099,
         dp_id_stage_regfile_DataPath_Physical_RF_n1098,
         dp_id_stage_regfile_DataPath_Physical_RF_n1097,
         dp_id_stage_regfile_DataPath_Physical_RF_n1096,
         dp_id_stage_regfile_DataPath_Physical_RF_n1095,
         dp_id_stage_regfile_DataPath_Physical_RF_n1094,
         dp_id_stage_regfile_DataPath_Physical_RF_n1093,
         dp_id_stage_regfile_DataPath_Physical_RF_n1092,
         dp_id_stage_regfile_DataPath_Physical_RF_n1091,
         dp_id_stage_regfile_DataPath_Physical_RF_n1090,
         dp_id_stage_regfile_DataPath_Physical_RF_n1089,
         dp_id_stage_regfile_DataPath_Physical_RF_n1088,
         dp_id_stage_regfile_DataPath_Physical_RF_n1087,
         dp_id_stage_regfile_DataPath_Physical_RF_n1086,
         dp_id_stage_regfile_DataPath_Physical_RF_n1085,
         dp_id_stage_regfile_DataPath_Physical_RF_n1084,
         dp_id_stage_regfile_DataPath_Physical_RF_n1083,
         dp_id_stage_regfile_DataPath_Physical_RF_n1082,
         dp_id_stage_regfile_DataPath_Physical_RF_n1081,
         dp_id_stage_regfile_DataPath_Physical_RF_n1080,
         dp_id_stage_regfile_DataPath_Physical_RF_n1079,
         dp_id_stage_regfile_DataPath_Physical_RF_n1078,
         dp_id_stage_regfile_DataPath_Physical_RF_n1077,
         dp_id_stage_regfile_DataPath_Physical_RF_n1076,
         dp_id_stage_regfile_DataPath_Physical_RF_n1075,
         dp_id_stage_regfile_DataPath_Physical_RF_n1074,
         dp_id_stage_regfile_DataPath_Physical_RF_n1073,
         dp_id_stage_regfile_DataPath_Physical_RF_n1072,
         dp_id_stage_regfile_DataPath_Physical_RF_n1071,
         dp_id_stage_regfile_DataPath_Physical_RF_n1070,
         dp_id_stage_regfile_DataPath_Physical_RF_n1069,
         dp_id_stage_regfile_DataPath_Physical_RF_n1068,
         dp_id_stage_regfile_DataPath_Physical_RF_n1067,
         dp_id_stage_regfile_DataPath_Physical_RF_n1066,
         dp_id_stage_regfile_DataPath_Physical_RF_n1065,
         dp_id_stage_regfile_DataPath_Physical_RF_n1064,
         dp_id_stage_regfile_DataPath_Physical_RF_n1063,
         dp_id_stage_regfile_DataPath_Physical_RF_n1062,
         dp_id_stage_regfile_DataPath_Physical_RF_n1061,
         dp_id_stage_regfile_DataPath_Physical_RF_n1060,
         dp_id_stage_regfile_DataPath_Physical_RF_n1059,
         dp_id_stage_regfile_DataPath_Physical_RF_n1058,
         dp_id_stage_regfile_DataPath_Physical_RF_n1057,
         dp_id_stage_regfile_DataPath_Physical_RF_n1056,
         dp_id_stage_regfile_DataPath_Physical_RF_n1055,
         dp_id_stage_regfile_DataPath_Physical_RF_n1054,
         dp_id_stage_regfile_DataPath_Physical_RF_n1053,
         dp_id_stage_regfile_DataPath_Physical_RF_n1052,
         dp_id_stage_regfile_DataPath_Physical_RF_n1051,
         dp_id_stage_regfile_DataPath_Physical_RF_n1050,
         dp_id_stage_regfile_DataPath_Physical_RF_n1049,
         dp_id_stage_regfile_DataPath_Physical_RF_n1048,
         dp_id_stage_regfile_DataPath_Physical_RF_n1047,
         dp_id_stage_regfile_DataPath_Physical_RF_n1046,
         dp_id_stage_regfile_DataPath_Physical_RF_n1045,
         dp_id_stage_regfile_DataPath_Physical_RF_n1044,
         dp_id_stage_regfile_DataPath_Physical_RF_n1043,
         dp_id_stage_regfile_DataPath_Physical_RF_n1042,
         dp_id_stage_regfile_DataPath_Physical_RF_n1041,
         dp_id_stage_regfile_DataPath_Physical_RF_n1040,
         dp_id_stage_regfile_DataPath_Physical_RF_n1039,
         dp_id_stage_regfile_DataPath_Physical_RF_n1038,
         dp_id_stage_regfile_DataPath_Physical_RF_n1037,
         dp_id_stage_regfile_DataPath_Physical_RF_n1036,
         dp_id_stage_regfile_DataPath_Physical_RF_n1035,
         dp_id_stage_regfile_DataPath_Physical_RF_n1034,
         dp_id_stage_regfile_DataPath_Physical_RF_n1033,
         dp_id_stage_regfile_DataPath_Physical_RF_n1032,
         dp_id_stage_regfile_DataPath_Physical_RF_n1031,
         dp_id_stage_regfile_DataPath_Physical_RF_n1030,
         dp_id_stage_regfile_DataPath_Physical_RF_n1029,
         dp_id_stage_regfile_DataPath_Physical_RF_n1028,
         dp_id_stage_regfile_DataPath_Physical_RF_n1027,
         dp_id_stage_regfile_DataPath_Physical_RF_n1026,
         dp_id_stage_regfile_DataPath_Physical_RF_n1025,
         dp_id_stage_regfile_DataPath_Physical_RF_n1024,
         dp_id_stage_regfile_DataPath_Physical_RF_n1023,
         dp_id_stage_regfile_DataPath_Physical_RF_n1022,
         dp_id_stage_regfile_DataPath_Physical_RF_n1021,
         dp_id_stage_regfile_DataPath_Physical_RF_n1020,
         dp_id_stage_regfile_DataPath_Physical_RF_n1019,
         dp_id_stage_regfile_DataPath_Physical_RF_n1018,
         dp_id_stage_regfile_DataPath_Physical_RF_n1017,
         dp_id_stage_regfile_DataPath_Physical_RF_n1016,
         dp_id_stage_regfile_DataPath_Physical_RF_n1015,
         dp_id_stage_regfile_DataPath_Physical_RF_n1014,
         dp_id_stage_regfile_DataPath_Physical_RF_n1013,
         dp_id_stage_regfile_DataPath_Physical_RF_n1012,
         dp_id_stage_regfile_DataPath_Physical_RF_n1011,
         dp_id_stage_regfile_DataPath_Physical_RF_n1010,
         dp_id_stage_regfile_DataPath_Physical_RF_n1009,
         dp_id_stage_regfile_DataPath_Physical_RF_n1008,
         dp_id_stage_regfile_DataPath_Physical_RF_n1007,
         dp_id_stage_regfile_DataPath_Physical_RF_n1006,
         dp_id_stage_regfile_DataPath_Physical_RF_n1005,
         dp_id_stage_regfile_DataPath_Physical_RF_n1004,
         dp_id_stage_regfile_DataPath_Physical_RF_n1003,
         dp_id_stage_regfile_DataPath_Physical_RF_n1002,
         dp_id_stage_regfile_DataPath_Physical_RF_n1001,
         dp_id_stage_regfile_DataPath_Physical_RF_n1000,
         dp_id_stage_regfile_DataPath_Physical_RF_n999,
         dp_id_stage_regfile_DataPath_Physical_RF_n998,
         dp_id_stage_regfile_DataPath_Physical_RF_n997,
         dp_id_stage_regfile_DataPath_Physical_RF_n996,
         dp_id_stage_regfile_DataPath_Physical_RF_n995,
         dp_id_stage_regfile_DataPath_Physical_RF_n994,
         dp_id_stage_regfile_DataPath_Physical_RF_n993,
         dp_id_stage_regfile_DataPath_Physical_RF_n992,
         dp_id_stage_regfile_DataPath_Physical_RF_n991,
         dp_id_stage_regfile_DataPath_Physical_RF_n990,
         dp_id_stage_regfile_DataPath_Physical_RF_n989,
         dp_id_stage_regfile_DataPath_Physical_RF_n988,
         dp_id_stage_regfile_DataPath_Physical_RF_n987,
         dp_id_stage_regfile_DataPath_Physical_RF_n986,
         dp_id_stage_regfile_DataPath_Physical_RF_n985,
         dp_id_stage_regfile_DataPath_Physical_RF_n984,
         dp_id_stage_regfile_DataPath_Physical_RF_n983,
         dp_id_stage_regfile_DataPath_Physical_RF_n982,
         dp_id_stage_regfile_DataPath_Physical_RF_n981,
         dp_id_stage_regfile_DataPath_Physical_RF_n980,
         dp_id_stage_regfile_DataPath_Physical_RF_n979,
         dp_id_stage_regfile_DataPath_Physical_RF_n978,
         dp_id_stage_regfile_DataPath_Physical_RF_n977,
         dp_id_stage_regfile_DataPath_Physical_RF_n976,
         dp_id_stage_regfile_DataPath_Physical_RF_n975,
         dp_id_stage_regfile_DataPath_Physical_RF_n974,
         dp_id_stage_regfile_DataPath_Physical_RF_n973,
         dp_id_stage_regfile_DataPath_Physical_RF_n972,
         dp_id_stage_regfile_DataPath_Physical_RF_n971,
         dp_id_stage_regfile_DataPath_Physical_RF_n970,
         dp_id_stage_regfile_DataPath_Physical_RF_n969,
         dp_id_stage_regfile_DataPath_Physical_RF_n968,
         dp_id_stage_regfile_DataPath_Physical_RF_n967,
         dp_id_stage_regfile_DataPath_Physical_RF_n966,
         dp_id_stage_regfile_DataPath_Physical_RF_n965,
         dp_id_stage_regfile_DataPath_Physical_RF_n964,
         dp_id_stage_regfile_DataPath_Physical_RF_n963,
         dp_id_stage_regfile_DataPath_Physical_RF_n962,
         dp_id_stage_regfile_DataPath_Physical_RF_n961,
         dp_id_stage_regfile_DataPath_Physical_RF_n960,
         dp_id_stage_regfile_DataPath_Physical_RF_n959,
         dp_id_stage_regfile_DataPath_Physical_RF_n958,
         dp_id_stage_regfile_DataPath_Physical_RF_n957,
         dp_id_stage_regfile_DataPath_Physical_RF_n956,
         dp_id_stage_regfile_DataPath_Physical_RF_n955,
         dp_id_stage_regfile_DataPath_Physical_RF_n954,
         dp_id_stage_regfile_DataPath_Physical_RF_n953,
         dp_id_stage_regfile_DataPath_Physical_RF_n952,
         dp_id_stage_regfile_DataPath_Physical_RF_n951,
         dp_id_stage_regfile_DataPath_Physical_RF_n950,
         dp_id_stage_regfile_DataPath_Physical_RF_n949,
         dp_id_stage_regfile_DataPath_Physical_RF_n948,
         dp_id_stage_regfile_DataPath_Physical_RF_n947,
         dp_id_stage_regfile_DataPath_Physical_RF_n946,
         dp_id_stage_regfile_DataPath_Physical_RF_n945,
         dp_id_stage_regfile_DataPath_Physical_RF_n944,
         dp_id_stage_regfile_DataPath_Physical_RF_n943,
         dp_id_stage_regfile_DataPath_Physical_RF_n942,
         dp_id_stage_regfile_DataPath_Physical_RF_n941,
         dp_id_stage_regfile_DataPath_Physical_RF_n940,
         dp_id_stage_regfile_DataPath_Physical_RF_n939,
         dp_id_stage_regfile_DataPath_Physical_RF_n938,
         dp_id_stage_regfile_DataPath_Physical_RF_n937,
         dp_id_stage_regfile_DataPath_Physical_RF_n936,
         dp_id_stage_regfile_DataPath_Physical_RF_n935,
         dp_id_stage_regfile_DataPath_Physical_RF_n934,
         dp_id_stage_regfile_DataPath_Physical_RF_n933,
         dp_id_stage_regfile_DataPath_Physical_RF_n932,
         dp_id_stage_regfile_DataPath_Physical_RF_n931,
         dp_id_stage_regfile_DataPath_Physical_RF_n930,
         dp_id_stage_regfile_DataPath_Physical_RF_n929,
         dp_id_stage_regfile_DataPath_Physical_RF_n928,
         dp_id_stage_regfile_DataPath_Physical_RF_n927,
         dp_id_stage_regfile_DataPath_Physical_RF_n926,
         dp_id_stage_regfile_DataPath_Physical_RF_n925,
         dp_id_stage_regfile_DataPath_Physical_RF_n924,
         dp_id_stage_regfile_DataPath_Physical_RF_n923,
         dp_id_stage_regfile_DataPath_Physical_RF_n922,
         dp_id_stage_regfile_DataPath_Physical_RF_n921,
         dp_id_stage_regfile_DataPath_Physical_RF_n920,
         dp_id_stage_regfile_DataPath_Physical_RF_n919,
         dp_id_stage_regfile_DataPath_Physical_RF_n918,
         dp_id_stage_regfile_DataPath_Physical_RF_n917,
         dp_id_stage_regfile_DataPath_Physical_RF_n916,
         dp_id_stage_regfile_DataPath_Physical_RF_n915,
         dp_id_stage_regfile_DataPath_Physical_RF_n914,
         dp_id_stage_regfile_DataPath_Physical_RF_n913,
         dp_id_stage_regfile_DataPath_Physical_RF_n912,
         dp_id_stage_regfile_DataPath_Physical_RF_n911,
         dp_id_stage_regfile_DataPath_Physical_RF_n910,
         dp_id_stage_regfile_DataPath_Physical_RF_n909,
         dp_id_stage_regfile_DataPath_Physical_RF_n908,
         dp_id_stage_regfile_DataPath_Physical_RF_n907,
         dp_id_stage_regfile_DataPath_Physical_RF_n906,
         dp_id_stage_regfile_DataPath_Physical_RF_n905,
         dp_id_stage_regfile_DataPath_Physical_RF_n904,
         dp_id_stage_regfile_DataPath_Physical_RF_n903,
         dp_id_stage_regfile_DataPath_Physical_RF_n902,
         dp_id_stage_regfile_DataPath_Physical_RF_n901,
         dp_id_stage_regfile_DataPath_Physical_RF_n900,
         dp_id_stage_regfile_DataPath_Physical_RF_n899,
         dp_id_stage_regfile_DataPath_Physical_RF_n898,
         dp_id_stage_regfile_DataPath_Physical_RF_n897,
         dp_id_stage_regfile_DataPath_Physical_RF_n896,
         dp_id_stage_regfile_DataPath_Physical_RF_n895,
         dp_id_stage_regfile_DataPath_Physical_RF_n894,
         dp_id_stage_regfile_DataPath_Physical_RF_n893,
         dp_id_stage_regfile_DataPath_Physical_RF_n892,
         dp_id_stage_regfile_DataPath_Physical_RF_n891,
         dp_id_stage_regfile_DataPath_Physical_RF_n890,
         dp_id_stage_regfile_DataPath_Physical_RF_n889,
         dp_id_stage_regfile_DataPath_Physical_RF_n888,
         dp_id_stage_regfile_DataPath_Physical_RF_n887,
         dp_id_stage_regfile_DataPath_Physical_RF_n886,
         dp_id_stage_regfile_DataPath_Physical_RF_n885,
         dp_id_stage_regfile_DataPath_Physical_RF_n884,
         dp_id_stage_regfile_DataPath_Physical_RF_n883,
         dp_id_stage_regfile_DataPath_Physical_RF_n882,
         dp_id_stage_regfile_DataPath_Physical_RF_n881,
         dp_id_stage_regfile_DataPath_Physical_RF_n880,
         dp_id_stage_regfile_DataPath_Physical_RF_n879,
         dp_id_stage_regfile_DataPath_Physical_RF_n878,
         dp_id_stage_regfile_DataPath_Physical_RF_n877,
         dp_id_stage_regfile_DataPath_Physical_RF_n876,
         dp_id_stage_regfile_DataPath_Physical_RF_n875,
         dp_id_stage_regfile_DataPath_Physical_RF_n874,
         dp_id_stage_regfile_DataPath_Physical_RF_n873,
         dp_id_stage_regfile_DataPath_Physical_RF_n872,
         dp_id_stage_regfile_DataPath_Physical_RF_n871,
         dp_id_stage_regfile_DataPath_Physical_RF_n870,
         dp_id_stage_regfile_DataPath_Physical_RF_n869,
         dp_id_stage_regfile_DataPath_Physical_RF_n868,
         dp_id_stage_regfile_DataPath_Physical_RF_n867,
         dp_id_stage_regfile_DataPath_Physical_RF_n866,
         dp_id_stage_regfile_DataPath_Physical_RF_n865,
         dp_id_stage_regfile_DataPath_Physical_RF_n864,
         dp_id_stage_regfile_DataPath_Physical_RF_n863,
         dp_id_stage_regfile_DataPath_Physical_RF_n862,
         dp_id_stage_regfile_DataPath_Physical_RF_n861,
         dp_id_stage_regfile_DataPath_Physical_RF_n860,
         dp_id_stage_regfile_DataPath_Physical_RF_n859,
         dp_id_stage_regfile_DataPath_Physical_RF_n858,
         dp_id_stage_regfile_DataPath_Physical_RF_n857,
         dp_id_stage_regfile_DataPath_Physical_RF_n856,
         dp_id_stage_regfile_DataPath_Physical_RF_n855,
         dp_id_stage_regfile_DataPath_Physical_RF_n854,
         dp_id_stage_regfile_DataPath_Physical_RF_n853,
         dp_id_stage_regfile_DataPath_Physical_RF_n852,
         dp_id_stage_regfile_DataPath_Physical_RF_n851,
         dp_id_stage_regfile_DataPath_Physical_RF_n850,
         dp_id_stage_regfile_DataPath_Physical_RF_n849,
         dp_id_stage_regfile_DataPath_Physical_RF_n848,
         dp_id_stage_regfile_DataPath_Physical_RF_n847,
         dp_id_stage_regfile_DataPath_Physical_RF_n846,
         dp_id_stage_regfile_DataPath_Physical_RF_n845,
         dp_id_stage_regfile_DataPath_Physical_RF_n844,
         dp_id_stage_regfile_DataPath_Physical_RF_n843,
         dp_id_stage_regfile_DataPath_Physical_RF_n842,
         dp_id_stage_regfile_DataPath_Physical_RF_n841,
         dp_id_stage_regfile_DataPath_Physical_RF_n840,
         dp_id_stage_regfile_DataPath_Physical_RF_n839,
         dp_id_stage_regfile_DataPath_Physical_RF_n838,
         dp_id_stage_regfile_DataPath_Physical_RF_n837,
         dp_id_stage_regfile_DataPath_Physical_RF_n836,
         dp_id_stage_regfile_DataPath_Physical_RF_n835,
         dp_id_stage_regfile_DataPath_Physical_RF_n834,
         dp_id_stage_regfile_DataPath_Physical_RF_n833,
         dp_id_stage_regfile_DataPath_Physical_RF_n832,
         dp_id_stage_regfile_DataPath_Physical_RF_n831,
         dp_id_stage_regfile_DataPath_Physical_RF_n830,
         dp_id_stage_regfile_DataPath_Physical_RF_n829,
         dp_id_stage_regfile_DataPath_Physical_RF_n828,
         dp_id_stage_regfile_DataPath_Physical_RF_n827,
         dp_id_stage_regfile_DataPath_Physical_RF_n826,
         dp_id_stage_regfile_DataPath_Physical_RF_n825,
         dp_id_stage_regfile_DataPath_Physical_RF_n824,
         dp_id_stage_regfile_DataPath_Physical_RF_n823,
         dp_id_stage_regfile_DataPath_Physical_RF_n822,
         dp_id_stage_regfile_DataPath_Physical_RF_n821,
         dp_id_stage_regfile_DataPath_Physical_RF_n820,
         dp_id_stage_regfile_DataPath_Physical_RF_n819,
         dp_id_stage_regfile_DataPath_Physical_RF_n818,
         dp_id_stage_regfile_DataPath_Physical_RF_n817,
         dp_id_stage_regfile_DataPath_Physical_RF_n816,
         dp_id_stage_regfile_DataPath_Physical_RF_n815,
         dp_id_stage_regfile_DataPath_Physical_RF_n814,
         dp_id_stage_regfile_DataPath_Physical_RF_n813,
         dp_id_stage_regfile_DataPath_Physical_RF_n812,
         dp_id_stage_regfile_DataPath_Physical_RF_n811,
         dp_id_stage_regfile_DataPath_Physical_RF_n810,
         dp_id_stage_regfile_DataPath_Physical_RF_n809,
         dp_id_stage_regfile_DataPath_Physical_RF_n808,
         dp_id_stage_regfile_DataPath_Physical_RF_n807,
         dp_id_stage_regfile_DataPath_Physical_RF_n806,
         dp_id_stage_regfile_DataPath_Physical_RF_n805,
         dp_id_stage_regfile_DataPath_Physical_RF_n804,
         dp_id_stage_regfile_DataPath_Physical_RF_n803,
         dp_id_stage_regfile_DataPath_Physical_RF_n802,
         dp_id_stage_regfile_DataPath_Physical_RF_n801,
         dp_id_stage_regfile_DataPath_Physical_RF_n800,
         dp_id_stage_regfile_DataPath_Physical_RF_n799,
         dp_id_stage_regfile_DataPath_Physical_RF_n798,
         dp_id_stage_regfile_DataPath_Physical_RF_n797,
         dp_id_stage_regfile_DataPath_Physical_RF_n796,
         dp_id_stage_regfile_DataPath_Physical_RF_n795,
         dp_id_stage_regfile_DataPath_Physical_RF_n794,
         dp_id_stage_regfile_DataPath_Physical_RF_n793,
         dp_id_stage_regfile_DataPath_Physical_RF_n792,
         dp_id_stage_regfile_DataPath_Physical_RF_n791,
         dp_id_stage_regfile_DataPath_Physical_RF_n790,
         dp_id_stage_regfile_DataPath_Physical_RF_n789,
         dp_id_stage_regfile_DataPath_Physical_RF_n788,
         dp_id_stage_regfile_DataPath_Physical_RF_n787,
         dp_id_stage_regfile_DataPath_Physical_RF_n786,
         dp_id_stage_regfile_DataPath_Physical_RF_n785,
         dp_id_stage_regfile_DataPath_Physical_RF_n784,
         dp_id_stage_regfile_DataPath_Physical_RF_n783,
         dp_id_stage_regfile_DataPath_Physical_RF_n782,
         dp_id_stage_regfile_DataPath_Physical_RF_n781,
         dp_id_stage_regfile_DataPath_Physical_RF_n780,
         dp_id_stage_regfile_DataPath_Physical_RF_n779,
         dp_id_stage_regfile_DataPath_Physical_RF_n778,
         dp_id_stage_regfile_DataPath_Physical_RF_n777,
         dp_id_stage_regfile_DataPath_Physical_RF_n776,
         dp_id_stage_regfile_DataPath_Physical_RF_n775,
         dp_id_stage_regfile_DataPath_Physical_RF_n774,
         dp_id_stage_regfile_DataPath_Physical_RF_n773,
         dp_id_stage_regfile_DataPath_Physical_RF_n772,
         dp_id_stage_regfile_DataPath_Physical_RF_n771,
         dp_id_stage_regfile_DataPath_Physical_RF_n770,
         dp_id_stage_regfile_DataPath_Physical_RF_n769,
         dp_id_stage_regfile_DataPath_Physical_RF_n768,
         dp_id_stage_regfile_DataPath_Physical_RF_n767,
         dp_id_stage_regfile_DataPath_Physical_RF_n766,
         dp_id_stage_regfile_DataPath_Physical_RF_n765,
         dp_id_stage_regfile_DataPath_Physical_RF_n764,
         dp_id_stage_regfile_DataPath_Physical_RF_n763,
         dp_id_stage_regfile_DataPath_Physical_RF_n762,
         dp_id_stage_regfile_DataPath_Physical_RF_n761,
         dp_id_stage_regfile_DataPath_Physical_RF_n760,
         dp_id_stage_regfile_DataPath_Physical_RF_n759,
         dp_id_stage_regfile_DataPath_Physical_RF_n758,
         dp_id_stage_regfile_DataPath_Physical_RF_n757,
         dp_id_stage_regfile_DataPath_Physical_RF_n756,
         dp_id_stage_regfile_DataPath_Physical_RF_n755,
         dp_id_stage_regfile_DataPath_Physical_RF_n754,
         dp_id_stage_regfile_DataPath_Physical_RF_n753,
         dp_id_stage_regfile_DataPath_Physical_RF_n752,
         dp_id_stage_regfile_DataPath_Physical_RF_n751,
         dp_id_stage_regfile_DataPath_Physical_RF_n750,
         dp_id_stage_regfile_DataPath_Physical_RF_n749,
         dp_id_stage_regfile_DataPath_Physical_RF_n748,
         dp_id_stage_regfile_DataPath_Physical_RF_n747,
         dp_id_stage_regfile_DataPath_Physical_RF_n746,
         dp_id_stage_regfile_DataPath_Physical_RF_n745,
         dp_id_stage_regfile_DataPath_Physical_RF_n744,
         dp_id_stage_regfile_DataPath_Physical_RF_n743,
         dp_id_stage_regfile_DataPath_Physical_RF_n742,
         dp_id_stage_regfile_DataPath_Physical_RF_n741,
         dp_id_stage_regfile_DataPath_Physical_RF_n740,
         dp_id_stage_regfile_DataPath_Physical_RF_n739,
         dp_id_stage_regfile_DataPath_Physical_RF_n738,
         dp_id_stage_regfile_DataPath_Physical_RF_n737,
         dp_id_stage_regfile_DataPath_Physical_RF_n736,
         dp_id_stage_regfile_DataPath_Physical_RF_n735,
         dp_id_stage_regfile_DataPath_Physical_RF_n734,
         dp_id_stage_regfile_DataPath_Physical_RF_n733,
         dp_id_stage_regfile_DataPath_Physical_RF_n732,
         dp_id_stage_regfile_DataPath_Physical_RF_n731,
         dp_id_stage_regfile_DataPath_Physical_RF_n730,
         dp_id_stage_regfile_DataPath_Physical_RF_n729,
         dp_id_stage_regfile_DataPath_Physical_RF_n728,
         dp_id_stage_regfile_DataPath_Physical_RF_n727,
         dp_id_stage_regfile_DataPath_Physical_RF_n726,
         dp_id_stage_regfile_DataPath_Physical_RF_n725,
         dp_id_stage_regfile_DataPath_Physical_RF_n724,
         dp_id_stage_regfile_DataPath_Physical_RF_n723,
         dp_id_stage_regfile_DataPath_Physical_RF_n722,
         dp_id_stage_regfile_DataPath_Physical_RF_n721,
         dp_id_stage_regfile_DataPath_Physical_RF_n720,
         dp_id_stage_regfile_DataPath_Physical_RF_n719,
         dp_id_stage_regfile_DataPath_Physical_RF_n718,
         dp_id_stage_regfile_DataPath_Physical_RF_n717,
         dp_id_stage_regfile_DataPath_Physical_RF_n716,
         dp_id_stage_regfile_DataPath_Physical_RF_n715,
         dp_id_stage_regfile_DataPath_Physical_RF_n714,
         dp_id_stage_regfile_DataPath_Physical_RF_n713,
         dp_id_stage_regfile_DataPath_Physical_RF_n712,
         dp_id_stage_regfile_DataPath_Physical_RF_n711,
         dp_id_stage_regfile_DataPath_Physical_RF_n710,
         dp_id_stage_regfile_DataPath_Physical_RF_n709,
         dp_id_stage_regfile_DataPath_Physical_RF_n708,
         dp_id_stage_regfile_DataPath_Physical_RF_n707,
         dp_id_stage_regfile_DataPath_Physical_RF_n706,
         dp_id_stage_regfile_DataPath_Physical_RF_n705,
         dp_id_stage_regfile_DataPath_Physical_RF_n704,
         dp_id_stage_regfile_DataPath_Physical_RF_n703,
         dp_id_stage_regfile_DataPath_Physical_RF_n702,
         dp_id_stage_regfile_DataPath_Physical_RF_n701,
         dp_id_stage_regfile_DataPath_Physical_RF_n700,
         dp_id_stage_regfile_DataPath_Physical_RF_n699,
         dp_id_stage_regfile_DataPath_Physical_RF_n698,
         dp_id_stage_regfile_DataPath_Physical_RF_n697,
         dp_id_stage_regfile_DataPath_Physical_RF_n696,
         dp_id_stage_regfile_DataPath_Physical_RF_n695,
         dp_id_stage_regfile_DataPath_Physical_RF_n694,
         dp_id_stage_regfile_DataPath_Physical_RF_n693,
         dp_id_stage_regfile_DataPath_Physical_RF_n692,
         dp_id_stage_regfile_DataPath_Physical_RF_n691,
         dp_id_stage_regfile_DataPath_Physical_RF_n690,
         dp_id_stage_regfile_DataPath_Physical_RF_n689,
         dp_id_stage_regfile_DataPath_Physical_RF_n688,
         dp_id_stage_regfile_DataPath_Physical_RF_n687,
         dp_id_stage_regfile_DataPath_Physical_RF_n686,
         dp_id_stage_regfile_DataPath_Physical_RF_n685,
         dp_id_stage_regfile_DataPath_Physical_RF_n684,
         dp_id_stage_regfile_DataPath_Physical_RF_n683,
         dp_id_stage_regfile_DataPath_Physical_RF_n682,
         dp_id_stage_regfile_DataPath_Physical_RF_n681,
         dp_id_stage_regfile_DataPath_Physical_RF_n680,
         dp_id_stage_regfile_DataPath_Physical_RF_n679,
         dp_id_stage_regfile_DataPath_Physical_RF_n678,
         dp_id_stage_regfile_DataPath_Physical_RF_n677,
         dp_id_stage_regfile_DataPath_Physical_RF_n676,
         dp_id_stage_regfile_DataPath_Physical_RF_n675,
         dp_id_stage_regfile_DataPath_Physical_RF_n674,
         dp_id_stage_regfile_DataPath_Physical_RF_n673,
         dp_id_stage_regfile_DataPath_Physical_RF_n672,
         dp_id_stage_regfile_DataPath_Physical_RF_n671,
         dp_id_stage_regfile_DataPath_Physical_RF_n670,
         dp_id_stage_regfile_DataPath_Physical_RF_n669,
         dp_id_stage_regfile_DataPath_Physical_RF_n668,
         dp_id_stage_regfile_DataPath_Physical_RF_n667,
         dp_id_stage_regfile_DataPath_Physical_RF_n666,
         dp_id_stage_regfile_DataPath_Physical_RF_n665,
         dp_id_stage_regfile_DataPath_Physical_RF_n664,
         dp_id_stage_regfile_DataPath_Physical_RF_n663,
         dp_id_stage_regfile_DataPath_Physical_RF_n662,
         dp_id_stage_regfile_DataPath_Physical_RF_n661,
         dp_id_stage_regfile_DataPath_Physical_RF_n660,
         dp_id_stage_regfile_DataPath_Physical_RF_n659,
         dp_id_stage_regfile_DataPath_Physical_RF_n658,
         dp_id_stage_regfile_DataPath_Physical_RF_n657,
         dp_id_stage_regfile_DataPath_Physical_RF_n656,
         dp_id_stage_regfile_DataPath_Physical_RF_n655,
         dp_id_stage_regfile_DataPath_Physical_RF_n654,
         dp_id_stage_regfile_DataPath_Physical_RF_n653,
         dp_id_stage_regfile_DataPath_Physical_RF_n652,
         dp_id_stage_regfile_DataPath_Physical_RF_n651,
         dp_id_stage_regfile_DataPath_Physical_RF_n650,
         dp_id_stage_regfile_DataPath_Physical_RF_n649,
         dp_id_stage_regfile_DataPath_Physical_RF_n648,
         dp_id_stage_regfile_DataPath_Physical_RF_n647,
         dp_id_stage_regfile_DataPath_Physical_RF_n646,
         dp_id_stage_regfile_DataPath_Physical_RF_n645,
         dp_id_stage_regfile_DataPath_Physical_RF_n644,
         dp_id_stage_regfile_DataPath_Physical_RF_n643,
         dp_id_stage_regfile_DataPath_Physical_RF_n642,
         dp_id_stage_regfile_DataPath_Physical_RF_n641,
         dp_id_stage_regfile_DataPath_Physical_RF_n640,
         dp_id_stage_regfile_DataPath_Physical_RF_n639,
         dp_id_stage_regfile_DataPath_Physical_RF_n638,
         dp_id_stage_regfile_DataPath_Physical_RF_n637,
         dp_id_stage_regfile_DataPath_Physical_RF_n636,
         dp_id_stage_regfile_DataPath_Physical_RF_n635,
         dp_id_stage_regfile_DataPath_Physical_RF_n634,
         dp_id_stage_regfile_DataPath_Physical_RF_n633,
         dp_id_stage_regfile_DataPath_Physical_RF_n632,
         dp_id_stage_regfile_DataPath_Physical_RF_n631,
         dp_id_stage_regfile_DataPath_Physical_RF_n630,
         dp_id_stage_regfile_DataPath_Physical_RF_n629,
         dp_id_stage_regfile_DataPath_Physical_RF_n628,
         dp_id_stage_regfile_DataPath_Physical_RF_n627,
         dp_id_stage_regfile_DataPath_Physical_RF_n626,
         dp_id_stage_regfile_DataPath_Physical_RF_n625,
         dp_id_stage_regfile_DataPath_Physical_RF_n624,
         dp_id_stage_regfile_DataPath_Physical_RF_n623,
         dp_id_stage_regfile_DataPath_Physical_RF_n622,
         dp_id_stage_regfile_DataPath_Physical_RF_n621,
         dp_id_stage_regfile_DataPath_Physical_RF_n620,
         dp_id_stage_regfile_DataPath_Physical_RF_n619,
         dp_id_stage_regfile_DataPath_Physical_RF_n618,
         dp_id_stage_regfile_DataPath_Physical_RF_n617,
         dp_id_stage_regfile_DataPath_Physical_RF_n616,
         dp_id_stage_regfile_DataPath_Physical_RF_n615,
         dp_id_stage_regfile_DataPath_Physical_RF_n614,
         dp_id_stage_regfile_DataPath_Physical_RF_n613,
         dp_id_stage_regfile_DataPath_Physical_RF_n612,
         dp_id_stage_regfile_DataPath_Physical_RF_n611,
         dp_id_stage_regfile_DataPath_Physical_RF_n610,
         dp_id_stage_regfile_DataPath_Physical_RF_n609,
         dp_id_stage_regfile_DataPath_Physical_RF_n608,
         dp_id_stage_regfile_DataPath_Physical_RF_n607,
         dp_id_stage_regfile_DataPath_Physical_RF_n606,
         dp_id_stage_regfile_DataPath_Physical_RF_n605,
         dp_id_stage_regfile_DataPath_Physical_RF_n604,
         dp_id_stage_regfile_DataPath_Physical_RF_n603,
         dp_id_stage_regfile_DataPath_Physical_RF_n602,
         dp_id_stage_regfile_DataPath_Physical_RF_n601,
         dp_id_stage_regfile_DataPath_Physical_RF_n600,
         dp_id_stage_regfile_DataPath_Physical_RF_n599,
         dp_id_stage_regfile_DataPath_Physical_RF_n598,
         dp_id_stage_regfile_DataPath_Physical_RF_n597,
         dp_id_stage_regfile_DataPath_Physical_RF_n596,
         dp_id_stage_regfile_DataPath_Physical_RF_n595,
         dp_id_stage_regfile_DataPath_Physical_RF_n594,
         dp_id_stage_regfile_DataPath_Physical_RF_n593,
         dp_id_stage_regfile_DataPath_Physical_RF_n592,
         dp_id_stage_regfile_DataPath_Physical_RF_n591,
         dp_id_stage_regfile_DataPath_Physical_RF_n590,
         dp_id_stage_regfile_DataPath_Physical_RF_n589,
         dp_id_stage_regfile_DataPath_Physical_RF_n588,
         dp_id_stage_regfile_DataPath_Physical_RF_n587,
         dp_id_stage_regfile_DataPath_Physical_RF_n586,
         dp_id_stage_regfile_DataPath_Physical_RF_n585,
         dp_id_stage_regfile_DataPath_Physical_RF_n584,
         dp_id_stage_regfile_DataPath_Physical_RF_n583,
         dp_id_stage_regfile_DataPath_Physical_RF_n582,
         dp_id_stage_regfile_DataPath_Physical_RF_n581,
         dp_id_stage_regfile_DataPath_Physical_RF_n580,
         dp_id_stage_regfile_DataPath_Physical_RF_n579,
         dp_id_stage_regfile_DataPath_Physical_RF_n578,
         dp_id_stage_regfile_DataPath_Physical_RF_n577,
         dp_id_stage_regfile_DataPath_Physical_RF_n576,
         dp_id_stage_regfile_DataPath_Physical_RF_n575,
         dp_id_stage_regfile_DataPath_Physical_RF_n574,
         dp_id_stage_regfile_DataPath_Physical_RF_n573,
         dp_id_stage_regfile_DataPath_Physical_RF_n572,
         dp_id_stage_regfile_DataPath_Physical_RF_n571,
         dp_id_stage_regfile_DataPath_Physical_RF_n570,
         dp_id_stage_regfile_DataPath_Physical_RF_n569,
         dp_id_stage_regfile_DataPath_Physical_RF_n568,
         dp_id_stage_regfile_DataPath_Physical_RF_n567,
         dp_id_stage_regfile_DataPath_Physical_RF_n566,
         dp_id_stage_regfile_DataPath_Physical_RF_n565,
         dp_id_stage_regfile_DataPath_Physical_RF_n564,
         dp_id_stage_regfile_DataPath_Physical_RF_n563,
         dp_id_stage_regfile_DataPath_Physical_RF_n562,
         dp_id_stage_regfile_DataPath_Physical_RF_n561,
         dp_id_stage_regfile_DataPath_Physical_RF_n560,
         dp_id_stage_regfile_DataPath_Physical_RF_n559,
         dp_id_stage_regfile_DataPath_Physical_RF_n558,
         dp_id_stage_regfile_DataPath_Physical_RF_n557,
         dp_id_stage_regfile_DataPath_Physical_RF_n556,
         dp_id_stage_regfile_DataPath_Physical_RF_n555,
         dp_id_stage_regfile_DataPath_Physical_RF_n554,
         dp_id_stage_regfile_DataPath_Physical_RF_n553,
         dp_id_stage_regfile_DataPath_Physical_RF_n552,
         dp_id_stage_regfile_DataPath_Physical_RF_n551,
         dp_id_stage_regfile_DataPath_Physical_RF_n550,
         dp_id_stage_regfile_DataPath_Physical_RF_n549,
         dp_id_stage_regfile_DataPath_Physical_RF_n548,
         dp_id_stage_regfile_DataPath_Physical_RF_n547,
         dp_id_stage_regfile_DataPath_Physical_RF_n546,
         dp_id_stage_regfile_DataPath_Physical_RF_n545,
         dp_id_stage_regfile_DataPath_Physical_RF_n544,
         dp_id_stage_regfile_DataPath_Physical_RF_n543,
         dp_id_stage_regfile_DataPath_Physical_RF_n542,
         dp_id_stage_regfile_DataPath_Physical_RF_n541,
         dp_id_stage_regfile_DataPath_Physical_RF_n540,
         dp_id_stage_regfile_DataPath_Physical_RF_n539,
         dp_id_stage_regfile_DataPath_Physical_RF_n538,
         dp_id_stage_regfile_DataPath_Physical_RF_n537,
         dp_id_stage_regfile_DataPath_Physical_RF_n536,
         dp_id_stage_regfile_DataPath_Physical_RF_n535,
         dp_id_stage_regfile_DataPath_Physical_RF_n534,
         dp_id_stage_regfile_DataPath_Physical_RF_n533,
         dp_id_stage_regfile_DataPath_Physical_RF_n532,
         dp_id_stage_regfile_DataPath_Physical_RF_n531,
         dp_id_stage_regfile_DataPath_Physical_RF_n530,
         dp_id_stage_regfile_DataPath_Physical_RF_n529,
         dp_id_stage_regfile_DataPath_Physical_RF_n528,
         dp_id_stage_regfile_DataPath_Physical_RF_n527,
         dp_id_stage_regfile_DataPath_Physical_RF_n526,
         dp_id_stage_regfile_DataPath_Physical_RF_n525,
         dp_id_stage_regfile_DataPath_Physical_RF_n524,
         dp_id_stage_regfile_DataPath_Physical_RF_n523,
         dp_id_stage_regfile_DataPath_Physical_RF_n522,
         dp_id_stage_regfile_DataPath_Physical_RF_n521,
         dp_id_stage_regfile_DataPath_Physical_RF_n520,
         dp_id_stage_regfile_DataPath_Physical_RF_n519,
         dp_id_stage_regfile_DataPath_Physical_RF_n518,
         dp_id_stage_regfile_DataPath_Physical_RF_n517,
         dp_id_stage_regfile_DataPath_Physical_RF_n516,
         dp_id_stage_regfile_DataPath_Physical_RF_n515,
         dp_id_stage_regfile_DataPath_Physical_RF_n514,
         dp_id_stage_regfile_DataPath_Physical_RF_n513,
         dp_id_stage_regfile_DataPath_Physical_RF_n512,
         dp_id_stage_regfile_DataPath_Physical_RF_n511,
         dp_id_stage_regfile_DataPath_Physical_RF_n510,
         dp_id_stage_regfile_DataPath_Physical_RF_n509,
         dp_id_stage_regfile_DataPath_Physical_RF_n508,
         dp_id_stage_regfile_DataPath_Physical_RF_n507,
         dp_id_stage_regfile_DataPath_Physical_RF_n506,
         dp_id_stage_regfile_DataPath_Physical_RF_n505,
         dp_id_stage_regfile_DataPath_Physical_RF_n504,
         dp_id_stage_regfile_DataPath_Physical_RF_n503,
         dp_id_stage_regfile_DataPath_Physical_RF_n502,
         dp_id_stage_regfile_DataPath_Physical_RF_n501,
         dp_id_stage_regfile_DataPath_Physical_RF_n500,
         dp_id_stage_regfile_DataPath_Physical_RF_n499,
         dp_id_stage_regfile_DataPath_Physical_RF_n498,
         dp_id_stage_regfile_DataPath_Physical_RF_n497,
         dp_id_stage_regfile_DataPath_Physical_RF_n496,
         dp_id_stage_regfile_DataPath_Physical_RF_n495,
         dp_id_stage_regfile_DataPath_Physical_RF_n494,
         dp_id_stage_regfile_DataPath_Physical_RF_n493,
         dp_id_stage_regfile_DataPath_Physical_RF_n492,
         dp_id_stage_regfile_DataPath_Physical_RF_n491,
         dp_id_stage_regfile_DataPath_Physical_RF_n490,
         dp_id_stage_regfile_DataPath_Physical_RF_n489,
         dp_id_stage_regfile_DataPath_Physical_RF_n488,
         dp_id_stage_regfile_DataPath_Physical_RF_n487,
         dp_id_stage_regfile_DataPath_Physical_RF_n486,
         dp_id_stage_regfile_DataPath_Physical_RF_n485,
         dp_id_stage_regfile_DataPath_Physical_RF_n484,
         dp_id_stage_regfile_DataPath_Physical_RF_n483,
         dp_id_stage_regfile_DataPath_Physical_RF_n482,
         dp_id_stage_regfile_DataPath_Physical_RF_n481,
         dp_id_stage_regfile_DataPath_Physical_RF_n480,
         dp_id_stage_regfile_DataPath_Physical_RF_n479,
         dp_id_stage_regfile_DataPath_Physical_RF_n478,
         dp_id_stage_regfile_DataPath_Physical_RF_n477,
         dp_id_stage_regfile_DataPath_Physical_RF_n476,
         dp_id_stage_regfile_DataPath_Physical_RF_n475,
         dp_id_stage_regfile_DataPath_Physical_RF_n474,
         dp_id_stage_regfile_DataPath_Physical_RF_n473,
         dp_id_stage_regfile_DataPath_Physical_RF_n472,
         dp_id_stage_regfile_DataPath_Physical_RF_n471,
         dp_id_stage_regfile_DataPath_Physical_RF_n470,
         dp_id_stage_regfile_DataPath_Physical_RF_n469,
         dp_id_stage_regfile_DataPath_Physical_RF_n468,
         dp_id_stage_regfile_DataPath_Physical_RF_n467,
         dp_id_stage_regfile_DataPath_Physical_RF_n466,
         dp_id_stage_regfile_DataPath_Physical_RF_n465,
         dp_id_stage_regfile_DataPath_Physical_RF_n464,
         dp_id_stage_regfile_DataPath_Physical_RF_n463,
         dp_id_stage_regfile_DataPath_Physical_RF_n462,
         dp_id_stage_regfile_DataPath_Physical_RF_n461,
         dp_id_stage_regfile_DataPath_Physical_RF_n460,
         dp_id_stage_regfile_DataPath_Physical_RF_n459,
         dp_id_stage_regfile_DataPath_Physical_RF_n458,
         dp_id_stage_regfile_DataPath_Physical_RF_n457,
         dp_id_stage_regfile_DataPath_Physical_RF_n456,
         dp_id_stage_regfile_DataPath_Physical_RF_n455,
         dp_id_stage_regfile_DataPath_Physical_RF_n454,
         dp_id_stage_regfile_DataPath_Physical_RF_n453,
         dp_id_stage_regfile_DataPath_Physical_RF_n452,
         dp_id_stage_regfile_DataPath_Physical_RF_n451,
         dp_id_stage_regfile_DataPath_Physical_RF_n450,
         dp_id_stage_regfile_DataPath_Physical_RF_n449,
         dp_id_stage_regfile_DataPath_Physical_RF_n448,
         dp_id_stage_regfile_DataPath_Physical_RF_n447,
         dp_id_stage_regfile_DataPath_Physical_RF_n446,
         dp_id_stage_regfile_DataPath_Physical_RF_n445,
         dp_id_stage_regfile_DataPath_Physical_RF_n444,
         dp_id_stage_regfile_DataPath_Physical_RF_n443,
         dp_id_stage_regfile_DataPath_Physical_RF_n442,
         dp_id_stage_regfile_DataPath_Physical_RF_n441,
         dp_id_stage_regfile_DataPath_Physical_RF_n440,
         dp_id_stage_regfile_DataPath_Physical_RF_n439,
         dp_id_stage_regfile_DataPath_Physical_RF_n438,
         dp_id_stage_regfile_DataPath_Physical_RF_n437,
         dp_id_stage_regfile_DataPath_Physical_RF_n436,
         dp_id_stage_regfile_DataPath_Physical_RF_n435,
         dp_id_stage_regfile_DataPath_Physical_RF_n434,
         dp_id_stage_regfile_DataPath_Physical_RF_n433,
         dp_id_stage_regfile_DataPath_Physical_RF_n432,
         dp_id_stage_regfile_DataPath_Physical_RF_n431,
         dp_id_stage_regfile_DataPath_Physical_RF_n430,
         dp_id_stage_regfile_DataPath_Physical_RF_n429,
         dp_id_stage_regfile_DataPath_Physical_RF_n428,
         dp_id_stage_regfile_DataPath_Physical_RF_n427,
         dp_id_stage_regfile_DataPath_Physical_RF_n426,
         dp_id_stage_regfile_DataPath_Physical_RF_n425,
         dp_id_stage_regfile_DataPath_Physical_RF_n424,
         dp_id_stage_regfile_DataPath_Physical_RF_n423,
         dp_id_stage_regfile_DataPath_Physical_RF_n422,
         dp_id_stage_regfile_DataPath_Physical_RF_n421,
         dp_id_stage_regfile_DataPath_Physical_RF_n420,
         dp_id_stage_regfile_DataPath_Physical_RF_n419,
         dp_id_stage_regfile_DataPath_Physical_RF_n418,
         dp_id_stage_regfile_DataPath_Physical_RF_n417,
         dp_id_stage_regfile_DataPath_Physical_RF_n416,
         dp_id_stage_regfile_DataPath_Physical_RF_n415,
         dp_id_stage_regfile_DataPath_Physical_RF_n414,
         dp_id_stage_regfile_DataPath_Physical_RF_n413,
         dp_id_stage_regfile_DataPath_Physical_RF_n412,
         dp_id_stage_regfile_DataPath_Physical_RF_n411,
         dp_id_stage_regfile_DataPath_Physical_RF_n410,
         dp_id_stage_regfile_DataPath_Physical_RF_n409,
         dp_id_stage_regfile_DataPath_Physical_RF_n408,
         dp_id_stage_regfile_DataPath_Physical_RF_n407,
         dp_id_stage_regfile_DataPath_Physical_RF_n406,
         dp_id_stage_regfile_DataPath_Physical_RF_n405,
         dp_id_stage_regfile_DataPath_Physical_RF_n404,
         dp_id_stage_regfile_DataPath_Physical_RF_n403,
         dp_id_stage_regfile_DataPath_Physical_RF_n402,
         dp_id_stage_regfile_DataPath_Physical_RF_n401,
         dp_id_stage_regfile_DataPath_Physical_RF_n400,
         dp_id_stage_regfile_DataPath_Physical_RF_n399,
         dp_id_stage_regfile_DataPath_Physical_RF_n398,
         dp_id_stage_regfile_DataPath_Physical_RF_n397,
         dp_id_stage_regfile_DataPath_Physical_RF_n396,
         dp_id_stage_regfile_DataPath_Physical_RF_n395,
         dp_id_stage_regfile_DataPath_Physical_RF_n394,
         dp_id_stage_regfile_DataPath_Physical_RF_n393,
         dp_id_stage_regfile_DataPath_Physical_RF_n392,
         dp_id_stage_regfile_DataPath_Physical_RF_n391,
         dp_id_stage_regfile_DataPath_Physical_RF_n390,
         dp_id_stage_regfile_DataPath_Physical_RF_n389,
         dp_id_stage_regfile_DataPath_Physical_RF_n388,
         dp_id_stage_regfile_DataPath_Physical_RF_n387,
         dp_id_stage_regfile_DataPath_Physical_RF_n386,
         dp_id_stage_regfile_DataPath_Physical_RF_n385,
         dp_id_stage_regfile_DataPath_Physical_RF_n384,
         dp_id_stage_regfile_DataPath_Physical_RF_n383,
         dp_id_stage_regfile_DataPath_Physical_RF_n382,
         dp_id_stage_regfile_DataPath_Physical_RF_n381,
         dp_id_stage_regfile_DataPath_Physical_RF_n380,
         dp_id_stage_regfile_DataPath_Physical_RF_n379,
         dp_id_stage_regfile_DataPath_Physical_RF_n378,
         dp_id_stage_regfile_DataPath_Physical_RF_n377,
         dp_id_stage_regfile_DataPath_Physical_RF_n376,
         dp_id_stage_regfile_DataPath_Physical_RF_n375,
         dp_id_stage_regfile_DataPath_Physical_RF_n374,
         dp_id_stage_regfile_DataPath_Physical_RF_n373,
         dp_id_stage_regfile_DataPath_Physical_RF_n372,
         dp_id_stage_regfile_DataPath_Physical_RF_n371,
         dp_id_stage_regfile_DataPath_Physical_RF_n370,
         dp_id_stage_regfile_DataPath_Physical_RF_n369,
         dp_id_stage_regfile_DataPath_Physical_RF_n368,
         dp_id_stage_regfile_DataPath_Physical_RF_n367,
         dp_id_stage_regfile_DataPath_Physical_RF_n366,
         dp_id_stage_regfile_DataPath_Physical_RF_n365,
         dp_id_stage_regfile_DataPath_Physical_RF_n364,
         dp_id_stage_regfile_DataPath_Physical_RF_n363,
         dp_id_stage_regfile_DataPath_Physical_RF_n362,
         dp_id_stage_regfile_DataPath_Physical_RF_n361,
         dp_id_stage_regfile_DataPath_Physical_RF_n360,
         dp_id_stage_regfile_DataPath_Physical_RF_n359,
         dp_id_stage_regfile_DataPath_Physical_RF_n358,
         dp_id_stage_regfile_DataPath_Physical_RF_n357,
         dp_id_stage_regfile_DataPath_Physical_RF_n356,
         dp_id_stage_regfile_DataPath_Physical_RF_n355,
         dp_id_stage_regfile_DataPath_Physical_RF_n354,
         dp_id_stage_regfile_DataPath_Physical_RF_n353,
         dp_id_stage_regfile_DataPath_Physical_RF_n352,
         dp_id_stage_regfile_DataPath_Physical_RF_n351,
         dp_id_stage_regfile_DataPath_Physical_RF_n350,
         dp_id_stage_regfile_DataPath_Physical_RF_n349,
         dp_id_stage_regfile_DataPath_Physical_RF_n348,
         dp_id_stage_regfile_DataPath_Physical_RF_n347,
         dp_id_stage_regfile_DataPath_Physical_RF_n346,
         dp_id_stage_regfile_DataPath_Physical_RF_n345,
         dp_id_stage_regfile_DataPath_Physical_RF_n344,
         dp_id_stage_regfile_DataPath_Physical_RF_n343,
         dp_id_stage_regfile_DataPath_Physical_RF_n342,
         dp_id_stage_regfile_DataPath_Physical_RF_n341,
         dp_id_stage_regfile_DataPath_Physical_RF_n340,
         dp_id_stage_regfile_DataPath_Physical_RF_n339,
         dp_id_stage_regfile_DataPath_Physical_RF_n338,
         dp_id_stage_regfile_DataPath_Physical_RF_n337,
         dp_id_stage_regfile_DataPath_Physical_RF_n336,
         dp_id_stage_regfile_DataPath_Physical_RF_n335,
         dp_id_stage_regfile_DataPath_Physical_RF_n334,
         dp_id_stage_regfile_DataPath_Physical_RF_n333,
         dp_id_stage_regfile_DataPath_Physical_RF_n332,
         dp_id_stage_regfile_DataPath_Physical_RF_n331,
         dp_id_stage_regfile_DataPath_Physical_RF_n330,
         dp_id_stage_regfile_DataPath_Physical_RF_n329,
         dp_id_stage_regfile_DataPath_Physical_RF_n328,
         dp_id_stage_regfile_DataPath_Physical_RF_n327,
         dp_id_stage_regfile_DataPath_Physical_RF_n326,
         dp_id_stage_regfile_DataPath_Physical_RF_n325,
         dp_id_stage_regfile_DataPath_Physical_RF_n324,
         dp_id_stage_regfile_DataPath_Physical_RF_n323,
         dp_id_stage_regfile_DataPath_Physical_RF_n322,
         dp_id_stage_regfile_DataPath_Physical_RF_n321,
         dp_id_stage_regfile_DataPath_Physical_RF_n320,
         dp_id_stage_regfile_DataPath_Physical_RF_n319,
         dp_id_stage_regfile_DataPath_Physical_RF_n318,
         dp_id_stage_regfile_DataPath_Physical_RF_n317,
         dp_id_stage_regfile_DataPath_Physical_RF_n316,
         dp_id_stage_regfile_DataPath_Physical_RF_n315,
         dp_id_stage_regfile_DataPath_Physical_RF_n314,
         dp_id_stage_regfile_DataPath_Physical_RF_n313,
         dp_id_stage_regfile_DataPath_Physical_RF_n312,
         dp_id_stage_regfile_DataPath_Physical_RF_n311,
         dp_id_stage_regfile_DataPath_Physical_RF_n310,
         dp_id_stage_regfile_DataPath_Physical_RF_n309,
         dp_id_stage_regfile_DataPath_Physical_RF_n308,
         dp_id_stage_regfile_DataPath_Physical_RF_n307,
         dp_id_stage_regfile_DataPath_Physical_RF_n306,
         dp_id_stage_regfile_DataPath_Physical_RF_n305,
         dp_id_stage_regfile_DataPath_Physical_RF_n304,
         dp_id_stage_regfile_DataPath_Physical_RF_n303,
         dp_id_stage_regfile_DataPath_Physical_RF_n302,
         dp_id_stage_regfile_DataPath_Physical_RF_n301,
         dp_id_stage_regfile_DataPath_Physical_RF_n300,
         dp_id_stage_regfile_DataPath_Physical_RF_n299,
         dp_id_stage_regfile_DataPath_Physical_RF_n298,
         dp_id_stage_regfile_DataPath_Physical_RF_n297,
         dp_id_stage_regfile_DataPath_Physical_RF_n296,
         dp_id_stage_regfile_DataPath_Physical_RF_n295,
         dp_id_stage_regfile_DataPath_Physical_RF_n294,
         dp_id_stage_regfile_DataPath_Physical_RF_n293,
         dp_id_stage_regfile_DataPath_Physical_RF_n292,
         dp_id_stage_regfile_DataPath_Physical_RF_n291,
         dp_id_stage_regfile_DataPath_Physical_RF_n290,
         dp_id_stage_regfile_DataPath_Physical_RF_n289,
         dp_id_stage_regfile_DataPath_Physical_RF_n288,
         dp_id_stage_regfile_DataPath_Physical_RF_n287,
         dp_id_stage_regfile_DataPath_Physical_RF_n286,
         dp_id_stage_regfile_DataPath_Physical_RF_n285,
         dp_id_stage_regfile_DataPath_Physical_RF_n284,
         dp_id_stage_regfile_DataPath_Physical_RF_n283,
         dp_id_stage_regfile_DataPath_Physical_RF_n282,
         dp_id_stage_regfile_DataPath_Physical_RF_n281,
         dp_id_stage_regfile_DataPath_Physical_RF_n280,
         dp_id_stage_regfile_DataPath_Physical_RF_n279,
         dp_id_stage_regfile_DataPath_Physical_RF_n278,
         dp_id_stage_regfile_DataPath_Physical_RF_n277,
         dp_id_stage_regfile_DataPath_Physical_RF_n276,
         dp_id_stage_regfile_DataPath_Physical_RF_n275,
         dp_id_stage_regfile_DataPath_Physical_RF_n274,
         dp_id_stage_regfile_DataPath_Physical_RF_n273,
         dp_id_stage_regfile_DataPath_Physical_RF_n272,
         dp_id_stage_regfile_DataPath_Physical_RF_n271,
         dp_id_stage_regfile_DataPath_Physical_RF_n270,
         dp_id_stage_regfile_DataPath_Physical_RF_n269,
         dp_id_stage_regfile_DataPath_Physical_RF_n268,
         dp_id_stage_regfile_DataPath_Physical_RF_n267,
         dp_id_stage_regfile_DataPath_Physical_RF_n266,
         dp_id_stage_regfile_DataPath_Physical_RF_n265,
         dp_id_stage_regfile_DataPath_Physical_RF_n264,
         dp_id_stage_regfile_DataPath_Physical_RF_n263,
         dp_id_stage_regfile_DataPath_Physical_RF_n262,
         dp_id_stage_regfile_DataPath_Physical_RF_n261,
         dp_id_stage_regfile_DataPath_Physical_RF_n260,
         dp_id_stage_regfile_DataPath_Physical_RF_n259,
         dp_id_stage_regfile_DataPath_Physical_RF_n258,
         dp_id_stage_regfile_DataPath_Physical_RF_n257,
         dp_id_stage_regfile_DataPath_Physical_RF_n256,
         dp_id_stage_regfile_DataPath_Physical_RF_n255,
         dp_id_stage_regfile_DataPath_Physical_RF_n254,
         dp_id_stage_regfile_DataPath_Physical_RF_n253,
         dp_id_stage_regfile_DataPath_Physical_RF_n252,
         dp_id_stage_regfile_DataPath_Physical_RF_n251,
         dp_id_stage_regfile_DataPath_Physical_RF_n250,
         dp_id_stage_regfile_DataPath_Physical_RF_n249,
         dp_id_stage_regfile_DataPath_Physical_RF_n248,
         dp_id_stage_regfile_DataPath_Physical_RF_n247,
         dp_id_stage_regfile_DataPath_Physical_RF_n246,
         dp_id_stage_regfile_DataPath_Physical_RF_n245,
         dp_id_stage_regfile_DataPath_Physical_RF_n244,
         dp_id_stage_regfile_DataPath_Physical_RF_n243,
         dp_id_stage_regfile_DataPath_Physical_RF_n242,
         dp_id_stage_regfile_DataPath_Physical_RF_n241,
         dp_id_stage_regfile_DataPath_Physical_RF_n240,
         dp_id_stage_regfile_DataPath_Physical_RF_n239,
         dp_id_stage_regfile_DataPath_Physical_RF_n238,
         dp_id_stage_regfile_DataPath_Physical_RF_n237,
         dp_id_stage_regfile_DataPath_Physical_RF_n236,
         dp_id_stage_regfile_DataPath_Physical_RF_n235,
         dp_id_stage_regfile_DataPath_Physical_RF_n234,
         dp_id_stage_regfile_DataPath_Physical_RF_n233,
         dp_id_stage_regfile_DataPath_Physical_RF_n232,
         dp_id_stage_regfile_DataPath_Physical_RF_n231,
         dp_id_stage_regfile_DataPath_Physical_RF_n230,
         dp_id_stage_regfile_DataPath_Physical_RF_n229,
         dp_id_stage_regfile_DataPath_Physical_RF_n228,
         dp_id_stage_regfile_DataPath_Physical_RF_n227,
         dp_id_stage_regfile_DataPath_Physical_RF_n226,
         dp_id_stage_regfile_DataPath_Physical_RF_n225,
         dp_id_stage_regfile_DataPath_Physical_RF_n224,
         dp_id_stage_regfile_DataPath_Physical_RF_n223,
         dp_id_stage_regfile_DataPath_Physical_RF_n222,
         dp_id_stage_regfile_DataPath_Physical_RF_n221,
         dp_id_stage_regfile_DataPath_Physical_RF_n220,
         dp_id_stage_regfile_DataPath_Physical_RF_n219,
         dp_id_stage_regfile_DataPath_Physical_RF_n218,
         dp_id_stage_regfile_DataPath_Physical_RF_n217,
         dp_id_stage_regfile_DataPath_Physical_RF_n216,
         dp_id_stage_regfile_DataPath_Physical_RF_n215,
         dp_id_stage_regfile_DataPath_Physical_RF_n214,
         dp_id_stage_regfile_DataPath_Physical_RF_n213,
         dp_id_stage_regfile_DataPath_Physical_RF_n212,
         dp_id_stage_regfile_DataPath_Physical_RF_n211,
         dp_id_stage_regfile_DataPath_Physical_RF_n210,
         dp_id_stage_regfile_DataPath_Physical_RF_n209,
         dp_id_stage_regfile_DataPath_Physical_RF_n208,
         dp_id_stage_regfile_DataPath_Physical_RF_n207,
         dp_id_stage_regfile_DataPath_Physical_RF_n206,
         dp_id_stage_regfile_DataPath_Physical_RF_n205,
         dp_id_stage_regfile_DataPath_Physical_RF_n204,
         dp_id_stage_regfile_DataPath_Physical_RF_n203,
         dp_id_stage_regfile_DataPath_Physical_RF_n202,
         dp_id_stage_regfile_DataPath_Physical_RF_n201,
         dp_id_stage_regfile_DataPath_Physical_RF_n200,
         dp_id_stage_regfile_DataPath_Physical_RF_n199,
         dp_id_stage_regfile_DataPath_Physical_RF_n198,
         dp_id_stage_regfile_DataPath_Physical_RF_n197,
         dp_id_stage_regfile_DataPath_Physical_RF_n196,
         dp_id_stage_regfile_DataPath_Physical_RF_n195,
         dp_id_stage_regfile_DataPath_Physical_RF_n194,
         dp_id_stage_regfile_DataPath_Physical_RF_n193,
         dp_id_stage_regfile_DataPath_Physical_RF_n192,
         dp_id_stage_regfile_DataPath_Physical_RF_n191,
         dp_id_stage_regfile_DataPath_Physical_RF_n190,
         dp_id_stage_regfile_DataPath_Physical_RF_n189,
         dp_id_stage_regfile_DataPath_Physical_RF_n188,
         dp_id_stage_regfile_DataPath_Physical_RF_n187,
         dp_id_stage_regfile_DataPath_Physical_RF_n186,
         dp_id_stage_regfile_DataPath_Physical_RF_n185,
         dp_id_stage_regfile_DataPath_Physical_RF_n184,
         dp_id_stage_regfile_DataPath_Physical_RF_n183,
         dp_id_stage_regfile_DataPath_Physical_RF_n182,
         dp_id_stage_regfile_DataPath_Physical_RF_n181,
         dp_id_stage_regfile_DataPath_Physical_RF_n180,
         dp_id_stage_regfile_DataPath_Physical_RF_n179,
         dp_id_stage_regfile_DataPath_Physical_RF_n178,
         dp_id_stage_regfile_DataPath_Physical_RF_n177,
         dp_id_stage_regfile_DataPath_Physical_RF_n176,
         dp_id_stage_regfile_DataPath_Physical_RF_n175,
         dp_id_stage_regfile_DataPath_Physical_RF_n174,
         dp_id_stage_regfile_DataPath_Physical_RF_n173,
         dp_id_stage_regfile_DataPath_Physical_RF_n172,
         dp_id_stage_regfile_DataPath_Physical_RF_n171,
         dp_id_stage_regfile_DataPath_Physical_RF_n170,
         dp_id_stage_regfile_DataPath_Physical_RF_n169,
         dp_id_stage_regfile_DataPath_Physical_RF_n168,
         dp_id_stage_regfile_DataPath_Physical_RF_n167,
         dp_id_stage_regfile_DataPath_Physical_RF_n166,
         dp_id_stage_regfile_DataPath_Physical_RF_n165,
         dp_id_stage_regfile_DataPath_Physical_RF_n164,
         dp_id_stage_regfile_DataPath_Physical_RF_n163,
         dp_id_stage_regfile_DataPath_Physical_RF_n162,
         dp_id_stage_regfile_DataPath_Physical_RF_n161,
         dp_id_stage_regfile_DataPath_Physical_RF_n160,
         dp_id_stage_regfile_DataPath_Physical_RF_n159,
         dp_id_stage_regfile_DataPath_Physical_RF_n158,
         dp_id_stage_regfile_DataPath_Physical_RF_n157,
         dp_id_stage_regfile_DataPath_Physical_RF_n156,
         dp_id_stage_regfile_DataPath_Physical_RF_n155,
         dp_id_stage_regfile_DataPath_Physical_RF_n154,
         dp_id_stage_regfile_DataPath_Physical_RF_n153,
         dp_id_stage_regfile_DataPath_Physical_RF_n152,
         dp_id_stage_regfile_DataPath_Physical_RF_n151,
         dp_id_stage_regfile_DataPath_Physical_RF_n150,
         dp_id_stage_regfile_DataPath_Physical_RF_n149,
         dp_id_stage_regfile_DataPath_Physical_RF_n148,
         dp_id_stage_regfile_DataPath_Physical_RF_n147,
         dp_id_stage_regfile_DataPath_Physical_RF_n146,
         dp_id_stage_regfile_DataPath_Physical_RF_n145,
         dp_id_stage_regfile_DataPath_Physical_RF_n144,
         dp_id_stage_regfile_DataPath_Physical_RF_n143,
         dp_id_stage_regfile_DataPath_Physical_RF_n142,
         dp_id_stage_regfile_DataPath_Physical_RF_n141,
         dp_id_stage_regfile_DataPath_Physical_RF_n140,
         dp_id_stage_regfile_DataPath_Physical_RF_n139,
         dp_id_stage_regfile_DataPath_Physical_RF_n138,
         dp_id_stage_regfile_DataPath_Physical_RF_n137,
         dp_id_stage_regfile_DataPath_Physical_RF_n136,
         dp_id_stage_regfile_DataPath_Physical_RF_n135,
         dp_id_stage_regfile_DataPath_Physical_RF_n134,
         dp_id_stage_regfile_DataPath_Physical_RF_n133,
         dp_id_stage_regfile_DataPath_Physical_RF_n132,
         dp_id_stage_regfile_DataPath_Physical_RF_n131,
         dp_id_stage_regfile_DataPath_Physical_RF_n130,
         dp_id_stage_regfile_DataPath_Physical_RF_n129,
         dp_id_stage_regfile_DataPath_Physical_RF_n128,
         dp_id_stage_regfile_DataPath_Physical_RF_n127,
         dp_id_stage_regfile_DataPath_Physical_RF_n126,
         dp_id_stage_regfile_DataPath_Physical_RF_n125,
         dp_id_stage_regfile_DataPath_Physical_RF_n124,
         dp_id_stage_regfile_DataPath_Physical_RF_n123,
         dp_id_stage_regfile_DataPath_Physical_RF_n122,
         dp_id_stage_regfile_DataPath_Physical_RF_n121,
         dp_id_stage_regfile_DataPath_Physical_RF_n120,
         dp_id_stage_regfile_DataPath_Physical_RF_n119,
         dp_id_stage_regfile_DataPath_Physical_RF_n118,
         dp_id_stage_regfile_DataPath_Physical_RF_n117,
         dp_id_stage_regfile_DataPath_Physical_RF_n116,
         dp_id_stage_regfile_DataPath_Physical_RF_n115,
         dp_id_stage_regfile_DataPath_Physical_RF_n114,
         dp_id_stage_regfile_DataPath_Physical_RF_n113,
         dp_id_stage_regfile_DataPath_Physical_RF_n112,
         dp_id_stage_regfile_DataPath_Physical_RF_n111,
         dp_id_stage_regfile_DataPath_Physical_RF_n110,
         dp_id_stage_regfile_DataPath_Physical_RF_n109,
         dp_id_stage_regfile_DataPath_Physical_RF_n108,
         dp_id_stage_regfile_DataPath_Physical_RF_n107,
         dp_id_stage_regfile_DataPath_Physical_RF_n106,
         dp_id_stage_regfile_DataPath_Physical_RF_n105,
         dp_id_stage_regfile_DataPath_Physical_RF_n104,
         dp_id_stage_regfile_DataPath_Physical_RF_n103,
         dp_id_stage_regfile_DataPath_Physical_RF_n102,
         dp_id_stage_regfile_DataPath_Physical_RF_n101,
         dp_id_stage_regfile_DataPath_Physical_RF_n100,
         dp_id_stage_regfile_DataPath_Physical_RF_n99,
         dp_id_stage_regfile_DataPath_Physical_RF_n98,
         dp_id_stage_regfile_DataPath_Physical_RF_n97,
         dp_id_stage_regfile_DataPath_Physical_RF_n96,
         dp_id_stage_regfile_DataPath_Physical_RF_n95,
         dp_id_stage_regfile_DataPath_Physical_RF_n94,
         dp_id_stage_regfile_DataPath_Physical_RF_n93,
         dp_id_stage_regfile_DataPath_Physical_RF_n92,
         dp_id_stage_regfile_DataPath_Physical_RF_n91,
         dp_id_stage_regfile_DataPath_Physical_RF_n90,
         dp_id_stage_regfile_DataPath_Physical_RF_n89,
         dp_id_stage_regfile_DataPath_Physical_RF_n88,
         dp_id_stage_regfile_DataPath_Physical_RF_n87,
         dp_id_stage_regfile_DataPath_Physical_RF_n86,
         dp_id_stage_regfile_DataPath_Physical_RF_n85,
         dp_id_stage_regfile_DataPath_Physical_RF_n84,
         dp_id_stage_regfile_DataPath_Physical_RF_n83,
         dp_id_stage_regfile_DataPath_Physical_RF_n82,
         dp_id_stage_regfile_DataPath_Physical_RF_n81,
         dp_id_stage_regfile_DataPath_Physical_RF_n80,
         dp_id_stage_regfile_DataPath_Physical_RF_n79,
         dp_id_stage_regfile_DataPath_Physical_RF_n78,
         dp_id_stage_regfile_DataPath_Physical_RF_n77,
         dp_id_stage_regfile_DataPath_Physical_RF_n76,
         dp_id_stage_regfile_DataPath_Physical_RF_n75,
         dp_id_stage_regfile_DataPath_Physical_RF_n74,
         dp_id_stage_regfile_DataPath_Physical_RF_n73,
         dp_id_stage_regfile_DataPath_Physical_RF_n72,
         dp_id_stage_regfile_DataPath_Physical_RF_n71,
         dp_id_stage_regfile_DataPath_Physical_RF_n70,
         dp_id_stage_regfile_DataPath_Physical_RF_n69,
         dp_id_stage_regfile_DataPath_Physical_RF_n68,
         dp_id_stage_regfile_DataPath_Physical_RF_n67,
         dp_id_stage_regfile_DataPath_Physical_RF_n66,
         dp_id_stage_regfile_DataPath_Physical_RF_n65,
         dp_id_stage_regfile_DataPath_Physical_RF_n64,
         dp_id_stage_regfile_DataPath_Physical_RF_n63,
         dp_id_stage_regfile_DataPath_Physical_RF_n62,
         dp_id_stage_regfile_DataPath_Physical_RF_n61,
         dp_id_stage_regfile_DataPath_Physical_RF_n60,
         dp_id_stage_regfile_DataPath_Physical_RF_n59,
         dp_id_stage_regfile_DataPath_Physical_RF_n58,
         dp_id_stage_regfile_DataPath_Physical_RF_n57,
         dp_id_stage_regfile_DataPath_Physical_RF_n56,
         dp_id_stage_regfile_DataPath_Physical_RF_n55,
         dp_id_stage_regfile_DataPath_Physical_RF_n54,
         dp_id_stage_regfile_DataPath_Physical_RF_n53,
         dp_id_stage_regfile_DataPath_Physical_RF_n52,
         dp_id_stage_regfile_DataPath_Physical_RF_n51,
         dp_id_stage_regfile_DataPath_Physical_RF_n50,
         dp_id_stage_regfile_DataPath_Physical_RF_n49,
         dp_id_stage_regfile_DataPath_Physical_RF_n48,
         dp_id_stage_regfile_DataPath_Physical_RF_n47,
         dp_id_stage_regfile_DataPath_Physical_RF_n46,
         dp_id_stage_regfile_DataPath_Physical_RF_n45,
         dp_id_stage_regfile_DataPath_Physical_RF_n44,
         dp_id_stage_regfile_DataPath_Physical_RF_n43,
         dp_id_stage_regfile_DataPath_Physical_RF_n42,
         dp_id_stage_regfile_DataPath_Physical_RF_n41,
         dp_id_stage_regfile_DataPath_Physical_RF_n40,
         dp_id_stage_regfile_DataPath_Physical_RF_n39,
         dp_id_stage_regfile_DataPath_Physical_RF_n38,
         dp_id_stage_regfile_DataPath_Physical_RF_n37,
         dp_id_stage_regfile_DataPath_Physical_RF_n36,
         dp_id_stage_regfile_DataPath_Physical_RF_n35,
         dp_id_stage_regfile_DataPath_Physical_RF_n34,
         dp_id_stage_regfile_DataPath_Physical_RF_n33,
         dp_id_stage_regfile_DataPath_Physical_RF_n32,
         dp_id_stage_regfile_DataPath_Physical_RF_n31,
         dp_id_stage_regfile_DataPath_Physical_RF_n30,
         dp_id_stage_regfile_DataPath_Physical_RF_n29,
         dp_id_stage_regfile_DataPath_Physical_RF_n28,
         dp_id_stage_regfile_DataPath_Physical_RF_n27,
         dp_id_stage_regfile_DataPath_Physical_RF_n26,
         dp_id_stage_regfile_DataPath_Physical_RF_n25,
         dp_id_stage_regfile_DataPath_Physical_RF_n24,
         dp_id_stage_regfile_DataPath_Physical_RF_n23,
         dp_id_stage_regfile_DataPath_Physical_RF_n22,
         dp_id_stage_regfile_DataPath_Physical_RF_n21,
         dp_id_stage_regfile_DataPath_Physical_RF_n20,
         dp_id_stage_regfile_DataPath_Physical_RF_n19,
         dp_id_stage_regfile_DataPath_Physical_RF_n18,
         dp_id_stage_regfile_DataPath_Physical_RF_n17,
         dp_id_stage_regfile_DataPath_Physical_RF_n16,
         dp_id_stage_regfile_DataPath_Physical_RF_n15,
         dp_id_stage_regfile_DataPath_Physical_RF_n14,
         dp_id_stage_regfile_DataPath_Physical_RF_n13,
         dp_id_stage_regfile_DataPath_Physical_RF_n12,
         dp_id_stage_regfile_DataPath_Physical_RF_n11,
         dp_id_stage_regfile_DataPath_Physical_RF_n10,
         dp_id_stage_regfile_DataPath_Physical_RF_n9,
         dp_id_stage_regfile_DataPath_Physical_RF_n8,
         dp_id_stage_regfile_DataPath_Physical_RF_n7,
         dp_id_stage_regfile_DataPath_Physical_RF_n6,
         dp_id_stage_regfile_DataPath_Physical_RF_n5,
         dp_id_stage_regfile_DataPath_Physical_RF_n4,
         dp_id_stage_regfile_DataPath_Physical_RF_n3,
         dp_id_stage_regfile_DataPath_Physical_RF_n2,
         dp_id_stage_regfile_DataPath_Physical_RF_N429,
         dp_id_stage_regfile_DataPath_Physical_RF_N428,
         dp_id_stage_regfile_DataPath_Physical_RF_N427,
         dp_id_stage_regfile_DataPath_Physical_RF_N426,
         dp_id_stage_regfile_DataPath_Physical_RF_N425,
         dp_id_stage_regfile_DataPath_Physical_RF_N424,
         dp_id_stage_regfile_DataPath_Physical_RF_N423,
         dp_id_stage_regfile_DataPath_Physical_RF_N422,
         dp_id_stage_regfile_DataPath_Physical_RF_N421,
         dp_id_stage_regfile_DataPath_Physical_RF_N420,
         dp_id_stage_regfile_DataPath_Physical_RF_N419,
         dp_id_stage_regfile_DataPath_Physical_RF_N418,
         dp_id_stage_regfile_DataPath_Physical_RF_N417,
         dp_id_stage_regfile_DataPath_Physical_RF_N416,
         dp_id_stage_regfile_DataPath_Physical_RF_N415,
         dp_id_stage_regfile_DataPath_Physical_RF_N414,
         dp_id_stage_regfile_DataPath_Physical_RF_N413,
         dp_id_stage_regfile_DataPath_Physical_RF_N412,
         dp_id_stage_regfile_DataPath_Physical_RF_N411,
         dp_id_stage_regfile_DataPath_Physical_RF_N410,
         dp_id_stage_regfile_DataPath_Physical_RF_N409,
         dp_id_stage_regfile_DataPath_Physical_RF_N408,
         dp_id_stage_regfile_DataPath_Physical_RF_N407,
         dp_id_stage_regfile_DataPath_Physical_RF_N406,
         dp_id_stage_regfile_DataPath_Physical_RF_N405,
         dp_id_stage_regfile_DataPath_Physical_RF_N404,
         dp_id_stage_regfile_DataPath_Physical_RF_N403,
         dp_id_stage_regfile_DataPath_Physical_RF_N402,
         dp_id_stage_regfile_DataPath_Physical_RF_N401,
         dp_id_stage_regfile_DataPath_Physical_RF_N400,
         dp_id_stage_regfile_DataPath_Physical_RF_N399,
         dp_id_stage_regfile_DataPath_Physical_RF_N398,
         dp_id_stage_regfile_DataPath_Physical_RF_N397,
         dp_id_stage_regfile_DataPath_Physical_RF_N396,
         dp_id_stage_regfile_DataPath_Physical_RF_N359,
         dp_id_stage_regfile_DataPath_Physical_RF_N358,
         dp_id_stage_regfile_DataPath_Physical_RF_N357,
         dp_id_stage_regfile_DataPath_Physical_RF_N356,
         dp_id_stage_regfile_DataPath_Physical_RF_N355,
         dp_id_stage_regfile_DataPath_Physical_RF_N354,
         dp_id_stage_regfile_DataPath_Physical_RF_N353,
         dp_id_stage_regfile_DataPath_Physical_RF_N352,
         dp_id_stage_regfile_DataPath_Physical_RF_N351,
         dp_id_stage_regfile_DataPath_Physical_RF_N350,
         dp_id_stage_regfile_DataPath_Physical_RF_N349,
         dp_id_stage_regfile_DataPath_Physical_RF_N348,
         dp_id_stage_regfile_DataPath_Physical_RF_N347,
         dp_id_stage_regfile_DataPath_Physical_RF_N346,
         dp_id_stage_regfile_DataPath_Physical_RF_N345,
         dp_id_stage_regfile_DataPath_Physical_RF_N344,
         dp_id_stage_regfile_DataPath_Physical_RF_N343,
         dp_id_stage_regfile_DataPath_Physical_RF_N342,
         dp_id_stage_regfile_DataPath_Physical_RF_N341,
         dp_id_stage_regfile_DataPath_Physical_RF_N340,
         dp_id_stage_regfile_DataPath_Physical_RF_N339,
         dp_id_stage_regfile_DataPath_Physical_RF_N338,
         dp_id_stage_regfile_DataPath_Physical_RF_N337,
         dp_id_stage_regfile_DataPath_Physical_RF_N336,
         dp_id_stage_regfile_DataPath_Physical_RF_N335,
         dp_id_stage_regfile_DataPath_Physical_RF_N334,
         dp_id_stage_regfile_DataPath_Physical_RF_N333,
         dp_id_stage_regfile_DataPath_Physical_RF_N332,
         dp_id_stage_regfile_DataPath_Physical_RF_N331,
         dp_id_stage_regfile_DataPath_Physical_RF_N330,
         dp_id_stage_regfile_DataPath_Physical_RF_N329,
         dp_id_stage_regfile_DataPath_Physical_RF_N328,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__31_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__0_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__1_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__2_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__3_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__4_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__5_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__6_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__7_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__8_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__9_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__10_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__11_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__12_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__13_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__14_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__15_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__16_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__17_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__18_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__19_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__20_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__21_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__22_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__23_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__24_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__25_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__26_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__27_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__28_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__29_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__30_,
         dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__31_,
         dp_ex_stage_n10, dp_ex_stage_n9, dp_ex_stage_n8, dp_ex_stage_n7,
         dp_ex_stage_n6, dp_ex_stage_n5, dp_ex_stage_n4, dp_ex_stage_n3,
         dp_ex_stage_n2, dp_ex_stage_n1, dp_ex_stage_muxA_n27,
         dp_ex_stage_muxA_n8, dp_ex_stage_muxA_n7, dp_ex_stage_muxA_n6,
         dp_ex_stage_muxA_n5, dp_ex_stage_muxA_n4, dp_ex_stage_muxA_n3,
         dp_ex_stage_muxA_n2, dp_ex_stage_muxB_n8, dp_ex_stage_muxB_n7,
         dp_ex_stage_muxB_n6, dp_ex_stage_muxB_n5, dp_ex_stage_muxB_n4,
         dp_ex_stage_muxB_n3, dp_ex_stage_muxB_n2, dp_ex_stage_muxB_n1,
         dp_ex_stage_alu_n311, dp_ex_stage_alu_n310, dp_ex_stage_alu_n309,
         dp_ex_stage_alu_n308, dp_ex_stage_alu_n307, dp_ex_stage_alu_n306,
         dp_ex_stage_alu_n305, dp_ex_stage_alu_n304, dp_ex_stage_alu_n303,
         dp_ex_stage_alu_n302, dp_ex_stage_alu_n301, dp_ex_stage_alu_n300,
         dp_ex_stage_alu_n299, dp_ex_stage_alu_n298, dp_ex_stage_alu_n297,
         dp_ex_stage_alu_n296, dp_ex_stage_alu_n295, dp_ex_stage_alu_n294,
         dp_ex_stage_alu_n293, dp_ex_stage_alu_n292, dp_ex_stage_alu_n291,
         dp_ex_stage_alu_n290, dp_ex_stage_alu_n289, dp_ex_stage_alu_n288,
         dp_ex_stage_alu_n287, dp_ex_stage_alu_n286, dp_ex_stage_alu_n285,
         dp_ex_stage_alu_n284, dp_ex_stage_alu_n283, dp_ex_stage_alu_n282,
         dp_ex_stage_alu_n281, dp_ex_stage_alu_n280, dp_ex_stage_alu_n279,
         dp_ex_stage_alu_n278, dp_ex_stage_alu_n277, dp_ex_stage_alu_n276,
         dp_ex_stage_alu_n275, dp_ex_stage_alu_n274, dp_ex_stage_alu_n273,
         dp_ex_stage_alu_n272, dp_ex_stage_alu_n271, dp_ex_stage_alu_n270,
         dp_ex_stage_alu_n269, dp_ex_stage_alu_n268, dp_ex_stage_alu_n267,
         dp_ex_stage_alu_n266, dp_ex_stage_alu_n265, dp_ex_stage_alu_n264,
         dp_ex_stage_alu_n263, dp_ex_stage_alu_n262, dp_ex_stage_alu_n261,
         dp_ex_stage_alu_n260, dp_ex_stage_alu_n259, dp_ex_stage_alu_n258,
         dp_ex_stage_alu_n257, dp_ex_stage_alu_n256, dp_ex_stage_alu_n255,
         dp_ex_stage_alu_n254, dp_ex_stage_alu_n253, dp_ex_stage_alu_n252,
         dp_ex_stage_alu_n251, dp_ex_stage_alu_n250, dp_ex_stage_alu_n249,
         dp_ex_stage_alu_n248, dp_ex_stage_alu_n247, dp_ex_stage_alu_n246,
         dp_ex_stage_alu_n245, dp_ex_stage_alu_n244, dp_ex_stage_alu_n243,
         dp_ex_stage_alu_n242, dp_ex_stage_alu_n241, dp_ex_stage_alu_n240,
         dp_ex_stage_alu_n239, dp_ex_stage_alu_n238, dp_ex_stage_alu_n237,
         dp_ex_stage_alu_n236, dp_ex_stage_alu_n235, dp_ex_stage_alu_n234,
         dp_ex_stage_alu_n233, dp_ex_stage_alu_n232, dp_ex_stage_alu_n231,
         dp_ex_stage_alu_n230, dp_ex_stage_alu_n229, dp_ex_stage_alu_n228,
         dp_ex_stage_alu_n227, dp_ex_stage_alu_n226, dp_ex_stage_alu_n225,
         dp_ex_stage_alu_n224, dp_ex_stage_alu_n223, dp_ex_stage_alu_n222,
         dp_ex_stage_alu_n221, dp_ex_stage_alu_n220, dp_ex_stage_alu_n219,
         dp_ex_stage_alu_n218, dp_ex_stage_alu_n217, dp_ex_stage_alu_n216,
         dp_ex_stage_alu_n215, dp_ex_stage_alu_n214, dp_ex_stage_alu_n213,
         dp_ex_stage_alu_n212, dp_ex_stage_alu_n211, dp_ex_stage_alu_n210,
         dp_ex_stage_alu_n209, dp_ex_stage_alu_n207, dp_ex_stage_alu_n204,
         dp_ex_stage_alu_n203, dp_ex_stage_alu_n202, dp_ex_stage_alu_n201,
         dp_ex_stage_alu_n200, dp_ex_stage_alu_n199, dp_ex_stage_alu_n198,
         dp_ex_stage_alu_n197, dp_ex_stage_alu_n196, dp_ex_stage_alu_n195,
         dp_ex_stage_alu_n194, dp_ex_stage_alu_n193, dp_ex_stage_alu_n192,
         dp_ex_stage_alu_n191, dp_ex_stage_alu_n93, dp_ex_stage_alu_n92,
         dp_ex_stage_alu_n89, dp_ex_stage_alu_n88, dp_ex_stage_alu_n87,
         dp_ex_stage_alu_n86, dp_ex_stage_alu_n85, dp_ex_stage_alu_n84,
         dp_ex_stage_alu_n83, dp_ex_stage_alu_n82, dp_ex_stage_alu_n81,
         dp_ex_stage_alu_n80, dp_ex_stage_alu_n79, dp_ex_stage_alu_n78,
         dp_ex_stage_alu_n77, dp_ex_stage_alu_n76, dp_ex_stage_alu_n74,
         dp_ex_stage_alu_n73, dp_ex_stage_alu_n72, dp_ex_stage_alu_n71,
         dp_ex_stage_alu_n70, dp_ex_stage_alu_n69, dp_ex_stage_alu_n68,
         dp_ex_stage_alu_n67, dp_ex_stage_alu_n66, dp_ex_stage_alu_n65,
         dp_ex_stage_alu_n64, dp_ex_stage_alu_n63, dp_ex_stage_alu_n62,
         dp_ex_stage_alu_n61, dp_ex_stage_alu_n60, dp_ex_stage_alu_n59,
         dp_ex_stage_alu_n58, dp_ex_stage_alu_n57, dp_ex_stage_alu_n56,
         dp_ex_stage_alu_n55, dp_ex_stage_alu_n54, dp_ex_stage_alu_n53,
         dp_ex_stage_alu_n52, dp_ex_stage_alu_n51, dp_ex_stage_alu_n50,
         dp_ex_stage_alu_n49, dp_ex_stage_alu_n48, dp_ex_stage_alu_n47,
         dp_ex_stage_alu_n46, dp_ex_stage_alu_n45, dp_ex_stage_alu_n44,
         dp_ex_stage_alu_n43, dp_ex_stage_alu_n42, dp_ex_stage_alu_n41,
         dp_ex_stage_alu_n40, dp_ex_stage_alu_n39, dp_ex_stage_alu_n38,
         dp_ex_stage_alu_n37, dp_ex_stage_alu_n36, dp_ex_stage_alu_n35,
         dp_ex_stage_alu_n34, dp_ex_stage_alu_n33, dp_ex_stage_alu_n32,
         dp_ex_stage_alu_n31, dp_ex_stage_alu_n30, dp_ex_stage_alu_n29,
         dp_ex_stage_alu_n28, dp_ex_stage_alu_n27, dp_ex_stage_alu_n26,
         dp_ex_stage_alu_n25, dp_ex_stage_alu_n24, dp_ex_stage_alu_n23,
         dp_ex_stage_alu_n22, dp_ex_stage_alu_n21, dp_ex_stage_alu_n20,
         dp_ex_stage_alu_n19, dp_ex_stage_alu_n18, dp_ex_stage_alu_n17,
         dp_ex_stage_alu_n16, dp_ex_stage_alu_n15, dp_ex_stage_alu_n14,
         dp_ex_stage_alu_n11, dp_ex_stage_alu_n10, dp_ex_stage_alu_n9,
         dp_ex_stage_alu_n8, dp_ex_stage_alu_n7, dp_ex_stage_alu_n6,
         dp_ex_stage_alu_n5, dp_ex_stage_alu_n4, dp_ex_stage_alu_n3,
         dp_ex_stage_alu_n2, dp_ex_stage_alu_n1, dp_ex_stage_alu_n208,
         dp_ex_stage_alu_n206, dp_ex_stage_alu_n205, dp_ex_stage_alu_n190,
         dp_ex_stage_alu_n189, dp_ex_stage_alu_n188, dp_ex_stage_alu_n187,
         dp_ex_stage_alu_n186, dp_ex_stage_alu_n185, dp_ex_stage_alu_n184,
         dp_ex_stage_alu_n183, dp_ex_stage_alu_n182, dp_ex_stage_alu_n181,
         dp_ex_stage_alu_n180, dp_ex_stage_alu_n179, dp_ex_stage_alu_n178,
         dp_ex_stage_alu_n177, dp_ex_stage_alu_n176, dp_ex_stage_alu_n175,
         dp_ex_stage_alu_n174, dp_ex_stage_alu_n173, dp_ex_stage_alu_n172,
         dp_ex_stage_alu_n171, dp_ex_stage_alu_n170, dp_ex_stage_alu_n169,
         dp_ex_stage_alu_n168, dp_ex_stage_alu_n167, dp_ex_stage_alu_n166,
         dp_ex_stage_alu_n165, dp_ex_stage_alu_n164, dp_ex_stage_alu_n163,
         dp_ex_stage_alu_n162, dp_ex_stage_alu_n161, dp_ex_stage_alu_n160,
         dp_ex_stage_alu_n159, dp_ex_stage_alu_n158, dp_ex_stage_alu_n157,
         dp_ex_stage_alu_n156, dp_ex_stage_alu_n155, dp_ex_stage_alu_n154,
         dp_ex_stage_alu_n153, dp_ex_stage_alu_n152, dp_ex_stage_alu_n151,
         dp_ex_stage_alu_n150, dp_ex_stage_alu_n149, dp_ex_stage_alu_n148,
         dp_ex_stage_alu_n147, dp_ex_stage_alu_n146, dp_ex_stage_alu_n145,
         dp_ex_stage_alu_n144, dp_ex_stage_alu_n143, dp_ex_stage_alu_n142,
         dp_ex_stage_alu_n141, dp_ex_stage_alu_n140, dp_ex_stage_alu_n139,
         dp_ex_stage_alu_n138, dp_ex_stage_alu_n137, dp_ex_stage_alu_n136,
         dp_ex_stage_alu_n135, dp_ex_stage_alu_n134, dp_ex_stage_alu_n133,
         dp_ex_stage_alu_n132, dp_ex_stage_alu_n131, dp_ex_stage_alu_n130,
         dp_ex_stage_alu_n129, dp_ex_stage_alu_n128, dp_ex_stage_alu_n127,
         dp_ex_stage_alu_n126, dp_ex_stage_alu_n125, dp_ex_stage_alu_n124,
         dp_ex_stage_alu_n123, dp_ex_stage_alu_n122, dp_ex_stage_alu_n121,
         dp_ex_stage_alu_n120, dp_ex_stage_alu_n119, dp_ex_stage_alu_n118,
         dp_ex_stage_alu_n117, dp_ex_stage_alu_n116, dp_ex_stage_alu_n115,
         dp_ex_stage_alu_n114, dp_ex_stage_alu_n113, dp_ex_stage_alu_n112,
         dp_ex_stage_alu_n111, dp_ex_stage_alu_n110, dp_ex_stage_alu_n109,
         dp_ex_stage_alu_n108, dp_ex_stage_alu_n107, dp_ex_stage_alu_n106,
         dp_ex_stage_alu_n105, dp_ex_stage_alu_n104, dp_ex_stage_alu_n103,
         dp_ex_stage_alu_n102, dp_ex_stage_alu_n101, dp_ex_stage_alu_n100,
         dp_ex_stage_alu_n99, dp_ex_stage_alu_n98, dp_ex_stage_alu_n97,
         dp_ex_stage_alu_n96, dp_ex_stage_alu_n95, dp_ex_stage_alu_n94,
         dp_ex_stage_alu_n91, dp_ex_stage_alu_n90, dp_ex_stage_alu_N23,
         dp_ex_stage_alu_shift_arith_i, dp_ex_stage_alu_N22,
         dp_ex_stage_alu_N21, dp_ex_stage_alu_N20, dp_ex_stage_alu_N19,
         dp_ex_stage_alu_N18, dp_ex_stage_alu_N17, dp_ex_stage_alu_N16,
         dp_ex_stage_alu_adder_n23, dp_ex_stage_alu_adder_n22,
         dp_ex_stage_alu_adder_n21, dp_ex_stage_alu_adder_n20,
         dp_ex_stage_alu_adder_n19, dp_ex_stage_alu_adder_n18,
         dp_ex_stage_alu_adder_n17, dp_ex_stage_alu_adder_n16,
         dp_ex_stage_alu_adder_n15, dp_ex_stage_alu_adder_n14,
         dp_ex_stage_alu_adder_n13, dp_ex_stage_alu_adder_n12,
         dp_ex_stage_alu_adder_n11, dp_ex_stage_alu_adder_n10,
         dp_ex_stage_alu_adder_n9, dp_ex_stage_alu_adder_n8,
         dp_ex_stage_alu_adder_n7, dp_ex_stage_alu_adder_n6,
         dp_ex_stage_alu_adder_n5, dp_ex_stage_alu_adder_n4,
         dp_ex_stage_alu_adder_n3, dp_ex_stage_alu_adder_n2,
         dp_ex_stage_alu_adder_n1, dp_ex_stage_alu_adder_B_xor_0_,
         dp_ex_stage_alu_adder_B_xor_1_, dp_ex_stage_alu_adder_B_xor_2_,
         dp_ex_stage_alu_adder_B_xor_3_, dp_ex_stage_alu_adder_B_xor_4_,
         dp_ex_stage_alu_adder_B_xor_6_, dp_ex_stage_alu_adder_B_xor_8_,
         dp_ex_stage_alu_adder_B_xor_9_, dp_ex_stage_alu_adder_B_xor_10_,
         dp_ex_stage_alu_adder_B_xor_11_, dp_ex_stage_alu_adder_B_xor_12_,
         dp_ex_stage_alu_adder_B_xor_13_, dp_ex_stage_alu_adder_B_xor_14_,
         dp_ex_stage_alu_adder_B_xor_16_, dp_ex_stage_alu_adder_B_xor_17_,
         dp_ex_stage_alu_adder_B_xor_18_, dp_ex_stage_alu_adder_B_xor_19_,
         dp_ex_stage_alu_adder_B_xor_20_, dp_ex_stage_alu_adder_B_xor_21_,
         dp_ex_stage_alu_adder_B_xor_22_, dp_ex_stage_alu_adder_B_xor_23_,
         dp_ex_stage_alu_adder_B_xor_24_, dp_ex_stage_alu_adder_B_xor_25_,
         dp_ex_stage_alu_adder_B_xor_26_, dp_ex_stage_alu_adder_B_xor_27_,
         dp_ex_stage_alu_adder_B_xor_28_, dp_ex_stage_alu_adder_B_xor_29_,
         dp_ex_stage_alu_adder_B_xor_30_, dp_ex_stage_alu_adder_B_xor_31_,
         dp_ex_stage_alu_adder_Cout, dp_ex_stage_alu_adder_SparseTree_n4,
         dp_ex_stage_alu_adder_SparseTree_n3,
         dp_ex_stage_alu_adder_SparseTree_n1,
         dp_ex_stage_alu_adder_SparseTree_prop_2__2_,
         dp_ex_stage_alu_adder_SparseTree_prop_3__3_,
         dp_ex_stage_alu_adder_SparseTree_prop_4__3_,
         dp_ex_stage_alu_adder_SparseTree_prop_4__4_,
         dp_ex_stage_alu_adder_SparseTree_prop_5__5_,
         dp_ex_stage_alu_adder_SparseTree_prop_6__5_,
         dp_ex_stage_alu_adder_SparseTree_prop_6__6_,
         dp_ex_stage_alu_adder_SparseTree_prop_7__7_,
         dp_ex_stage_alu_adder_SparseTree_prop_8__5_,
         dp_ex_stage_alu_adder_SparseTree_prop_8__7_,
         dp_ex_stage_alu_adder_SparseTree_prop_8__8_,
         dp_ex_stage_alu_adder_SparseTree_prop_9__9_,
         dp_ex_stage_alu_adder_SparseTree_prop_10__9_,
         dp_ex_stage_alu_adder_SparseTree_prop_10__10_,
         dp_ex_stage_alu_adder_SparseTree_prop_11__11_,
         dp_ex_stage_alu_adder_SparseTree_prop_12__9_,
         dp_ex_stage_alu_adder_SparseTree_prop_12__11_,
         dp_ex_stage_alu_adder_SparseTree_prop_12__12_,
         dp_ex_stage_alu_adder_SparseTree_prop_13__13_,
         dp_ex_stage_alu_adder_SparseTree_prop_14__13_,
         dp_ex_stage_alu_adder_SparseTree_prop_14__14_,
         dp_ex_stage_alu_adder_SparseTree_prop_15__15_,
         dp_ex_stage_alu_adder_SparseTree_prop_16__9_,
         dp_ex_stage_alu_adder_SparseTree_prop_16__13_,
         dp_ex_stage_alu_adder_SparseTree_prop_16__15_,
         dp_ex_stage_alu_adder_SparseTree_prop_16__16_,
         dp_ex_stage_alu_adder_SparseTree_prop_17__17_,
         dp_ex_stage_alu_adder_SparseTree_prop_18__17_,
         dp_ex_stage_alu_adder_SparseTree_prop_18__18_,
         dp_ex_stage_alu_adder_SparseTree_prop_19__19_,
         dp_ex_stage_alu_adder_SparseTree_prop_20__17_,
         dp_ex_stage_alu_adder_SparseTree_prop_20__19_,
         dp_ex_stage_alu_adder_SparseTree_prop_20__20_,
         dp_ex_stage_alu_adder_SparseTree_prop_21__21_,
         dp_ex_stage_alu_adder_SparseTree_prop_22__21_,
         dp_ex_stage_alu_adder_SparseTree_prop_22__22_,
         dp_ex_stage_alu_adder_SparseTree_prop_23__23_,
         dp_ex_stage_alu_adder_SparseTree_prop_24__17_,
         dp_ex_stage_alu_adder_SparseTree_prop_24__21_,
         dp_ex_stage_alu_adder_SparseTree_prop_24__23_,
         dp_ex_stage_alu_adder_SparseTree_prop_24__24_,
         dp_ex_stage_alu_adder_SparseTree_prop_25__25_,
         dp_ex_stage_alu_adder_SparseTree_prop_26__25_,
         dp_ex_stage_alu_adder_SparseTree_prop_26__26_,
         dp_ex_stage_alu_adder_SparseTree_prop_27__27_,
         dp_ex_stage_alu_adder_SparseTree_prop_28__17_,
         dp_ex_stage_alu_adder_SparseTree_prop_28__25_,
         dp_ex_stage_alu_adder_SparseTree_prop_28__27_,
         dp_ex_stage_alu_adder_SparseTree_prop_28__28_,
         dp_ex_stage_alu_adder_SparseTree_prop_29__29_,
         dp_ex_stage_alu_adder_SparseTree_prop_30__29_,
         dp_ex_stage_alu_adder_SparseTree_prop_30__30_,
         dp_ex_stage_alu_adder_SparseTree_prop_31__31_,
         dp_ex_stage_alu_adder_SparseTree_prop_32__17_,
         dp_ex_stage_alu_adder_SparseTree_prop_32__25_,
         dp_ex_stage_alu_adder_SparseTree_prop_32__29_,
         dp_ex_stage_alu_adder_SparseTree_prop_32__31_,
         dp_ex_stage_alu_adder_SparseTree_prop_32__32_,
         dp_ex_stage_alu_adder_SparseTree_prop_1__1_,
         dp_ex_stage_alu_adder_SparseTree_gen_2__0_,
         dp_ex_stage_alu_adder_SparseTree_gen_2__2_,
         dp_ex_stage_alu_adder_SparseTree_gen_3__3_,
         dp_ex_stage_alu_adder_SparseTree_gen_4__3_,
         dp_ex_stage_alu_adder_SparseTree_gen_4__4_,
         dp_ex_stage_alu_adder_SparseTree_gen_5__5_,
         dp_ex_stage_alu_adder_SparseTree_gen_6__5_,
         dp_ex_stage_alu_adder_SparseTree_gen_6__6_,
         dp_ex_stage_alu_adder_SparseTree_gen_7__7_,
         dp_ex_stage_alu_adder_SparseTree_gen_8__5_,
         dp_ex_stage_alu_adder_SparseTree_gen_8__7_,
         dp_ex_stage_alu_adder_SparseTree_gen_8__8_,
         dp_ex_stage_alu_adder_SparseTree_gen_9__9_,
         dp_ex_stage_alu_adder_SparseTree_gen_10__9_,
         dp_ex_stage_alu_adder_SparseTree_gen_10__10_,
         dp_ex_stage_alu_adder_SparseTree_gen_11__11_,
         dp_ex_stage_alu_adder_SparseTree_gen_12__9_,
         dp_ex_stage_alu_adder_SparseTree_gen_12__11_,
         dp_ex_stage_alu_adder_SparseTree_gen_12__12_,
         dp_ex_stage_alu_adder_SparseTree_gen_13__13_,
         dp_ex_stage_alu_adder_SparseTree_gen_14__13_,
         dp_ex_stage_alu_adder_SparseTree_gen_14__14_,
         dp_ex_stage_alu_adder_SparseTree_gen_15__15_,
         dp_ex_stage_alu_adder_SparseTree_gen_16__9_,
         dp_ex_stage_alu_adder_SparseTree_gen_16__13_,
         dp_ex_stage_alu_adder_SparseTree_gen_16__15_,
         dp_ex_stage_alu_adder_SparseTree_gen_16__16_,
         dp_ex_stage_alu_adder_SparseTree_gen_17__17_,
         dp_ex_stage_alu_adder_SparseTree_gen_18__17_,
         dp_ex_stage_alu_adder_SparseTree_gen_18__18_,
         dp_ex_stage_alu_adder_SparseTree_gen_19__19_,
         dp_ex_stage_alu_adder_SparseTree_gen_20__17_,
         dp_ex_stage_alu_adder_SparseTree_gen_20__19_,
         dp_ex_stage_alu_adder_SparseTree_gen_20__20_,
         dp_ex_stage_alu_adder_SparseTree_gen_21__21_,
         dp_ex_stage_alu_adder_SparseTree_gen_22__21_,
         dp_ex_stage_alu_adder_SparseTree_gen_22__22_,
         dp_ex_stage_alu_adder_SparseTree_gen_23__23_,
         dp_ex_stage_alu_adder_SparseTree_gen_24__17_,
         dp_ex_stage_alu_adder_SparseTree_gen_24__21_,
         dp_ex_stage_alu_adder_SparseTree_gen_24__23_,
         dp_ex_stage_alu_adder_SparseTree_gen_24__24_,
         dp_ex_stage_alu_adder_SparseTree_gen_25__25_,
         dp_ex_stage_alu_adder_SparseTree_gen_26__25_,
         dp_ex_stage_alu_adder_SparseTree_gen_26__26_,
         dp_ex_stage_alu_adder_SparseTree_gen_27__27_,
         dp_ex_stage_alu_adder_SparseTree_gen_28__17_,
         dp_ex_stage_alu_adder_SparseTree_gen_28__25_,
         dp_ex_stage_alu_adder_SparseTree_gen_28__27_,
         dp_ex_stage_alu_adder_SparseTree_gen_28__28_,
         dp_ex_stage_alu_adder_SparseTree_gen_29__29_,
         dp_ex_stage_alu_adder_SparseTree_gen_30__29_,
         dp_ex_stage_alu_adder_SparseTree_gen_30__30_,
         dp_ex_stage_alu_adder_SparseTree_gen_31__31_,
         dp_ex_stage_alu_adder_SparseTree_gen_32__17_,
         dp_ex_stage_alu_adder_SparseTree_gen_32__25_,
         dp_ex_stage_alu_adder_SparseTree_gen_32__29_,
         dp_ex_stage_alu_adder_SparseTree_gen_32__31_,
         dp_ex_stage_alu_adder_SparseTree_gen_32__32_,
         dp_ex_stage_alu_adder_SparseTree_gen_1__0_,
         dp_ex_stage_alu_adder_SparseTree_gen_1__1_,
         dp_ex_stage_alu_adder_SparseTree_n9,
         dp_ex_stage_alu_adder_SparseTree_n8,
         dp_ex_stage_alu_adder_SparseTree_n7,
         dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_n1,
         dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_n1,
         dp_ex_stage_alu_adder_SparseTree_G10_n2,
         dp_ex_stage_alu_adder_SparseTree_G20_1_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_n2,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_n3,
         dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_n3,
         dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_n3,
         dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_n3,
         dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_n3,
         dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_n3,
         dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_n3,
         dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_n3,
         dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_n3,
         dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_n3,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n9,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n8,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n7,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n6,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n13,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n12,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n11,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n10,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n13,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n12,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n11,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n10,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n13,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n12,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n11,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n10,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n13,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n12,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n11,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n10,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n14,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n13,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n12,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n11,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n10,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n1,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n4,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n3,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n2,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n1,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_3_,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_1_,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n14,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n13,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n12,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n11,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n10,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n1,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_Co,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n14,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n13,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n12,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n11,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n10,
         dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n1,
         dp_ex_stage_alu_shifter_n118, dp_ex_stage_alu_shifter_n117,
         dp_ex_stage_alu_shifter_n116, dp_ex_stage_alu_shifter_n115,
         dp_ex_stage_alu_shifter_n114, dp_ex_stage_alu_shifter_n113,
         dp_ex_stage_alu_shifter_n112, dp_ex_stage_alu_shifter_n111,
         dp_ex_stage_alu_shifter_n110, dp_ex_stage_alu_shifter_n109,
         dp_ex_stage_alu_shifter_n108, dp_ex_stage_alu_shifter_n107,
         dp_ex_stage_alu_shifter_n106, dp_ex_stage_alu_shifter_n105,
         dp_ex_stage_alu_shifter_n104, dp_ex_stage_alu_shifter_n103,
         dp_ex_stage_alu_shifter_n102, dp_ex_stage_alu_shifter_n101,
         dp_ex_stage_alu_shifter_n100, dp_ex_stage_alu_shifter_n99,
         dp_ex_stage_alu_shifter_n98, dp_ex_stage_alu_shifter_n97,
         dp_ex_stage_alu_shifter_n96, dp_ex_stage_alu_shifter_n95,
         dp_ex_stage_alu_shifter_n94, dp_ex_stage_alu_shifter_n93,
         dp_ex_stage_alu_shifter_n20, dp_ex_stage_alu_shifter_n19,
         dp_ex_stage_alu_shifter_n12, dp_ex_stage_alu_shifter_n11,
         dp_ex_stage_alu_shifter_n10, dp_ex_stage_alu_shifter_n9,
         dp_ex_stage_alu_shifter_n8, dp_ex_stage_alu_shifter_n7,
         dp_ex_stage_alu_shifter_n6, dp_ex_stage_alu_shifter_n5,
         dp_ex_stage_alu_shifter_n4, dp_ex_stage_alu_shifter_n3,
         dp_ex_stage_alu_shifter_n2, dp_ex_stage_alu_shifter_n1,
         dp_ex_stage_alu_shifter_n92, dp_ex_stage_alu_shifter_n91,
         dp_ex_stage_alu_shifter_n90, dp_ex_stage_alu_shifter_n89,
         dp_ex_stage_alu_shifter_n88, dp_ex_stage_alu_shifter_n87,
         dp_ex_stage_alu_shifter_n86, dp_ex_stage_alu_shifter_n85,
         dp_ex_stage_alu_shifter_n84, dp_ex_stage_alu_shifter_n83,
         dp_ex_stage_alu_shifter_n82, dp_ex_stage_alu_shifter_n81,
         dp_ex_stage_alu_shifter_n80, dp_ex_stage_alu_shifter_n79,
         dp_ex_stage_alu_shifter_n78, dp_ex_stage_alu_shifter_n77,
         dp_ex_stage_alu_shifter_n76, dp_ex_stage_alu_shifter_n75,
         dp_ex_stage_alu_shifter_n74, dp_ex_stage_alu_shifter_n73,
         dp_ex_stage_alu_shifter_n72, dp_ex_stage_alu_shifter_n71,
         dp_ex_stage_alu_shifter_n70, dp_ex_stage_alu_shifter_n69,
         dp_ex_stage_alu_shifter_n68, dp_ex_stage_alu_shifter_n67,
         dp_ex_stage_alu_shifter_n66, dp_ex_stage_alu_shifter_n65,
         dp_ex_stage_alu_shifter_n64, dp_ex_stage_alu_shifter_n63,
         dp_ex_stage_alu_shifter_n62, dp_ex_stage_alu_shifter_n61,
         dp_ex_stage_alu_shifter_n60, dp_ex_stage_alu_shifter_n59,
         dp_ex_stage_alu_shifter_n58, dp_ex_stage_alu_shifter_n57,
         dp_ex_stage_alu_shifter_n56, dp_ex_stage_alu_shifter_n55,
         dp_ex_stage_alu_shifter_n54, dp_ex_stage_alu_shifter_n53,
         dp_ex_stage_alu_shifter_n52, dp_ex_stage_alu_shifter_n51,
         dp_ex_stage_alu_shifter_n50, dp_ex_stage_alu_shifter_n49,
         dp_ex_stage_alu_shifter_n48, dp_ex_stage_alu_shifter_n47,
         dp_ex_stage_alu_shifter_n46, dp_ex_stage_alu_shifter_n45,
         dp_ex_stage_alu_shifter_n44, dp_ex_stage_alu_shifter_n43,
         dp_ex_stage_alu_shifter_n42, dp_ex_stage_alu_shifter_n41,
         dp_ex_stage_alu_shifter_n40, dp_ex_stage_alu_shifter_n39,
         dp_ex_stage_alu_shifter_n38, dp_ex_stage_alu_shifter_n37,
         dp_ex_stage_alu_shifter_n36, dp_ex_stage_alu_shifter_n35,
         dp_ex_stage_alu_shifter_n34, dp_ex_stage_alu_shifter_n33,
         dp_ex_stage_alu_shifter_n32, dp_ex_stage_alu_shifter_n31,
         dp_ex_stage_alu_shifter_n30, dp_ex_stage_alu_shifter_n29,
         dp_ex_stage_alu_shifter_n28, dp_ex_stage_alu_shifter_n27,
         dp_ex_stage_alu_shifter_n26, dp_ex_stage_alu_shifter_n25,
         dp_ex_stage_alu_shifter_n24, dp_ex_stage_alu_shifter_n23,
         dp_ex_stage_alu_shifter_n22, dp_ex_stage_alu_shifter_n21,
         dp_ex_stage_alu_shifter_N265, dp_ex_stage_alu_shifter_N264,
         dp_ex_stage_alu_shifter_N263, dp_ex_stage_alu_shifter_N262,
         dp_ex_stage_alu_shifter_N261, dp_ex_stage_alu_shifter_N260,
         dp_ex_stage_alu_shifter_N259, dp_ex_stage_alu_shifter_N258,
         dp_ex_stage_alu_shifter_N257, dp_ex_stage_alu_shifter_N256,
         dp_ex_stage_alu_shifter_N255, dp_ex_stage_alu_shifter_N254,
         dp_ex_stage_alu_shifter_N253, dp_ex_stage_alu_shifter_N252,
         dp_ex_stage_alu_shifter_N251, dp_ex_stage_alu_shifter_N250,
         dp_ex_stage_alu_shifter_N249, dp_ex_stage_alu_shifter_N248,
         dp_ex_stage_alu_shifter_N247, dp_ex_stage_alu_shifter_N246,
         dp_ex_stage_alu_shifter_N245, dp_ex_stage_alu_shifter_N244,
         dp_ex_stage_alu_shifter_N243, dp_ex_stage_alu_shifter_N242,
         dp_ex_stage_alu_shifter_N241, dp_ex_stage_alu_shifter_N240,
         dp_ex_stage_alu_shifter_N239, dp_ex_stage_alu_shifter_N238,
         dp_ex_stage_alu_shifter_N237, dp_ex_stage_alu_shifter_N236,
         dp_ex_stage_alu_shifter_N235, dp_ex_stage_alu_shifter_N234,
         dp_ex_stage_alu_shifter_N233, dp_ex_stage_alu_shifter_N232,
         dp_ex_stage_alu_shifter_N231, dp_ex_stage_alu_shifter_N230,
         dp_ex_stage_alu_shifter_N229, dp_ex_stage_alu_shifter_N228,
         dp_ex_stage_alu_shifter_N227, dp_ex_stage_alu_shifter_N226,
         dp_ex_stage_alu_shifter_N225, dp_ex_stage_alu_shifter_N224,
         dp_ex_stage_alu_shifter_N223, dp_ex_stage_alu_shifter_N222,
         dp_ex_stage_alu_shifter_N221, dp_ex_stage_alu_shifter_N220,
         dp_ex_stage_alu_shifter_N219, dp_ex_stage_alu_shifter_N218,
         dp_ex_stage_alu_shifter_N217, dp_ex_stage_alu_shifter_N216,
         dp_ex_stage_alu_shifter_N215, dp_ex_stage_alu_shifter_N214,
         dp_ex_stage_alu_shifter_N213, dp_ex_stage_alu_shifter_N212,
         dp_ex_stage_alu_shifter_N211, dp_ex_stage_alu_shifter_N210,
         dp_ex_stage_alu_shifter_N209, dp_ex_stage_alu_shifter_N208,
         dp_ex_stage_alu_shifter_N207, dp_ex_stage_alu_shifter_N206,
         dp_ex_stage_alu_shifter_N205, dp_ex_stage_alu_shifter_N204,
         dp_ex_stage_alu_shifter_N203, dp_ex_stage_alu_shifter_N202,
         dp_ex_stage_alu_shifter_N168, dp_ex_stage_alu_shifter_N167,
         dp_ex_stage_alu_shifter_N166, dp_ex_stage_alu_shifter_N165,
         dp_ex_stage_alu_shifter_N164, dp_ex_stage_alu_shifter_N163,
         dp_ex_stage_alu_shifter_N162, dp_ex_stage_alu_shifter_N161,
         dp_ex_stage_alu_shifter_N160, dp_ex_stage_alu_shifter_N159,
         dp_ex_stage_alu_shifter_N158, dp_ex_stage_alu_shifter_N157,
         dp_ex_stage_alu_shifter_N156, dp_ex_stage_alu_shifter_N155,
         dp_ex_stage_alu_shifter_N154, dp_ex_stage_alu_shifter_N153,
         dp_ex_stage_alu_shifter_N152, dp_ex_stage_alu_shifter_N151,
         dp_ex_stage_alu_shifter_N150, dp_ex_stage_alu_shifter_N149,
         dp_ex_stage_alu_shifter_N148, dp_ex_stage_alu_shifter_N147,
         dp_ex_stage_alu_shifter_N146, dp_ex_stage_alu_shifter_N145,
         dp_ex_stage_alu_shifter_N144, dp_ex_stage_alu_shifter_N143,
         dp_ex_stage_alu_shifter_N142, dp_ex_stage_alu_shifter_N141,
         dp_ex_stage_alu_shifter_N140, dp_ex_stage_alu_shifter_N139,
         dp_ex_stage_alu_shifter_N138, dp_ex_stage_alu_shifter_N137,
         dp_ex_stage_alu_shifter_N136, dp_ex_stage_alu_shifter_N135,
         dp_ex_stage_alu_shifter_N134, dp_ex_stage_alu_shifter_N133,
         dp_ex_stage_alu_shifter_N132, dp_ex_stage_alu_shifter_N131,
         dp_ex_stage_alu_shifter_N130, dp_ex_stage_alu_shifter_N129,
         dp_ex_stage_alu_shifter_N128, dp_ex_stage_alu_shifter_N127,
         dp_ex_stage_alu_shifter_N126, dp_ex_stage_alu_shifter_N125,
         dp_ex_stage_alu_shifter_N124, dp_ex_stage_alu_shifter_N123,
         dp_ex_stage_alu_shifter_N122, dp_ex_stage_alu_shifter_N121,
         dp_ex_stage_alu_shifter_N120, dp_ex_stage_alu_shifter_N119,
         dp_ex_stage_alu_shifter_N118, dp_ex_stage_alu_shifter_N117,
         dp_ex_stage_alu_shifter_N116, dp_ex_stage_alu_shifter_N115,
         dp_ex_stage_alu_shifter_N114, dp_ex_stage_alu_shifter_N113,
         dp_ex_stage_alu_shifter_N112, dp_ex_stage_alu_shifter_N111,
         dp_ex_stage_alu_shifter_N110, dp_ex_stage_alu_shifter_N109,
         dp_ex_stage_alu_shifter_N108, dp_ex_stage_alu_shifter_N107,
         dp_ex_stage_alu_shifter_N106, dp_ex_stage_alu_shifter_N105,
         dp_ex_stage_alu_shifter_N70, dp_ex_stage_alu_shifter_N69,
         dp_ex_stage_alu_shifter_N68, dp_ex_stage_alu_shifter_N67,
         dp_ex_stage_alu_shifter_N66, dp_ex_stage_alu_shifter_N65,
         dp_ex_stage_alu_shifter_N64, dp_ex_stage_alu_shifter_N63,
         dp_ex_stage_alu_shifter_N62, dp_ex_stage_alu_shifter_N61,
         dp_ex_stage_alu_shifter_N60, dp_ex_stage_alu_shifter_N59,
         dp_ex_stage_alu_shifter_N58, dp_ex_stage_alu_shifter_N57,
         dp_ex_stage_alu_shifter_N56, dp_ex_stage_alu_shifter_N55,
         dp_ex_stage_alu_shifter_N54, dp_ex_stage_alu_shifter_N53,
         dp_ex_stage_alu_shifter_N52, dp_ex_stage_alu_shifter_N51,
         dp_ex_stage_alu_shifter_N50, dp_ex_stage_alu_shifter_N49,
         dp_ex_stage_alu_shifter_N48, dp_ex_stage_alu_shifter_N47,
         dp_ex_stage_alu_shifter_N46, dp_ex_stage_alu_shifter_N45,
         dp_ex_stage_alu_shifter_N44, dp_ex_stage_alu_shifter_N43,
         dp_ex_stage_alu_shifter_N42, dp_ex_stage_alu_shifter_N41,
         dp_ex_stage_alu_shifter_N40, dp_ex_stage_alu_shifter_N39,
         dp_ex_stage_alu_shifter_N38, dp_ex_stage_alu_shifter_N37,
         dp_ex_stage_alu_shifter_N36, dp_ex_stage_alu_shifter_N35,
         dp_ex_stage_alu_shifter_N34, dp_ex_stage_alu_shifter_N33,
         dp_ex_stage_alu_shifter_N32, dp_ex_stage_alu_shifter_N31,
         dp_ex_stage_alu_shifter_N30, dp_ex_stage_alu_shifter_N29,
         dp_ex_stage_alu_shifter_N28, dp_ex_stage_alu_shifter_N27,
         dp_ex_stage_alu_shifter_N26, dp_ex_stage_alu_shifter_N25,
         dp_ex_stage_alu_shifter_N24, dp_ex_stage_alu_shifter_N23,
         dp_ex_stage_alu_shifter_N22, dp_ex_stage_alu_shifter_N21,
         dp_ex_stage_alu_shifter_N20, dp_ex_stage_alu_shifter_N19,
         dp_ex_stage_alu_shifter_N18, dp_ex_stage_alu_shifter_N17,
         dp_ex_stage_alu_shifter_N16, dp_ex_stage_alu_shifter_N15,
         dp_ex_stage_alu_shifter_N14, dp_ex_stage_alu_shifter_N13,
         dp_ex_stage_alu_shifter_N12, dp_ex_stage_alu_shifter_N11,
         dp_ex_stage_alu_shifter_N10, dp_ex_stage_alu_shifter_N9,
         dp_ex_stage_alu_shifter_N8, dp_ex_stage_alu_shifter_N7,
         dp_ex_stage_alu_shifter_sll_48_n34,
         dp_ex_stage_alu_shifter_sll_48_n33,
         dp_ex_stage_alu_shifter_sll_48_n32,
         dp_ex_stage_alu_shifter_sll_48_n31,
         dp_ex_stage_alu_shifter_sll_48_n30,
         dp_ex_stage_alu_shifter_sll_48_n29,
         dp_ex_stage_alu_shifter_sll_48_n28,
         dp_ex_stage_alu_shifter_sll_48_n27,
         dp_ex_stage_alu_shifter_sll_48_n26,
         dp_ex_stage_alu_shifter_sll_48_n25,
         dp_ex_stage_alu_shifter_sll_48_n24,
         dp_ex_stage_alu_shifter_sll_48_n23,
         dp_ex_stage_alu_shifter_sll_48_n22,
         dp_ex_stage_alu_shifter_sll_48_n21,
         dp_ex_stage_alu_shifter_sll_48_n20,
         dp_ex_stage_alu_shifter_sll_48_n19,
         dp_ex_stage_alu_shifter_sll_48_n18,
         dp_ex_stage_alu_shifter_sll_48_n17,
         dp_ex_stage_alu_shifter_sll_48_n16,
         dp_ex_stage_alu_shifter_sll_48_n15,
         dp_ex_stage_alu_shifter_sll_48_n14,
         dp_ex_stage_alu_shifter_sll_48_n13,
         dp_ex_stage_alu_shifter_sll_48_n12,
         dp_ex_stage_alu_shifter_sll_48_n11,
         dp_ex_stage_alu_shifter_sll_48_n10, dp_ex_stage_alu_shifter_sll_48_n9,
         dp_ex_stage_alu_shifter_sll_48_n8, dp_ex_stage_alu_shifter_sll_48_n7,
         dp_ex_stage_alu_shifter_sll_48_n6, dp_ex_stage_alu_shifter_sll_48_n5,
         dp_ex_stage_alu_shifter_sll_48_n4, dp_ex_stage_alu_shifter_sll_48_n3,
         dp_ex_stage_alu_shifter_sll_48_n2, dp_ex_stage_alu_shifter_sll_48_n1,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__8_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__9_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__10_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__11_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__12_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__13_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__14_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__15_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__16_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__17_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__18_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__19_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__20_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__21_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__22_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__23_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__24_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__25_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__26_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__27_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__28_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__29_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__30_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_4__31_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__0_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__1_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__2_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__3_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__4_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__5_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__6_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__7_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__8_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__9_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__10_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__11_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__12_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__13_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__14_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__15_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__16_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__17_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__18_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__19_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__20_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__21_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__22_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__23_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__24_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__25_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__26_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__27_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__28_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__29_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__30_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_3__31_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__0_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__1_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__2_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__3_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__4_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__5_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__6_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__7_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__8_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__9_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__10_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__11_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__12_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__13_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__14_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__15_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__16_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__17_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__18_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__19_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__20_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__21_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__22_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__23_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__24_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__25_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__26_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__27_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__28_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__29_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__30_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_2__31_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__0_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__1_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__2_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__3_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__4_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__5_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__6_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__7_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__8_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__9_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__10_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__11_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__12_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__13_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__14_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__15_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__16_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__17_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__18_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__19_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__20_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__21_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__22_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__23_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__24_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__25_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__26_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__27_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__28_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__29_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__30_,
         dp_ex_stage_alu_shifter_sll_48_ML_int_1__31_,
         dp_ex_stage_alu_shifter_sla_46_n193,
         dp_ex_stage_alu_shifter_sla_46_n192,
         dp_ex_stage_alu_shifter_sla_46_n191,
         dp_ex_stage_alu_shifter_sla_46_n190,
         dp_ex_stage_alu_shifter_sla_46_n189,
         dp_ex_stage_alu_shifter_sla_46_n188,
         dp_ex_stage_alu_shifter_sla_46_n187,
         dp_ex_stage_alu_shifter_sla_46_n186,
         dp_ex_stage_alu_shifter_sla_46_n185,
         dp_ex_stage_alu_shifter_sla_46_n184,
         dp_ex_stage_alu_shifter_sla_46_n183,
         dp_ex_stage_alu_shifter_sla_46_n182,
         dp_ex_stage_alu_shifter_sla_46_n181,
         dp_ex_stage_alu_shifter_sla_46_n180,
         dp_ex_stage_alu_shifter_sla_46_n179,
         dp_ex_stage_alu_shifter_sla_46_n178,
         dp_ex_stage_alu_shifter_sla_46_n177,
         dp_ex_stage_alu_shifter_sla_46_n176,
         dp_ex_stage_alu_shifter_sla_46_n175,
         dp_ex_stage_alu_shifter_sla_46_n174,
         dp_ex_stage_alu_shifter_sla_46_n173,
         dp_ex_stage_alu_shifter_sla_46_n172,
         dp_ex_stage_alu_shifter_sla_46_n171,
         dp_ex_stage_alu_shifter_sla_46_n170,
         dp_ex_stage_alu_shifter_sla_46_n169,
         dp_ex_stage_alu_shifter_sla_46_n168,
         dp_ex_stage_alu_shifter_sla_46_n167,
         dp_ex_stage_alu_shifter_sla_46_n166,
         dp_ex_stage_alu_shifter_sla_46_n165,
         dp_ex_stage_alu_shifter_sla_46_n164,
         dp_ex_stage_alu_shifter_sla_46_n163,
         dp_ex_stage_alu_shifter_sla_46_n162,
         dp_ex_stage_alu_shifter_sla_46_n161,
         dp_ex_stage_alu_shifter_sla_46_n160,
         dp_ex_stage_alu_shifter_sla_46_n159,
         dp_ex_stage_alu_shifter_sla_46_n158,
         dp_ex_stage_alu_shifter_sla_46_n157,
         dp_ex_stage_alu_shifter_sla_46_n156,
         dp_ex_stage_alu_shifter_sla_46_n155,
         dp_ex_stage_alu_shifter_sla_46_n154,
         dp_ex_stage_alu_shifter_sla_46_n153,
         dp_ex_stage_alu_shifter_sla_46_n152,
         dp_ex_stage_alu_shifter_sla_46_n151,
         dp_ex_stage_alu_shifter_sla_46_n150,
         dp_ex_stage_alu_shifter_sla_46_n149,
         dp_ex_stage_alu_shifter_sla_46_n148,
         dp_ex_stage_alu_shifter_sla_46_n147,
         dp_ex_stage_alu_shifter_sla_46_n146,
         dp_ex_stage_alu_shifter_sla_46_n145,
         dp_ex_stage_alu_shifter_sla_46_n144,
         dp_ex_stage_alu_shifter_sla_46_n143,
         dp_ex_stage_alu_shifter_sla_46_n142,
         dp_ex_stage_alu_shifter_sla_46_n141,
         dp_ex_stage_alu_shifter_sla_46_n140,
         dp_ex_stage_alu_shifter_sla_46_n139,
         dp_ex_stage_alu_shifter_sla_46_n138,
         dp_ex_stage_alu_shifter_sla_46_n137,
         dp_ex_stage_alu_shifter_sla_46_n136,
         dp_ex_stage_alu_shifter_sla_46_n135,
         dp_ex_stage_alu_shifter_sla_46_n134,
         dp_ex_stage_alu_shifter_sla_46_n133,
         dp_ex_stage_alu_shifter_sla_46_n132,
         dp_ex_stage_alu_shifter_sla_46_n131,
         dp_ex_stage_alu_shifter_sla_46_n130,
         dp_ex_stage_alu_shifter_sla_46_n129,
         dp_ex_stage_alu_shifter_sla_46_n128,
         dp_ex_stage_alu_shifter_sla_46_n127,
         dp_ex_stage_alu_shifter_sla_46_n126,
         dp_ex_stage_alu_shifter_sla_46_n125,
         dp_ex_stage_alu_shifter_sla_46_n124,
         dp_ex_stage_alu_shifter_sla_46_n123,
         dp_ex_stage_alu_shifter_sla_46_n122,
         dp_ex_stage_alu_shifter_sla_46_n121,
         dp_ex_stage_alu_shifter_sla_46_n120,
         dp_ex_stage_alu_shifter_sla_46_n119,
         dp_ex_stage_alu_shifter_sla_46_n118,
         dp_ex_stage_alu_shifter_sla_46_n117,
         dp_ex_stage_alu_shifter_sla_46_n116,
         dp_ex_stage_alu_shifter_sla_46_n115,
         dp_ex_stage_alu_shifter_sla_46_n114,
         dp_ex_stage_alu_shifter_sla_46_n113,
         dp_ex_stage_alu_shifter_sla_46_n112,
         dp_ex_stage_alu_shifter_sla_46_n111,
         dp_ex_stage_alu_shifter_sla_46_n110,
         dp_ex_stage_alu_shifter_sla_46_n109,
         dp_ex_stage_alu_shifter_sla_46_n108,
         dp_ex_stage_alu_shifter_sla_46_n107,
         dp_ex_stage_alu_shifter_sla_46_n106,
         dp_ex_stage_alu_shifter_sla_46_n105,
         dp_ex_stage_alu_shifter_sla_46_n104,
         dp_ex_stage_alu_shifter_sla_46_n103,
         dp_ex_stage_alu_shifter_sla_46_n102,
         dp_ex_stage_alu_shifter_sla_46_n101,
         dp_ex_stage_alu_shifter_sla_46_n100,
         dp_ex_stage_alu_shifter_sla_46_n99,
         dp_ex_stage_alu_shifter_sla_46_n98,
         dp_ex_stage_alu_shifter_sla_46_n97,
         dp_ex_stage_alu_shifter_sla_46_n96,
         dp_ex_stage_alu_shifter_sla_46_n95,
         dp_ex_stage_alu_shifter_sla_46_n94,
         dp_ex_stage_alu_shifter_sla_46_n93,
         dp_ex_stage_alu_shifter_sla_46_n92,
         dp_ex_stage_alu_shifter_sla_46_n91,
         dp_ex_stage_alu_shifter_sla_46_n90,
         dp_ex_stage_alu_shifter_sla_46_n89,
         dp_ex_stage_alu_shifter_sla_46_n88,
         dp_ex_stage_alu_shifter_sla_46_n87,
         dp_ex_stage_alu_shifter_sla_46_n86,
         dp_ex_stage_alu_shifter_sla_46_n85,
         dp_ex_stage_alu_shifter_sla_46_n84,
         dp_ex_stage_alu_shifter_sla_46_n83,
         dp_ex_stage_alu_shifter_sla_46_n82,
         dp_ex_stage_alu_shifter_sla_46_n81,
         dp_ex_stage_alu_shifter_sla_46_n80,
         dp_ex_stage_alu_shifter_sla_46_n79,
         dp_ex_stage_alu_shifter_sla_46_n78,
         dp_ex_stage_alu_shifter_sla_46_n77,
         dp_ex_stage_alu_shifter_sla_46_n76,
         dp_ex_stage_alu_shifter_sla_46_n75,
         dp_ex_stage_alu_shifter_sla_46_n74,
         dp_ex_stage_alu_shifter_sla_46_n73,
         dp_ex_stage_alu_shifter_sla_46_n72,
         dp_ex_stage_alu_shifter_sla_46_n71,
         dp_ex_stage_alu_shifter_sla_46_n70,
         dp_ex_stage_alu_shifter_sla_46_n69,
         dp_ex_stage_alu_shifter_sla_46_n68,
         dp_ex_stage_alu_shifter_sla_46_n67,
         dp_ex_stage_alu_shifter_sla_46_n66,
         dp_ex_stage_alu_shifter_sla_46_n65,
         dp_ex_stage_alu_shifter_sla_46_n64,
         dp_ex_stage_alu_shifter_sla_46_n63,
         dp_ex_stage_alu_shifter_sla_46_n62,
         dp_ex_stage_alu_shifter_sla_46_n61,
         dp_ex_stage_alu_shifter_sla_46_n60,
         dp_ex_stage_alu_shifter_sla_46_n59,
         dp_ex_stage_alu_shifter_sla_46_n58,
         dp_ex_stage_alu_shifter_sla_46_n57,
         dp_ex_stage_alu_shifter_sla_46_n56,
         dp_ex_stage_alu_shifter_sla_46_n55,
         dp_ex_stage_alu_shifter_sla_46_n54,
         dp_ex_stage_alu_shifter_sla_46_n53,
         dp_ex_stage_alu_shifter_sla_46_n52,
         dp_ex_stage_alu_shifter_sla_46_n51,
         dp_ex_stage_alu_shifter_sla_46_n50,
         dp_ex_stage_alu_shifter_sla_46_n49,
         dp_ex_stage_alu_shifter_sla_46_n48,
         dp_ex_stage_alu_shifter_sla_46_n47,
         dp_ex_stage_alu_shifter_sla_46_n46,
         dp_ex_stage_alu_shifter_sla_46_n45,
         dp_ex_stage_alu_shifter_sla_46_n44,
         dp_ex_stage_alu_shifter_sla_46_n43,
         dp_ex_stage_alu_shifter_sla_46_n42,
         dp_ex_stage_alu_shifter_sla_46_n41,
         dp_ex_stage_alu_shifter_sla_46_n40,
         dp_ex_stage_alu_shifter_sla_46_n39,
         dp_ex_stage_alu_shifter_sla_46_n38,
         dp_ex_stage_alu_shifter_sla_46_n37,
         dp_ex_stage_alu_shifter_sla_46_n36,
         dp_ex_stage_alu_shifter_sla_46_n35,
         dp_ex_stage_alu_shifter_sla_46_n34,
         dp_ex_stage_alu_shifter_sla_46_n33,
         dp_ex_stage_alu_shifter_sla_46_n32,
         dp_ex_stage_alu_shifter_sla_46_n31,
         dp_ex_stage_alu_shifter_sla_46_n30,
         dp_ex_stage_alu_shifter_sla_46_n29,
         dp_ex_stage_alu_shifter_sla_46_n28,
         dp_ex_stage_alu_shifter_sla_46_n27,
         dp_ex_stage_alu_shifter_sla_46_n26,
         dp_ex_stage_alu_shifter_sla_46_n25,
         dp_ex_stage_alu_shifter_sla_46_n24,
         dp_ex_stage_alu_shifter_sla_46_n23,
         dp_ex_stage_alu_shifter_sla_46_n22,
         dp_ex_stage_alu_shifter_sla_46_n21,
         dp_ex_stage_alu_shifter_sla_46_n20,
         dp_ex_stage_alu_shifter_sla_46_n19,
         dp_ex_stage_alu_shifter_sla_46_n18,
         dp_ex_stage_alu_shifter_sla_46_n17,
         dp_ex_stage_alu_shifter_sla_46_n16,
         dp_ex_stage_alu_shifter_sla_46_n15,
         dp_ex_stage_alu_shifter_sla_46_n14,
         dp_ex_stage_alu_shifter_sla_46_n13,
         dp_ex_stage_alu_shifter_sla_46_n12,
         dp_ex_stage_alu_shifter_sla_46_n11,
         dp_ex_stage_alu_shifter_sla_46_n10, dp_ex_stage_alu_shifter_sla_46_n9,
         dp_ex_stage_alu_shifter_sla_46_n8, dp_ex_stage_alu_shifter_sla_46_n7,
         dp_ex_stage_alu_shifter_sla_46_n6, dp_ex_stage_alu_shifter_sla_46_n5,
         dp_ex_stage_alu_shifter_sla_46_n4, dp_ex_stage_alu_shifter_sla_46_n3,
         dp_ex_stage_alu_shifter_sla_46_n2, dp_ex_stage_alu_shifter_sla_46_n1,
         dp_ex_stage_alu_shifter_srl_41_n189,
         dp_ex_stage_alu_shifter_srl_41_n188,
         dp_ex_stage_alu_shifter_srl_41_n187,
         dp_ex_stage_alu_shifter_srl_41_n186,
         dp_ex_stage_alu_shifter_srl_41_n185,
         dp_ex_stage_alu_shifter_srl_41_n184,
         dp_ex_stage_alu_shifter_srl_41_n183,
         dp_ex_stage_alu_shifter_srl_41_n182,
         dp_ex_stage_alu_shifter_srl_41_n181,
         dp_ex_stage_alu_shifter_srl_41_n180,
         dp_ex_stage_alu_shifter_srl_41_n179,
         dp_ex_stage_alu_shifter_srl_41_n178,
         dp_ex_stage_alu_shifter_srl_41_n177,
         dp_ex_stage_alu_shifter_srl_41_n176,
         dp_ex_stage_alu_shifter_srl_41_n175,
         dp_ex_stage_alu_shifter_srl_41_n174,
         dp_ex_stage_alu_shifter_srl_41_n173,
         dp_ex_stage_alu_shifter_srl_41_n172,
         dp_ex_stage_alu_shifter_srl_41_n171,
         dp_ex_stage_alu_shifter_srl_41_n170,
         dp_ex_stage_alu_shifter_srl_41_n169,
         dp_ex_stage_alu_shifter_srl_41_n168,
         dp_ex_stage_alu_shifter_srl_41_n167,
         dp_ex_stage_alu_shifter_srl_41_n166,
         dp_ex_stage_alu_shifter_srl_41_n165,
         dp_ex_stage_alu_shifter_srl_41_n164,
         dp_ex_stage_alu_shifter_srl_41_n163,
         dp_ex_stage_alu_shifter_srl_41_n162,
         dp_ex_stage_alu_shifter_srl_41_n161,
         dp_ex_stage_alu_shifter_srl_41_n160,
         dp_ex_stage_alu_shifter_srl_41_n159,
         dp_ex_stage_alu_shifter_srl_41_n158,
         dp_ex_stage_alu_shifter_srl_41_n157,
         dp_ex_stage_alu_shifter_srl_41_n156,
         dp_ex_stage_alu_shifter_srl_41_n155,
         dp_ex_stage_alu_shifter_srl_41_n154,
         dp_ex_stage_alu_shifter_srl_41_n153,
         dp_ex_stage_alu_shifter_srl_41_n152,
         dp_ex_stage_alu_shifter_srl_41_n151,
         dp_ex_stage_alu_shifter_srl_41_n150,
         dp_ex_stage_alu_shifter_srl_41_n149,
         dp_ex_stage_alu_shifter_srl_41_n148,
         dp_ex_stage_alu_shifter_srl_41_n147,
         dp_ex_stage_alu_shifter_srl_41_n146,
         dp_ex_stage_alu_shifter_srl_41_n145,
         dp_ex_stage_alu_shifter_srl_41_n144,
         dp_ex_stage_alu_shifter_srl_41_n143,
         dp_ex_stage_alu_shifter_srl_41_n142,
         dp_ex_stage_alu_shifter_srl_41_n141,
         dp_ex_stage_alu_shifter_srl_41_n140,
         dp_ex_stage_alu_shifter_srl_41_n139,
         dp_ex_stage_alu_shifter_srl_41_n138,
         dp_ex_stage_alu_shifter_srl_41_n137,
         dp_ex_stage_alu_shifter_srl_41_n136,
         dp_ex_stage_alu_shifter_srl_41_n135,
         dp_ex_stage_alu_shifter_srl_41_n134,
         dp_ex_stage_alu_shifter_srl_41_n133,
         dp_ex_stage_alu_shifter_srl_41_n132,
         dp_ex_stage_alu_shifter_srl_41_n131,
         dp_ex_stage_alu_shifter_srl_41_n130,
         dp_ex_stage_alu_shifter_srl_41_n129,
         dp_ex_stage_alu_shifter_srl_41_n128,
         dp_ex_stage_alu_shifter_srl_41_n127,
         dp_ex_stage_alu_shifter_srl_41_n126,
         dp_ex_stage_alu_shifter_srl_41_n125,
         dp_ex_stage_alu_shifter_srl_41_n124,
         dp_ex_stage_alu_shifter_srl_41_n123,
         dp_ex_stage_alu_shifter_srl_41_n122,
         dp_ex_stage_alu_shifter_srl_41_n121,
         dp_ex_stage_alu_shifter_srl_41_n120,
         dp_ex_stage_alu_shifter_srl_41_n119,
         dp_ex_stage_alu_shifter_srl_41_n118,
         dp_ex_stage_alu_shifter_srl_41_n117,
         dp_ex_stage_alu_shifter_srl_41_n116,
         dp_ex_stage_alu_shifter_srl_41_n115,
         dp_ex_stage_alu_shifter_srl_41_n114,
         dp_ex_stage_alu_shifter_srl_41_n113,
         dp_ex_stage_alu_shifter_srl_41_n112,
         dp_ex_stage_alu_shifter_srl_41_n111,
         dp_ex_stage_alu_shifter_srl_41_n110,
         dp_ex_stage_alu_shifter_srl_41_n109,
         dp_ex_stage_alu_shifter_srl_41_n108,
         dp_ex_stage_alu_shifter_srl_41_n107,
         dp_ex_stage_alu_shifter_srl_41_n106,
         dp_ex_stage_alu_shifter_srl_41_n105,
         dp_ex_stage_alu_shifter_srl_41_n104,
         dp_ex_stage_alu_shifter_srl_41_n103,
         dp_ex_stage_alu_shifter_srl_41_n102,
         dp_ex_stage_alu_shifter_srl_41_n101,
         dp_ex_stage_alu_shifter_srl_41_n100,
         dp_ex_stage_alu_shifter_srl_41_n99,
         dp_ex_stage_alu_shifter_srl_41_n98,
         dp_ex_stage_alu_shifter_srl_41_n97,
         dp_ex_stage_alu_shifter_srl_41_n96,
         dp_ex_stage_alu_shifter_srl_41_n95,
         dp_ex_stage_alu_shifter_srl_41_n94,
         dp_ex_stage_alu_shifter_srl_41_n93,
         dp_ex_stage_alu_shifter_srl_41_n92,
         dp_ex_stage_alu_shifter_srl_41_n91,
         dp_ex_stage_alu_shifter_srl_41_n90,
         dp_ex_stage_alu_shifter_srl_41_n89,
         dp_ex_stage_alu_shifter_srl_41_n88,
         dp_ex_stage_alu_shifter_srl_41_n87,
         dp_ex_stage_alu_shifter_srl_41_n86,
         dp_ex_stage_alu_shifter_srl_41_n85,
         dp_ex_stage_alu_shifter_srl_41_n84,
         dp_ex_stage_alu_shifter_srl_41_n83,
         dp_ex_stage_alu_shifter_srl_41_n82,
         dp_ex_stage_alu_shifter_srl_41_n81,
         dp_ex_stage_alu_shifter_srl_41_n80,
         dp_ex_stage_alu_shifter_srl_41_n79,
         dp_ex_stage_alu_shifter_srl_41_n78,
         dp_ex_stage_alu_shifter_srl_41_n77,
         dp_ex_stage_alu_shifter_srl_41_n76,
         dp_ex_stage_alu_shifter_srl_41_n75,
         dp_ex_stage_alu_shifter_srl_41_n74,
         dp_ex_stage_alu_shifter_srl_41_n73,
         dp_ex_stage_alu_shifter_srl_41_n72,
         dp_ex_stage_alu_shifter_srl_41_n71,
         dp_ex_stage_alu_shifter_srl_41_n70,
         dp_ex_stage_alu_shifter_srl_41_n69,
         dp_ex_stage_alu_shifter_srl_41_n68,
         dp_ex_stage_alu_shifter_srl_41_n67,
         dp_ex_stage_alu_shifter_srl_41_n66,
         dp_ex_stage_alu_shifter_srl_41_n65,
         dp_ex_stage_alu_shifter_srl_41_n64,
         dp_ex_stage_alu_shifter_srl_41_n63,
         dp_ex_stage_alu_shifter_srl_41_n62,
         dp_ex_stage_alu_shifter_srl_41_n60,
         dp_ex_stage_alu_shifter_srl_41_n59,
         dp_ex_stage_alu_shifter_srl_41_n58,
         dp_ex_stage_alu_shifter_srl_41_n57,
         dp_ex_stage_alu_shifter_srl_41_n56,
         dp_ex_stage_alu_shifter_srl_41_n55,
         dp_ex_stage_alu_shifter_srl_41_n54,
         dp_ex_stage_alu_shifter_srl_41_n53,
         dp_ex_stage_alu_shifter_srl_41_n52,
         dp_ex_stage_alu_shifter_srl_41_n51,
         dp_ex_stage_alu_shifter_srl_41_n50,
         dp_ex_stage_alu_shifter_srl_41_n49,
         dp_ex_stage_alu_shifter_srl_41_n48,
         dp_ex_stage_alu_shifter_srl_41_n47,
         dp_ex_stage_alu_shifter_srl_41_n46,
         dp_ex_stage_alu_shifter_srl_41_n45,
         dp_ex_stage_alu_shifter_srl_41_n44,
         dp_ex_stage_alu_shifter_srl_41_n43,
         dp_ex_stage_alu_shifter_srl_41_n42,
         dp_ex_stage_alu_shifter_srl_41_n41,
         dp_ex_stage_alu_shifter_srl_41_n40,
         dp_ex_stage_alu_shifter_srl_41_n39,
         dp_ex_stage_alu_shifter_srl_41_n38,
         dp_ex_stage_alu_shifter_srl_41_n37,
         dp_ex_stage_alu_shifter_srl_41_n36,
         dp_ex_stage_alu_shifter_srl_41_n35,
         dp_ex_stage_alu_shifter_srl_41_n34,
         dp_ex_stage_alu_shifter_srl_41_n33,
         dp_ex_stage_alu_shifter_srl_41_n32,
         dp_ex_stage_alu_shifter_srl_41_n31,
         dp_ex_stage_alu_shifter_srl_41_n30,
         dp_ex_stage_alu_shifter_srl_41_n29,
         dp_ex_stage_alu_shifter_srl_41_n28,
         dp_ex_stage_alu_shifter_srl_41_n27,
         dp_ex_stage_alu_shifter_srl_41_n26,
         dp_ex_stage_alu_shifter_srl_41_n25,
         dp_ex_stage_alu_shifter_srl_41_n24,
         dp_ex_stage_alu_shifter_srl_41_n23,
         dp_ex_stage_alu_shifter_srl_41_n22,
         dp_ex_stage_alu_shifter_srl_41_n21,
         dp_ex_stage_alu_shifter_srl_41_n20,
         dp_ex_stage_alu_shifter_srl_41_n19,
         dp_ex_stage_alu_shifter_srl_41_n18,
         dp_ex_stage_alu_shifter_srl_41_n17,
         dp_ex_stage_alu_shifter_srl_41_n16,
         dp_ex_stage_alu_shifter_srl_41_n15,
         dp_ex_stage_alu_shifter_srl_41_n14,
         dp_ex_stage_alu_shifter_srl_41_n13,
         dp_ex_stage_alu_shifter_srl_41_n12,
         dp_ex_stage_alu_shifter_srl_41_n11,
         dp_ex_stage_alu_shifter_srl_41_n10, dp_ex_stage_alu_shifter_srl_41_n9,
         dp_ex_stage_alu_shifter_srl_41_n8, dp_ex_stage_alu_shifter_srl_41_n7,
         dp_ex_stage_alu_shifter_srl_41_n6, dp_ex_stage_alu_shifter_srl_41_n5,
         dp_ex_stage_alu_shifter_srl_41_n4, dp_ex_stage_alu_shifter_srl_41_n3,
         dp_ex_stage_alu_shifter_srl_41_n2, dp_ex_stage_alu_shifter_srl_41_n1,
         dp_ex_stage_alu_shifter_sra_39_n193,
         dp_ex_stage_alu_shifter_sra_39_n192,
         dp_ex_stage_alu_shifter_sra_39_n191,
         dp_ex_stage_alu_shifter_sra_39_n190,
         dp_ex_stage_alu_shifter_sra_39_n189,
         dp_ex_stage_alu_shifter_sra_39_n188,
         dp_ex_stage_alu_shifter_sra_39_n187,
         dp_ex_stage_alu_shifter_sra_39_n186,
         dp_ex_stage_alu_shifter_sra_39_n185,
         dp_ex_stage_alu_shifter_sra_39_n184,
         dp_ex_stage_alu_shifter_sra_39_n183,
         dp_ex_stage_alu_shifter_sra_39_n182,
         dp_ex_stage_alu_shifter_sra_39_n181,
         dp_ex_stage_alu_shifter_sra_39_n180,
         dp_ex_stage_alu_shifter_sra_39_n179,
         dp_ex_stage_alu_shifter_sra_39_n178,
         dp_ex_stage_alu_shifter_sra_39_n177,
         dp_ex_stage_alu_shifter_sra_39_n176,
         dp_ex_stage_alu_shifter_sra_39_n175,
         dp_ex_stage_alu_shifter_sra_39_n174,
         dp_ex_stage_alu_shifter_sra_39_n173,
         dp_ex_stage_alu_shifter_sra_39_n172,
         dp_ex_stage_alu_shifter_sra_39_n171,
         dp_ex_stage_alu_shifter_sra_39_n170,
         dp_ex_stage_alu_shifter_sra_39_n169,
         dp_ex_stage_alu_shifter_sra_39_n168,
         dp_ex_stage_alu_shifter_sra_39_n167,
         dp_ex_stage_alu_shifter_sra_39_n166,
         dp_ex_stage_alu_shifter_sra_39_n165,
         dp_ex_stage_alu_shifter_sra_39_n164,
         dp_ex_stage_alu_shifter_sra_39_n163,
         dp_ex_stage_alu_shifter_sra_39_n162,
         dp_ex_stage_alu_shifter_sra_39_n161,
         dp_ex_stage_alu_shifter_sra_39_n160,
         dp_ex_stage_alu_shifter_sra_39_n159,
         dp_ex_stage_alu_shifter_sra_39_n158,
         dp_ex_stage_alu_shifter_sra_39_n157,
         dp_ex_stage_alu_shifter_sra_39_n156,
         dp_ex_stage_alu_shifter_sra_39_n155,
         dp_ex_stage_alu_shifter_sra_39_n154,
         dp_ex_stage_alu_shifter_sra_39_n153,
         dp_ex_stage_alu_shifter_sra_39_n152,
         dp_ex_stage_alu_shifter_sra_39_n151,
         dp_ex_stage_alu_shifter_sra_39_n150,
         dp_ex_stage_alu_shifter_sra_39_n149,
         dp_ex_stage_alu_shifter_sra_39_n148,
         dp_ex_stage_alu_shifter_sra_39_n147,
         dp_ex_stage_alu_shifter_sra_39_n146,
         dp_ex_stage_alu_shifter_sra_39_n145,
         dp_ex_stage_alu_shifter_sra_39_n144,
         dp_ex_stage_alu_shifter_sra_39_n143,
         dp_ex_stage_alu_shifter_sra_39_n142,
         dp_ex_stage_alu_shifter_sra_39_n141,
         dp_ex_stage_alu_shifter_sra_39_n140,
         dp_ex_stage_alu_shifter_sra_39_n139,
         dp_ex_stage_alu_shifter_sra_39_n138,
         dp_ex_stage_alu_shifter_sra_39_n137,
         dp_ex_stage_alu_shifter_sra_39_n136,
         dp_ex_stage_alu_shifter_sra_39_n135,
         dp_ex_stage_alu_shifter_sra_39_n134,
         dp_ex_stage_alu_shifter_sra_39_n133,
         dp_ex_stage_alu_shifter_sra_39_n132,
         dp_ex_stage_alu_shifter_sra_39_n131,
         dp_ex_stage_alu_shifter_sra_39_n130,
         dp_ex_stage_alu_shifter_sra_39_n129,
         dp_ex_stage_alu_shifter_sra_39_n128,
         dp_ex_stage_alu_shifter_sra_39_n127,
         dp_ex_stage_alu_shifter_sra_39_n126,
         dp_ex_stage_alu_shifter_sra_39_n125,
         dp_ex_stage_alu_shifter_sra_39_n124,
         dp_ex_stage_alu_shifter_sra_39_n123,
         dp_ex_stage_alu_shifter_sra_39_n122,
         dp_ex_stage_alu_shifter_sra_39_n121,
         dp_ex_stage_alu_shifter_sra_39_n120,
         dp_ex_stage_alu_shifter_sra_39_n119,
         dp_ex_stage_alu_shifter_sra_39_n118,
         dp_ex_stage_alu_shifter_sra_39_n117,
         dp_ex_stage_alu_shifter_sra_39_n116,
         dp_ex_stage_alu_shifter_sra_39_n115,
         dp_ex_stage_alu_shifter_sra_39_n114,
         dp_ex_stage_alu_shifter_sra_39_n113,
         dp_ex_stage_alu_shifter_sra_39_n112,
         dp_ex_stage_alu_shifter_sra_39_n111,
         dp_ex_stage_alu_shifter_sra_39_n110,
         dp_ex_stage_alu_shifter_sra_39_n109,
         dp_ex_stage_alu_shifter_sra_39_n108,
         dp_ex_stage_alu_shifter_sra_39_n107,
         dp_ex_stage_alu_shifter_sra_39_n106,
         dp_ex_stage_alu_shifter_sra_39_n105,
         dp_ex_stage_alu_shifter_sra_39_n104,
         dp_ex_stage_alu_shifter_sra_39_n103,
         dp_ex_stage_alu_shifter_sra_39_n102,
         dp_ex_stage_alu_shifter_sra_39_n101,
         dp_ex_stage_alu_shifter_sra_39_n100,
         dp_ex_stage_alu_shifter_sra_39_n99,
         dp_ex_stage_alu_shifter_sra_39_n98,
         dp_ex_stage_alu_shifter_sra_39_n97,
         dp_ex_stage_alu_shifter_sra_39_n96,
         dp_ex_stage_alu_shifter_sra_39_n95,
         dp_ex_stage_alu_shifter_sra_39_n94,
         dp_ex_stage_alu_shifter_sra_39_n93,
         dp_ex_stage_alu_shifter_sra_39_n92,
         dp_ex_stage_alu_shifter_sra_39_n91,
         dp_ex_stage_alu_shifter_sra_39_n90,
         dp_ex_stage_alu_shifter_sra_39_n89,
         dp_ex_stage_alu_shifter_sra_39_n88,
         dp_ex_stage_alu_shifter_sra_39_n87,
         dp_ex_stage_alu_shifter_sra_39_n86,
         dp_ex_stage_alu_shifter_sra_39_n85,
         dp_ex_stage_alu_shifter_sra_39_n84,
         dp_ex_stage_alu_shifter_sra_39_n83,
         dp_ex_stage_alu_shifter_sra_39_n82,
         dp_ex_stage_alu_shifter_sra_39_n81,
         dp_ex_stage_alu_shifter_sra_39_n80,
         dp_ex_stage_alu_shifter_sra_39_n79,
         dp_ex_stage_alu_shifter_sra_39_n78,
         dp_ex_stage_alu_shifter_sra_39_n77,
         dp_ex_stage_alu_shifter_sra_39_n76,
         dp_ex_stage_alu_shifter_sra_39_n75,
         dp_ex_stage_alu_shifter_sra_39_n74,
         dp_ex_stage_alu_shifter_sra_39_n73,
         dp_ex_stage_alu_shifter_sra_39_n72,
         dp_ex_stage_alu_shifter_sra_39_n71,
         dp_ex_stage_alu_shifter_sra_39_n70,
         dp_ex_stage_alu_shifter_sra_39_n69,
         dp_ex_stage_alu_shifter_sra_39_n68,
         dp_ex_stage_alu_shifter_sra_39_n67,
         dp_ex_stage_alu_shifter_sra_39_n66,
         dp_ex_stage_alu_shifter_sra_39_n65,
         dp_ex_stage_alu_shifter_sra_39_n64,
         dp_ex_stage_alu_shifter_sra_39_n63,
         dp_ex_stage_alu_shifter_sra_39_n62,
         dp_ex_stage_alu_shifter_sra_39_n61,
         dp_ex_stage_alu_shifter_sra_39_n60,
         dp_ex_stage_alu_shifter_sra_39_n59,
         dp_ex_stage_alu_shifter_sra_39_n58,
         dp_ex_stage_alu_shifter_sra_39_n57,
         dp_ex_stage_alu_shifter_sra_39_n56,
         dp_ex_stage_alu_shifter_sra_39_n55,
         dp_ex_stage_alu_shifter_sra_39_n54,
         dp_ex_stage_alu_shifter_sra_39_n53,
         dp_ex_stage_alu_shifter_sra_39_n52,
         dp_ex_stage_alu_shifter_sra_39_n51,
         dp_ex_stage_alu_shifter_sra_39_n50,
         dp_ex_stage_alu_shifter_sra_39_n49,
         dp_ex_stage_alu_shifter_sra_39_n48,
         dp_ex_stage_alu_shifter_sra_39_n47,
         dp_ex_stage_alu_shifter_sra_39_n46,
         dp_ex_stage_alu_shifter_sra_39_n45,
         dp_ex_stage_alu_shifter_sra_39_n43,
         dp_ex_stage_alu_shifter_sra_39_n42,
         dp_ex_stage_alu_shifter_sra_39_n41,
         dp_ex_stage_alu_shifter_sra_39_n40,
         dp_ex_stage_alu_shifter_sra_39_n39,
         dp_ex_stage_alu_shifter_sra_39_n38,
         dp_ex_stage_alu_shifter_sra_39_n37,
         dp_ex_stage_alu_shifter_sra_39_n36,
         dp_ex_stage_alu_shifter_sra_39_n35,
         dp_ex_stage_alu_shifter_sra_39_n34,
         dp_ex_stage_alu_shifter_sra_39_n33,
         dp_ex_stage_alu_shifter_sra_39_n32,
         dp_ex_stage_alu_shifter_sra_39_n31,
         dp_ex_stage_alu_shifter_sra_39_n30,
         dp_ex_stage_alu_shifter_sra_39_n29,
         dp_ex_stage_alu_shifter_sra_39_n28,
         dp_ex_stage_alu_shifter_sra_39_n27,
         dp_ex_stage_alu_shifter_sra_39_n26,
         dp_ex_stage_alu_shifter_sra_39_n25,
         dp_ex_stage_alu_shifter_sra_39_n24,
         dp_ex_stage_alu_shifter_sra_39_n23,
         dp_ex_stage_alu_shifter_sra_39_n22,
         dp_ex_stage_alu_shifter_sra_39_n21,
         dp_ex_stage_alu_shifter_sra_39_n20,
         dp_ex_stage_alu_shifter_sra_39_n19,
         dp_ex_stage_alu_shifter_sra_39_n18,
         dp_ex_stage_alu_shifter_sra_39_n17,
         dp_ex_stage_alu_shifter_sra_39_n16,
         dp_ex_stage_alu_shifter_sra_39_n15,
         dp_ex_stage_alu_shifter_sra_39_n14,
         dp_ex_stage_alu_shifter_sra_39_n13,
         dp_ex_stage_alu_shifter_sra_39_n12,
         dp_ex_stage_alu_shifter_sra_39_n11,
         dp_ex_stage_alu_shifter_sra_39_n10, dp_ex_stage_alu_shifter_sra_39_n9,
         dp_ex_stage_alu_shifter_sra_39_n8, dp_ex_stage_alu_shifter_sra_39_n7,
         dp_ex_stage_alu_shifter_sra_39_n6, dp_ex_stage_alu_shifter_sra_39_n5,
         dp_ex_stage_alu_shifter_sra_39_n4, dp_ex_stage_alu_shifter_sra_39_n3,
         dp_ex_stage_alu_shifter_sra_39_n2, dp_ex_stage_alu_shifter_sra_39_n1,
         dp_ex_stage_alu_shifter_rol_32_n15,
         dp_ex_stage_alu_shifter_rol_32_n14,
         dp_ex_stage_alu_shifter_rol_32_n13,
         dp_ex_stage_alu_shifter_rol_32_n12,
         dp_ex_stage_alu_shifter_rol_32_n11,
         dp_ex_stage_alu_shifter_rol_32_n10, dp_ex_stage_alu_shifter_rol_32_n9,
         dp_ex_stage_alu_shifter_rol_32_n8, dp_ex_stage_alu_shifter_rol_32_n7,
         dp_ex_stage_alu_shifter_rol_32_n6, dp_ex_stage_alu_shifter_rol_32_n5,
         dp_ex_stage_alu_shifter_rol_32_n4, dp_ex_stage_alu_shifter_rol_32_n3,
         dp_ex_stage_alu_shifter_rol_32_n2, dp_ex_stage_alu_shifter_rol_32_n1,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__0_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__1_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__2_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__3_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__4_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__5_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__6_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__7_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__8_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__9_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__10_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__11_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__12_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__13_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__14_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__15_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__16_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__17_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__18_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__19_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__20_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__21_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__22_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__23_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__24_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__25_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__26_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__27_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__28_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__29_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__30_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_4__31_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__0_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__1_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__2_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__3_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__4_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__5_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__6_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__7_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__8_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__9_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__10_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__11_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__12_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__13_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__14_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__15_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__16_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__17_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__18_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__19_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__20_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__21_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__22_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__23_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__24_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__25_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__26_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__27_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__28_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__29_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__30_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_3__31_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__0_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__1_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__2_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__3_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__4_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__5_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__6_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__7_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__8_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__9_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__10_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__11_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__12_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__13_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__14_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__15_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__16_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__17_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__18_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__19_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__20_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__21_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__22_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__23_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__24_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__25_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__26_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__27_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__28_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__29_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__30_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_2__31_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__0_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__1_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__2_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__3_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__4_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__5_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__6_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__7_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__8_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__9_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__10_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__11_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__12_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__13_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__14_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__15_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__16_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__17_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__18_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__19_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__20_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__21_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__22_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__23_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__24_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__25_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__26_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__27_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__28_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__29_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__30_,
         dp_ex_stage_alu_shifter_rol_32_ML_int_1__31_,
         dp_ex_stage_alu_shifter_ror_30_n15,
         dp_ex_stage_alu_shifter_ror_30_n14,
         dp_ex_stage_alu_shifter_ror_30_n13,
         dp_ex_stage_alu_shifter_ror_30_n12,
         dp_ex_stage_alu_shifter_ror_30_n11,
         dp_ex_stage_alu_shifter_ror_30_n10, dp_ex_stage_alu_shifter_ror_30_n9,
         dp_ex_stage_alu_shifter_ror_30_n8, dp_ex_stage_alu_shifter_ror_30_n7,
         dp_ex_stage_alu_shifter_ror_30_n6, dp_ex_stage_alu_shifter_ror_30_n5,
         dp_ex_stage_alu_shifter_ror_30_n4, dp_ex_stage_alu_shifter_ror_30_n3,
         dp_ex_stage_alu_shifter_ror_30_n2, dp_ex_stage_alu_shifter_ror_30_n1,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__0_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__1_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__2_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__3_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__4_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__5_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__6_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__7_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__8_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__9_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__10_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__11_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__12_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__13_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__14_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__15_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__16_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__17_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__18_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__19_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__20_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__21_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__22_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__23_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__24_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__25_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__26_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__27_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__28_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__29_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__30_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_4__31_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__0_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__1_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__2_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__3_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__4_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__5_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__6_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__7_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__8_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__9_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__10_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__11_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__12_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__13_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__14_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__15_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__16_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__17_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__18_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__19_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__20_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__21_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__22_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__23_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__24_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__25_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__26_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__27_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__28_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__29_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__30_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_3__31_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__0_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__1_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__2_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__3_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__4_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__5_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__6_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__7_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__8_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__9_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__10_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__11_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__12_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__13_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__14_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__15_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__16_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__17_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__18_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__19_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__20_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__21_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__22_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__23_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__24_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__25_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__26_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__27_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__28_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__29_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__30_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_2__31_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__0_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__1_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__2_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__3_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__4_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__5_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__6_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__7_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__8_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__9_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__10_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__11_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__12_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__13_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__14_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__15_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__16_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__17_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__18_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__19_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__20_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__21_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__22_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__23_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__24_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__25_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__26_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__27_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__28_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__29_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__30_,
         dp_ex_stage_alu_shifter_ror_30_MR_int_1__31_,
         dp_ex_stage_alu_r61_n222, dp_ex_stage_alu_r61_n221,
         dp_ex_stage_alu_r61_n220, dp_ex_stage_alu_r61_n219,
         dp_ex_stage_alu_r61_n218, dp_ex_stage_alu_r61_n217,
         dp_ex_stage_alu_r61_n216, dp_ex_stage_alu_r61_n215,
         dp_ex_stage_alu_r61_n214, dp_ex_stage_alu_r61_n213,
         dp_ex_stage_alu_r61_n212, dp_ex_stage_alu_r61_n211,
         dp_ex_stage_alu_r61_n210, dp_ex_stage_alu_r61_n209,
         dp_ex_stage_alu_r61_n208, dp_ex_stage_alu_r61_n207,
         dp_ex_stage_alu_r61_n206, dp_ex_stage_alu_r61_n205,
         dp_ex_stage_alu_r61_n204, dp_ex_stage_alu_r61_n203,
         dp_ex_stage_alu_r61_n202, dp_ex_stage_alu_r61_n201,
         dp_ex_stage_alu_r61_n200, dp_ex_stage_alu_r61_n199,
         dp_ex_stage_alu_r61_n198, dp_ex_stage_alu_r61_n197,
         dp_ex_stage_alu_r61_n196, dp_ex_stage_alu_r61_n195,
         dp_ex_stage_alu_r61_n194, dp_ex_stage_alu_r61_n193,
         dp_ex_stage_alu_r61_n192, dp_ex_stage_alu_r61_n191,
         dp_ex_stage_alu_r61_n190, dp_ex_stage_alu_r61_n189,
         dp_ex_stage_alu_r61_n188, dp_ex_stage_alu_r61_n187,
         dp_ex_stage_alu_r61_n186, dp_ex_stage_alu_r61_n185,
         dp_ex_stage_alu_r61_n184, dp_ex_stage_alu_r61_n183,
         dp_ex_stage_alu_r61_n182, dp_ex_stage_alu_r61_n181,
         dp_ex_stage_alu_r61_n180, dp_ex_stage_alu_r61_n179,
         dp_ex_stage_alu_r61_n178, dp_ex_stage_alu_r61_n177,
         dp_ex_stage_alu_r61_n176, dp_ex_stage_alu_r61_n175,
         dp_ex_stage_alu_r61_n174, dp_ex_stage_alu_r61_n173,
         dp_ex_stage_alu_r61_n172, dp_ex_stage_alu_r61_n171,
         dp_ex_stage_alu_r61_n170, dp_ex_stage_alu_r61_n169,
         dp_ex_stage_alu_r61_n168, dp_ex_stage_alu_r61_n167,
         dp_ex_stage_alu_r61_n166, dp_ex_stage_alu_r61_n165,
         dp_ex_stage_alu_r61_n164, dp_ex_stage_alu_r61_n163,
         dp_ex_stage_alu_r61_n162, dp_ex_stage_alu_r61_n161,
         dp_ex_stage_alu_r61_n160, dp_ex_stage_alu_r61_n159,
         dp_ex_stage_alu_r61_n158, dp_ex_stage_alu_r61_n157,
         dp_ex_stage_alu_r61_n156, dp_ex_stage_alu_r61_n155,
         dp_ex_stage_alu_r61_n154, dp_ex_stage_alu_r61_n153,
         dp_ex_stage_alu_r61_n152, dp_ex_stage_alu_r61_n151,
         dp_ex_stage_alu_r61_n150, dp_ex_stage_alu_r61_n149,
         dp_ex_stage_alu_r61_n148, dp_ex_stage_alu_r61_n147,
         dp_ex_stage_alu_r61_n146, dp_ex_stage_alu_r61_n145,
         dp_ex_stage_alu_r61_n144, dp_ex_stage_alu_r61_n143,
         dp_ex_stage_alu_r61_n142, dp_ex_stage_alu_r61_n141,
         dp_ex_stage_alu_r61_n140, dp_ex_stage_alu_r61_n139,
         dp_ex_stage_alu_r61_n138, dp_ex_stage_alu_r61_n137,
         dp_ex_stage_alu_r61_n136, dp_ex_stage_alu_r61_n135,
         dp_ex_stage_alu_r61_n134, dp_ex_stage_alu_r61_n133,
         dp_ex_stage_alu_r61_n132, dp_ex_stage_alu_r61_n131,
         dp_ex_stage_alu_r61_n130, dp_ex_stage_alu_r61_n129,
         dp_ex_stage_alu_r61_n128, dp_ex_stage_alu_r61_n127,
         dp_ex_stage_alu_r61_n126, dp_ex_stage_alu_r61_n125,
         dp_ex_stage_alu_r61_n124, dp_ex_stage_alu_r61_n123,
         dp_ex_stage_alu_r61_n122, dp_ex_stage_alu_r61_n121,
         dp_ex_stage_alu_r61_n120, dp_ex_stage_alu_r61_n119,
         dp_ex_stage_alu_r61_n118, dp_ex_stage_alu_r61_n117,
         dp_ex_stage_alu_r61_n116, dp_ex_stage_alu_r61_n115,
         dp_ex_stage_alu_r61_n114, dp_ex_stage_alu_r61_n113,
         dp_ex_stage_alu_r61_n112, dp_ex_stage_alu_r61_n111,
         dp_ex_stage_alu_r61_n110, dp_ex_stage_alu_r61_n109,
         dp_ex_stage_alu_r61_n108, dp_ex_stage_alu_r61_n107,
         dp_ex_stage_alu_r61_n106, dp_ex_stage_alu_r61_n105,
         dp_ex_stage_alu_r61_n104, dp_ex_stage_alu_r61_n103,
         dp_ex_stage_alu_r61_n102, dp_ex_stage_alu_r61_n101,
         dp_ex_stage_alu_r61_n100, dp_ex_stage_alu_r61_n99,
         dp_ex_stage_alu_r61_n98, dp_ex_stage_alu_r61_n97,
         dp_ex_stage_alu_r61_n96, dp_ex_stage_alu_r61_n95,
         dp_ex_stage_alu_r61_n94, dp_ex_stage_alu_r61_n93,
         dp_ex_stage_alu_r61_n92, dp_ex_stage_alu_r61_n91,
         dp_ex_stage_alu_r61_n90, dp_ex_stage_alu_r61_n89,
         dp_ex_stage_alu_r61_n88, dp_ex_stage_alu_r61_n87,
         dp_ex_stage_alu_r61_n86, dp_ex_stage_alu_r61_n85,
         dp_ex_stage_alu_r61_n84, dp_ex_stage_alu_r61_n83,
         dp_ex_stage_alu_r61_n82, dp_ex_stage_alu_r61_n81,
         dp_ex_stage_alu_r61_n80, dp_ex_stage_alu_r61_n79,
         dp_ex_stage_alu_r61_n78, dp_ex_stage_alu_r61_n77,
         dp_ex_stage_alu_r61_n76, dp_ex_stage_alu_r61_n75,
         dp_ex_stage_alu_r61_n74, dp_ex_stage_alu_r61_n73,
         dp_ex_stage_alu_r61_n72, dp_ex_stage_alu_r61_n71,
         dp_ex_stage_alu_r61_n70, dp_ex_stage_alu_r61_n69,
         dp_ex_stage_alu_r61_n68, dp_ex_stage_alu_r61_n67,
         dp_ex_stage_alu_r61_n66, dp_ex_stage_alu_r61_n65,
         dp_ex_stage_alu_r61_n64, dp_ex_stage_alu_r61_n63,
         dp_ex_stage_alu_r61_n62, dp_ex_stage_alu_r61_n61,
         dp_ex_stage_alu_r61_n60, dp_ex_stage_alu_r61_n59,
         dp_ex_stage_alu_r61_n58, dp_ex_stage_alu_r61_n57,
         dp_ex_stage_alu_r61_n56, dp_ex_stage_alu_r61_n55,
         dp_ex_stage_alu_r61_n54, dp_ex_stage_alu_r61_n53,
         dp_ex_stage_alu_r61_n52, dp_ex_stage_alu_r61_n51,
         dp_ex_stage_alu_r61_n50, dp_ex_stage_alu_r61_n49,
         dp_ex_stage_alu_r61_n48, dp_ex_stage_alu_r61_n47,
         dp_ex_stage_alu_r61_n46, dp_ex_stage_alu_r61_n45,
         dp_ex_stage_alu_r61_n44, dp_ex_stage_alu_r61_n43,
         dp_ex_stage_alu_r61_n42, dp_ex_stage_alu_r61_n41,
         dp_ex_stage_alu_r61_n40, dp_ex_stage_alu_r61_n39,
         dp_ex_stage_alu_r61_n38, dp_ex_stage_alu_r61_n37,
         dp_ex_stage_alu_r61_n36, dp_ex_stage_alu_r61_n35,
         dp_ex_stage_alu_r61_n34, dp_ex_stage_alu_r61_n33,
         dp_ex_stage_alu_r61_n32, dp_ex_stage_alu_r61_n31,
         dp_ex_stage_alu_r61_n30, dp_ex_stage_alu_r61_n29,
         dp_ex_stage_alu_r61_n28, dp_ex_stage_alu_r61_n27,
         dp_ex_stage_alu_r61_n26, dp_ex_stage_alu_r61_n25,
         dp_ex_stage_alu_r61_n24, dp_ex_stage_alu_r61_n23,
         dp_ex_stage_alu_r61_n22, dp_ex_stage_alu_r61_n21,
         dp_ex_stage_alu_r61_n20, dp_ex_stage_alu_r61_n19,
         dp_ex_stage_alu_r61_n18, dp_ex_stage_alu_r61_n17,
         dp_ex_stage_alu_r61_n16, dp_ex_stage_alu_r61_n15,
         dp_ex_stage_alu_r61_n14, dp_ex_stage_alu_r61_n13,
         dp_ex_stage_alu_r61_n12, dp_ex_stage_alu_r61_n11,
         dp_ex_stage_alu_r61_n10, dp_ex_stage_alu_r61_n9,
         dp_ex_stage_alu_r61_n8, dp_ex_stage_alu_r61_n7,
         dp_ex_stage_alu_r61_n6, dp_ex_stage_alu_r61_n5,
         dp_ex_stage_alu_r61_n4, dp_ex_stage_alu_r61_n3,
         dp_ex_stage_alu_r61_n2, dp_ex_stage_alu_r61_n1,
         dp_ex_stage_alu_r60_n315, dp_ex_stage_alu_r60_n314,
         dp_ex_stage_alu_r60_n313, dp_ex_stage_alu_r60_n312,
         dp_ex_stage_alu_r60_n311, dp_ex_stage_alu_r60_n310,
         dp_ex_stage_alu_r60_n309, dp_ex_stage_alu_r60_n308,
         dp_ex_stage_alu_r60_n307, dp_ex_stage_alu_r60_n306,
         dp_ex_stage_alu_r60_n305, dp_ex_stage_alu_r60_n304,
         dp_ex_stage_alu_r60_n303, dp_ex_stage_alu_r60_n302,
         dp_ex_stage_alu_r60_n301, dp_ex_stage_alu_r60_n300,
         dp_ex_stage_alu_r60_n299, dp_ex_stage_alu_r60_n298,
         dp_ex_stage_alu_r60_n297, dp_ex_stage_alu_r60_n296,
         dp_ex_stage_alu_r60_n295, dp_ex_stage_alu_r60_n294,
         dp_ex_stage_alu_r60_n293, dp_ex_stage_alu_r60_n292,
         dp_ex_stage_alu_r60_n291, dp_ex_stage_alu_r60_n290,
         dp_ex_stage_alu_r60_n289, dp_ex_stage_alu_r60_n288,
         dp_ex_stage_alu_r60_n287, dp_ex_stage_alu_r60_n286,
         dp_ex_stage_alu_r60_n285, dp_ex_stage_alu_r60_n284,
         dp_ex_stage_alu_r60_n283, dp_ex_stage_alu_r60_n282,
         dp_ex_stage_alu_r60_n281, dp_ex_stage_alu_r60_n280,
         dp_ex_stage_alu_r60_n279, dp_ex_stage_alu_r60_n278,
         dp_ex_stage_alu_r60_n277, dp_ex_stage_alu_r60_n276,
         dp_ex_stage_alu_r60_n275, dp_ex_stage_alu_r60_n274,
         dp_ex_stage_alu_r60_n273, dp_ex_stage_alu_r60_n272,
         dp_ex_stage_alu_r60_n271, dp_ex_stage_alu_r60_n270,
         dp_ex_stage_alu_r60_n269, dp_ex_stage_alu_r60_n268,
         dp_ex_stage_alu_r60_n267, dp_ex_stage_alu_r60_n266,
         dp_ex_stage_alu_r60_n265, dp_ex_stage_alu_r60_n264,
         dp_ex_stage_alu_r60_n263, dp_ex_stage_alu_r60_n262,
         dp_ex_stage_alu_r60_n261, dp_ex_stage_alu_r60_n260,
         dp_ex_stage_alu_r60_n259, dp_ex_stage_alu_r60_n258,
         dp_ex_stage_alu_r60_n257, dp_ex_stage_alu_r60_n256,
         dp_ex_stage_alu_r60_n255, dp_ex_stage_alu_r60_n254,
         dp_ex_stage_alu_r60_n253, dp_ex_stage_alu_r60_n252,
         dp_ex_stage_alu_r60_n251, dp_ex_stage_alu_r60_n250,
         dp_ex_stage_alu_r60_n249, dp_ex_stage_alu_r60_n248,
         dp_ex_stage_alu_r60_n247, dp_ex_stage_alu_r60_n246,
         dp_ex_stage_alu_r60_n245, dp_ex_stage_alu_r60_n244,
         dp_ex_stage_alu_r60_n243, dp_ex_stage_alu_r60_n242,
         dp_ex_stage_alu_r60_n241, dp_ex_stage_alu_r60_n240,
         dp_ex_stage_alu_r60_n239, dp_ex_stage_alu_r60_n238,
         dp_ex_stage_alu_r60_n237, dp_ex_stage_alu_r60_n236,
         dp_ex_stage_alu_r60_n235, dp_ex_stage_alu_r60_n234,
         dp_ex_stage_alu_r60_n233, dp_ex_stage_alu_r60_n232,
         dp_ex_stage_alu_r60_n231, dp_ex_stage_alu_r60_n230,
         dp_ex_stage_alu_r60_n229, dp_ex_stage_alu_r60_n228,
         dp_ex_stage_alu_r60_n227, dp_ex_stage_alu_r60_n226,
         dp_ex_stage_alu_r60_n225, dp_ex_stage_alu_r60_n224,
         dp_ex_stage_alu_r60_n223, dp_ex_stage_alu_r60_n222,
         dp_ex_stage_alu_r60_n221, dp_ex_stage_alu_r60_n220,
         dp_ex_stage_alu_r60_n219, dp_ex_stage_alu_r60_n218,
         dp_ex_stage_alu_r60_n217, dp_ex_stage_alu_r60_n216,
         dp_ex_stage_alu_r60_n215, dp_ex_stage_alu_r60_n214,
         dp_ex_stage_alu_r60_n213, dp_ex_stage_alu_r60_n212,
         dp_ex_stage_alu_r60_n211, dp_ex_stage_alu_r60_n210,
         dp_ex_stage_alu_r60_n209, dp_ex_stage_alu_r60_n208,
         dp_ex_stage_alu_r60_n207, dp_ex_stage_alu_r60_n206,
         dp_ex_stage_alu_r60_n205, dp_ex_stage_alu_r60_n204,
         dp_ex_stage_alu_r60_n203, dp_ex_stage_alu_r60_n202,
         dp_ex_stage_alu_r60_n201, dp_ex_stage_alu_r60_n200,
         dp_ex_stage_alu_r60_n199, dp_ex_stage_alu_r60_n198,
         dp_ex_stage_alu_r60_n197, dp_ex_stage_alu_r60_n196,
         dp_ex_stage_alu_r60_n195, dp_ex_stage_alu_r60_n194,
         dp_ex_stage_alu_r60_n193, dp_ex_stage_alu_r60_n192,
         dp_ex_stage_alu_r60_n191, dp_ex_stage_alu_r60_n190,
         dp_ex_stage_alu_r60_n189, dp_ex_stage_alu_r60_n188,
         dp_ex_stage_alu_r60_n187, dp_ex_stage_alu_r60_n186,
         dp_ex_stage_alu_r60_n185, dp_ex_stage_alu_r60_n184,
         dp_ex_stage_alu_r60_n183, dp_ex_stage_alu_r60_n182,
         dp_ex_stage_alu_r60_n181, dp_ex_stage_alu_r60_n180,
         dp_ex_stage_alu_r60_n179, dp_ex_stage_alu_r60_n178,
         dp_ex_stage_alu_r60_n177, dp_ex_stage_alu_r60_n176,
         dp_ex_stage_alu_r60_n175, dp_ex_stage_alu_r60_n174,
         dp_ex_stage_alu_r60_n173, dp_ex_stage_alu_r60_n172,
         dp_ex_stage_alu_r60_n171, dp_ex_stage_alu_r60_n170,
         dp_ex_stage_alu_r60_n169, dp_ex_stage_alu_r60_n168,
         dp_ex_stage_alu_r60_n167, dp_ex_stage_alu_r60_n166,
         dp_ex_stage_alu_r60_n165, dp_ex_stage_alu_r60_n164,
         dp_ex_stage_alu_r60_n163, dp_ex_stage_alu_r60_n162,
         dp_ex_stage_alu_r60_n161, dp_ex_stage_alu_r60_n160,
         dp_ex_stage_alu_r60_n159, dp_ex_stage_alu_r60_n158,
         dp_ex_stage_alu_r60_n157, dp_ex_stage_alu_r60_n156,
         dp_ex_stage_alu_r60_n155, dp_ex_stage_alu_r60_n154,
         dp_ex_stage_alu_r60_n153, dp_ex_stage_alu_r60_n152,
         dp_ex_stage_alu_r60_n151, dp_ex_stage_alu_r60_n150,
         dp_ex_stage_alu_r60_n149, dp_ex_stage_alu_r60_n148,
         dp_ex_stage_alu_r60_n147, dp_ex_stage_alu_r60_n146,
         dp_ex_stage_alu_r60_n145, dp_ex_stage_alu_r60_n144,
         dp_ex_stage_alu_r60_n143, dp_ex_stage_alu_r60_n142,
         dp_ex_stage_alu_r60_n141, dp_ex_stage_alu_r60_n140,
         dp_ex_stage_alu_r60_n139, dp_ex_stage_alu_r60_n138,
         dp_ex_stage_alu_r60_n137, dp_ex_stage_alu_r60_n136,
         dp_ex_stage_alu_r60_n135, dp_ex_stage_alu_r60_n134,
         dp_ex_stage_alu_r60_n133, dp_ex_stage_alu_r60_n132,
         dp_ex_stage_alu_r60_n131, dp_ex_stage_alu_r60_n130,
         dp_ex_stage_alu_r60_n129, dp_ex_stage_alu_r60_n128,
         dp_ex_stage_alu_r60_n127, dp_ex_stage_alu_r60_n126,
         dp_ex_stage_alu_r60_n125, dp_ex_stage_alu_r60_n124,
         dp_ex_stage_alu_r60_n123, dp_ex_stage_alu_r60_n122,
         dp_ex_stage_alu_r60_n121, dp_ex_stage_alu_r60_n120,
         dp_ex_stage_alu_r60_n119, dp_ex_stage_alu_r60_n118,
         dp_ex_stage_alu_r60_n117, dp_ex_stage_alu_r60_n116,
         dp_ex_stage_alu_r60_n115, dp_ex_stage_alu_r60_n114,
         dp_ex_stage_alu_r60_n113, dp_ex_stage_alu_r60_n112,
         dp_ex_stage_alu_r60_n111, dp_ex_stage_alu_r60_n110,
         dp_ex_stage_alu_r60_n109, dp_ex_stage_alu_r60_n108,
         dp_ex_stage_alu_r60_n107, dp_ex_stage_alu_r60_n106,
         dp_ex_stage_alu_r60_n105, dp_ex_stage_alu_r60_n104,
         dp_ex_stage_alu_r60_n103, dp_ex_stage_alu_r60_n102,
         dp_ex_stage_alu_r60_n101, dp_ex_stage_alu_r60_n100,
         dp_ex_stage_alu_r60_n99, dp_ex_stage_alu_r60_n98,
         dp_ex_stage_alu_r60_n97, dp_ex_stage_alu_r60_n96,
         dp_ex_stage_alu_r60_n95, dp_ex_stage_alu_r60_n94,
         dp_ex_stage_alu_r60_n93, dp_ex_stage_alu_r60_n92,
         dp_ex_stage_alu_r60_n91, dp_ex_stage_alu_r60_n90,
         dp_ex_stage_alu_r60_n89, dp_ex_stage_alu_r60_n88,
         dp_ex_stage_alu_r60_n87, dp_ex_stage_alu_r60_n86,
         dp_ex_stage_alu_r60_n85, dp_ex_stage_alu_r60_n84,
         dp_ex_stage_alu_r60_n83, dp_ex_stage_alu_r60_n82,
         dp_ex_stage_alu_r60_n81, dp_ex_stage_alu_r60_n80,
         dp_ex_stage_alu_r60_n79, dp_ex_stage_alu_r60_n78,
         dp_ex_stage_alu_r60_n77, dp_ex_stage_alu_r60_n76,
         dp_ex_stage_alu_r60_n75, dp_ex_stage_alu_r60_n74,
         dp_ex_stage_alu_r60_n73, dp_ex_stage_alu_r60_n72,
         dp_ex_stage_alu_r60_n71, dp_ex_stage_alu_r60_n70,
         dp_ex_stage_alu_r60_n69, dp_ex_stage_alu_r60_n68,
         dp_ex_stage_alu_r60_n67, dp_ex_stage_alu_r60_n66,
         dp_ex_stage_alu_r60_n65, dp_ex_stage_alu_r60_n64,
         dp_ex_stage_alu_r60_n63, dp_ex_stage_alu_r60_n62,
         dp_ex_stage_alu_r60_n61, dp_ex_stage_alu_r60_n60,
         dp_ex_stage_alu_r60_n59, dp_ex_stage_alu_r60_n58,
         dp_ex_stage_alu_r60_n57, dp_ex_stage_alu_r60_n56,
         dp_ex_stage_alu_r60_n55, dp_ex_stage_alu_r60_n54,
         dp_ex_stage_alu_r60_n53, dp_ex_stage_alu_r60_n52,
         dp_ex_stage_alu_r60_n51, dp_ex_stage_alu_r60_n50,
         dp_ex_stage_alu_r60_n49, dp_ex_stage_alu_r60_n48,
         dp_ex_stage_alu_r60_n47, dp_ex_stage_alu_r60_n46,
         dp_ex_stage_alu_r60_n45, dp_ex_stage_alu_r60_n44,
         dp_ex_stage_alu_r60_n43, dp_ex_stage_alu_r60_n42,
         dp_ex_stage_alu_r60_n41, dp_ex_stage_alu_r60_n40,
         dp_ex_stage_alu_r60_n39, dp_ex_stage_alu_r60_n38,
         dp_ex_stage_alu_r60_n37, dp_ex_stage_alu_r60_n36,
         dp_ex_stage_alu_r60_n35, dp_ex_stage_alu_r60_n34,
         dp_ex_stage_alu_r60_n33, dp_ex_stage_alu_r60_n32,
         dp_ex_stage_alu_r60_n31, dp_ex_stage_alu_r60_n30,
         dp_ex_stage_alu_r60_n29, dp_ex_stage_alu_r60_n28,
         dp_ex_stage_alu_r60_n27, dp_ex_stage_alu_r60_n26,
         dp_ex_stage_alu_r60_n25, dp_ex_stage_alu_r60_n24,
         dp_ex_stage_alu_r60_n23, dp_ex_stage_alu_r60_n22,
         dp_ex_stage_alu_r60_n21, dp_ex_stage_alu_r60_n20,
         dp_ex_stage_alu_r60_n19, dp_ex_stage_alu_r60_n17,
         dp_ex_stage_alu_r60_n16, dp_ex_stage_alu_r60_n15,
         dp_ex_stage_alu_r60_n14, dp_ex_stage_alu_r60_n13,
         dp_ex_stage_alu_r60_n12, dp_ex_stage_alu_r60_n11,
         dp_ex_stage_alu_r60_n10, dp_ex_stage_alu_r60_n9,
         dp_ex_stage_alu_r60_n8, dp_ex_stage_alu_r60_n7,
         dp_ex_stage_alu_r60_n6, dp_ex_stage_alu_r60_n5,
         dp_ex_stage_alu_r60_n4, dp_ex_stage_alu_r60_n3,
         dp_ex_stage_alu_r60_n2, dp_ex_stage_alu_r60_n1;
  wire   [4:0] alu_op_i;
  wire   [5:4] CU_I_cw2;
  wire   [4:0] dp_rd_fwd_ex_o;
  wire   [31:0] dp_data_mem_ex_o;
  wire   [31:0] dp_alu_out_ex_o;
  wire   [31:0] dp_npc_ex_i;
  wire   [31:0] dp_imm_ex_i;
  wire   [31:0] dp_rf_out1_ex_i;
  wire   [4:0] dp_rd_fwd_id_o;
  wire   [31:0] dp_npc_id_o;
  wire   [31:0] dp_imm_id_o;
  wire   [31:0] dp_rf_out2_id_o;
  wire   [31:0] dp_rf_out1_id_o;
  wire   [31:0] dp_wr_data_id_i;
  wire   [4:0] dp_rd_fwd_wb_i;
  wire   [31:0] dp_npc_if_o;
  wire   [31:0] dp_id_stage_out2_i;
  wire   [31:0] dp_id_stage_out1_i;
  wire   [4:0] dp_id_stage_p_addr_wRD;
  wire   [4:0] dp_id_stage_p_addr_wRS2;
  wire   [4:0] dp_id_stage_p_addr_wRS1;
  wire   [3:0] dp_id_stage_regfile_ControlUnit_next_state;
  wire   [5:0] dp_id_stage_regfile_DataPath_mux_wr_out;
  wire   [5:0] dp_id_stage_regfile_DataPath_mux_rd_out;
  wire   [5:0] dp_id_stage_regfile_DataPath_addr_w_p;
  wire   [5:0] dp_id_stage_regfile_DataPath_addr_rd2_p;
  wire   [5:0] dp_id_stage_regfile_DataPath_addr_rd1_p;
  wire   [31:0] dp_ex_stage_muxB_out;
  wire   [31:0] dp_ex_stage_muxA_out;
  wire   [31:0] dp_ex_stage_alu_shifter_out;
  wire   [31:0] dp_ex_stage_alu_adder_out;
  wire   [7:0] dp_ex_stage_alu_adder_carries;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry
;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry
;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry
;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry
;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry
;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry
;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry
;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry
;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry
;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry
;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry
;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry
;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry
;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1;
  wire   [3:0] dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry
;
  wire  
         [1:3] dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry
;
  tri   [31:0] DRAM_DATA;
  tri   [31:0] dp_z_word;

  INV_X2 CU_I_U264 ( .A(IRAM_DATA[0]), .ZN(CU_I_n291) );
  NAND2_X1 CU_I_U263 ( .A1(alu_op_i[1]), .A2(CU_I_n63), .ZN(CU_I_n79) );
  NAND2_X1 CU_I_U262 ( .A1(alu_op_i[3]), .A2(CU_I_n63), .ZN(CU_I_n82) );
  NAND2_X1 CU_I_U261 ( .A1(CU_I_n293), .A2(CU_I_n66), .ZN(CU_I_n167) );
  NAND2_X1 CU_I_U260 ( .A1(alu_op_i[2]), .A2(CU_I_n63), .ZN(CU_I_n81) );
  OAI211_X1 CU_I_U259 ( .C1(CU_I_n69), .C2(CU_I_n35), .A(CU_I_n80), .B(
        CU_I_n81), .ZN(CU_I_n213) );
  NAND2_X1 CU_I_U258 ( .A1(CU_I_n180), .A2(CU_I_n132), .ZN(CU_I_n102) );
  AND2_X1 CU_I_U257 ( .A1(CU_I_n102), .A2(CU_I_n127), .ZN(CU_I_n206) );
  AOI21_X1 CU_I_U256 ( .B1(CU_I_n117), .B2(CU_I_n180), .A(CU_I_n75), .ZN(
        CU_I_n145) );
  INV_X1 CU_I_U255 ( .A(CU_I_n47), .ZN(CU_I_n261) );
  OAI22_X1 CU_I_U254 ( .A1(pipe_if_id_en_i), .A2(CU_I_n8), .B1(CU_I_n175), 
        .B2(CU_I_n67), .ZN(CU_I_n241) );
  OAI21_X1 CU_I_U253 ( .B1(CU_I_n51), .B2(CU_I_n36), .A(CU_I_n79), .ZN(
        CU_I_n212) );
  NOR3_X1 CU_I_U252 ( .A1(CU_I_n157), .A2(IRAM_DATA[30]), .A3(CU_I_n276), .ZN(
        CU_I_n152) );
  AND2_X1 CU_I_U251 ( .A1(CU_I_n202), .A2(CU_I_n276), .ZN(CU_I_n176) );
  NOR3_X1 CU_I_U250 ( .A1(CU_I_n276), .A2(CU_I_n157), .A3(CU_I_n274), .ZN(
        CU_I_n207) );
  NOR4_X1 CU_I_U249 ( .A1(IRAM_DATA[30]), .A2(IRAM_DATA[29]), .A3(CU_I_n276), 
        .A4(CU_I_n279), .ZN(CU_I_n150) );
  AOI21_X1 CU_I_U248 ( .B1(CU_I_n278), .B2(CU_I_n276), .A(IRAM_DATA[30]), .ZN(
        CU_I_n162) );
  NAND4_X1 CU_I_U247 ( .A1(CU_I_n161), .A2(CU_I_n154), .A3(IRAM_DATA[29]), 
        .A4(CU_I_n276), .ZN(CU_I_n187) );
  AOI22_X1 CU_I_U246 ( .A1(CU_I_n259), .A2(CU_I_n276), .B1(IRAM_DATA[30]), 
        .B2(CU_I_n156), .ZN(CU_I_n147) );
  NOR3_X1 CU_I_U245 ( .A1(IRAM_DATA[28]), .A2(IRAM_DATA[30]), .A3(CU_I_n157), 
        .ZN(CU_I_n133) );
  NAND2_X1 CU_I_U244 ( .A1(CU_I_n154), .A2(CU_I_n133), .ZN(CU_I_n101) );
  NAND2_X1 CU_I_U243 ( .A1(CU_I_n38), .A2(CU_I_n117), .ZN(CU_I_n155) );
  AOI21_X1 CU_I_U242 ( .B1(CU_I_n132), .B2(CU_I_n38), .A(CU_I_n264), .ZN(
        CU_I_n131) );
  NOR2_X1 CU_I_U241 ( .A1(CU_I_n267), .A2(CU_I_n194), .ZN(CU_I_n192) );
  OAI211_X1 CU_I_U240 ( .C1(CU_I_n48), .C2(CU_I_n281), .A(CU_I_n130), .B(
        CU_I_n206), .ZN(CU_I_n111) );
  AOI211_X1 CU_I_U239 ( .C1(CU_I_n152), .C2(CU_I_n160), .A(CU_I_n111), .B(
        CU_I_n204), .ZN(CU_I_n87) );
  NOR3_X1 CU_I_U238 ( .A1(CU_I_n110), .A2(CU_I_n41), .A3(CU_I_n112), .ZN(
        CU_I_n109) );
  NAND2_X1 CU_I_U237 ( .A1(CU_I_n292), .A2(CU_I_n64), .ZN(CU_I_n166) );
  OAI211_X1 CU_I_U236 ( .C1(CU_I_n69), .C2(CU_I_n33), .A(CU_I_n80), .B(
        CU_I_n83), .ZN(CU_I_n215) );
  AOI22_X1 CU_I_U235 ( .A1(CU_I_n68), .A2(CU_I_cw1_1_), .B1(CU_I_n171), .B2(
        CU_I_n172), .ZN(CU_I_n170) );
  INV_X1 CU_I_U234 ( .A(CU_I_n170), .ZN(CU_I_n74) );
  AOI22_X1 CU_I_U233 ( .A1(CU_I_n291), .A2(IRAM_DATA[2]), .B1(CU_I_n289), .B2(
        CU_I_n94), .ZN(CU_I_n93) );
  OR2_X1 CU_I_U232 ( .A1(CU_I_n93), .A2(IRAM_DATA[3]), .ZN(CU_I_n88) );
  NAND2_X1 CU_I_U223 ( .A1(pipe_clear_n_i), .A2(CU_I_n30), .ZN(jump_en_i) );
  INV_X1 CU_I_U215 ( .A(IRAM_DATA[26]), .ZN(CU_I_n282) );
  INV_X1 CU_I_U214 ( .A(IRAM_DATA[4]), .ZN(CU_I_n286) );
  NAND2_X1 CU_I_U213 ( .A1(IRAM_READY), .A2(IRAM_ISSUE), .ZN(CU_I_n78) );
  INV_X1 CU_I_U212 ( .A(IRAM_DATA[27]), .ZN(CU_I_n279) );
  INV_X1 CU_I_U211 ( .A(IRAM_DATA[31]), .ZN(CU_I_n266) );
  INV_X1 CU_I_U210 ( .A(CU_I_n126), .ZN(CU_I_n285) );
  INV_X1 CU_I_U209 ( .A(CU_I_n185), .ZN(CU_I_n260) );
  NAND2_X1 CU_I_U208 ( .A1(regrd_sel_i), .A2(CU_I_n65), .ZN(CU_I_n190) );
  OAI21_X1 CU_I_U207 ( .B1(CU_I_n260), .B2(CU_I_n49), .A(CU_I_n190), .ZN(
        CU_I_n247) );
  AND3_X1 CU_I_U206 ( .A1(CU_I_n114), .A2(CU_I_n196), .A3(CU_I_n187), .ZN(
        CU_I_n197) );
  NAND2_X1 CU_I_U205 ( .A1(rf_rs2_en_i), .A2(CU_I_n66), .ZN(CU_I_n198) );
  OAI21_X1 CU_I_U204 ( .B1(CU_I_n197), .B2(CU_I_n49), .A(CU_I_n198), .ZN(
        CU_I_n251) );
  NAND2_X1 CU_I_U203 ( .A1(imm_isoff_i), .A2(CU_I_n66), .ZN(CU_I_n195) );
  OAI21_X1 CU_I_U202 ( .B1(CU_I_n268), .B2(CU_I_n49), .A(CU_I_n195), .ZN(
        CU_I_n250) );
  NAND2_X1 CU_I_U201 ( .A1(imm_uns_i), .A2(CU_I_n66), .ZN(CU_I_n193) );
  OAI21_X1 CU_I_U200 ( .B1(CU_I_n192), .B2(CU_I_n49), .A(CU_I_n193), .ZN(
        CU_I_n249) );
  NOR4_X1 CU_I_U199 ( .A1(CU_I_n267), .A2(CU_I_n179), .A3(CU_I_n184), .A4(
        CU_I_n181), .ZN(CU_I_n199) );
  NAND2_X1 CU_I_U198 ( .A1(rf_rs1_en_i), .A2(CU_I_n67), .ZN(CU_I_n200) );
  OAI21_X1 CU_I_U197 ( .B1(CU_I_n199), .B2(CU_I_n49), .A(CU_I_n200), .ZN(
        CU_I_n252) );
  OR3_X1 CU_I_U196 ( .A1(CU_I_n157), .A2(IRAM_DATA[28]), .A3(CU_I_n274), .ZN(
        CU_I_n116) );
  OAI21_X1 CU_I_U195 ( .B1(CU_I_n2), .B2(pipe_ex_mem_en_i), .A(CU_I_n182), 
        .ZN(CU_I_n248) );
  NAND2_X1 CU_I_U194 ( .A1(CU_I_n91), .A2(CU_I_n92), .ZN(CU_I_n90) );
  OAI21_X1 CU_I_U193 ( .B1(pipe_if_id_en_i), .B2(CU_I_n6), .A(CU_I_n182), .ZN(
        CU_I_n243) );
  NAND4_X1 CU_I_U192 ( .A1(CU_I_n91), .A2(IRAM_DATA[1]), .A3(IRAM_DATA[0]), 
        .A4(CU_I_n289), .ZN(CU_I_n128) );
  NAND2_X1 CU_I_U191 ( .A1(CU_I_n127), .A2(CU_I_n128), .ZN(CU_I_n105) );
  INV_X1 CU_I_U190 ( .A(IRAM_DATA[5]), .ZN(CU_I_n284) );
  NOR2_X1 CU_I_U189 ( .A1(IRAM_DATA[2]), .A2(CU_I_n291), .ZN(CU_I_n144) );
  NAND2_X1 CU_I_U188 ( .A1(DRAM_READNOTWRITE), .A2(CU_I_n67), .ZN(CU_I_n209)
         );
  OAI211_X1 CU_I_U187 ( .C1(CU_I_n69), .C2(CU_I_n16), .A(CU_I_n80), .B(
        CU_I_n209), .ZN(CU_I_n253) );
  OAI21_X1 CU_I_U186 ( .B1(CU_I_n51), .B2(CU_I_n3), .A(CU_I_n166), .ZN(
        CU_I_n226) );
  NAND2_X1 CU_I_U185 ( .A1(mem_in_en_i), .A2(CU_I_n65), .ZN(CU_I_n168) );
  OAI21_X1 CU_I_U184 ( .B1(CU_I_n51), .B2(CU_I_n5), .A(CU_I_n168), .ZN(
        CU_I_n228) );
  NAND2_X1 CU_I_U183 ( .A1(npc_wb_en_i), .A2(CU_I_n65), .ZN(CU_I_n169) );
  OAI21_X1 CU_I_U182 ( .B1(CU_I_n51), .B2(CU_I_n6), .A(CU_I_n169), .ZN(
        CU_I_n229) );
  NAND2_X1 CU_I_U181 ( .A1(wb_mux_sel_i), .A2(CU_I_n64), .ZN(CU_I_n165) );
  OAI21_X1 CU_I_U180 ( .B1(CU_I_n51), .B2(CU_I_n31), .A(CU_I_n165), .ZN(
        CU_I_n222) );
  NAND2_X1 CU_I_U179 ( .A1(rf_we_i), .A2(CU_I_n64), .ZN(CU_I_n164) );
  OAI21_X1 CU_I_U178 ( .B1(CU_I_n51), .B2(CU_I_n32), .A(CU_I_n164), .ZN(
        CU_I_n221) );
  OAI21_X1 CU_I_U177 ( .B1(CU_I_n51), .B2(CU_I_n34), .A(CU_I_n82), .ZN(
        CU_I_n214) );
  NAND2_X1 CU_I_U176 ( .A1(CU_I_n294), .A2(CU_I_n65), .ZN(CU_I_n77) );
  OAI21_X1 CU_I_U175 ( .B1(CU_I_n51), .B2(CU_I_n37), .A(CU_I_n77), .ZN(
        CU_I_n211) );
  OAI21_X1 CU_I_U174 ( .B1(CU_I_n51), .B2(CU_I_n4), .A(CU_I_n167), .ZN(
        CU_I_n227) );
  OAI22_X1 CU_I_U173 ( .A1(IRAM_DATA[0]), .A2(CU_I_n290), .B1(CU_I_n291), .B2(
        CU_I_n119), .ZN(CU_I_n135) );
  NAND4_X1 CU_I_U172 ( .A1(CU_I_n107), .A2(IRAM_DATA[5]), .A3(CU_I_n135), .A4(
        CU_I_n288), .ZN(CU_I_n129) );
  NAND4_X1 CU_I_U171 ( .A1(CU_I_n107), .A2(IRAM_DATA[5]), .A3(IRAM_DATA[0]), 
        .A4(CU_I_n108), .ZN(CU_I_n103) );
  INV_X1 CU_I_U170 ( .A(IRAM_DATA[1]), .ZN(CU_I_n290) );
  NAND2_X1 CU_I_U169 ( .A1(IRAM_DATA[2]), .A2(IRAM_DATA[1]), .ZN(CU_I_n108) );
  NAND2_X1 CU_I_U168 ( .A1(CU_I_n25), .A2(CU_I_n64), .ZN(CU_I_n83) );
  NOR2_X1 CU_I_U167 ( .A1(IRAM_DATA[28]), .A2(IRAM_DATA[29]), .ZN(CU_I_n201)
         );
  AOI21_X1 CU_I_U166 ( .B1(IRAM_DATA[29]), .B2(CU_I_n281), .A(CU_I_n274), .ZN(
        CU_I_n163) );
  INV_X1 CU_I_U165 ( .A(IRAM_DATA[2]), .ZN(CU_I_n289) );
  NOR4_X1 CU_I_U164 ( .A1(CU_I_n96), .A2(CU_I_n97), .A3(CU_I_n98), .A4(
        CU_I_n99), .ZN(CU_I_n95) );
  OAI22_X1 CU_I_U163 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n36), .B1(CU_I_n95), 
        .B2(CU_I_n49), .ZN(CU_I_n217) );
  INV_X1 CU_I_U162 ( .A(CU_I_n187), .ZN(CU_I_n257) );
  OAI22_X1 CU_I_U161 ( .A1(pipe_if_id_en_i), .A2(CU_I_n4), .B1(CU_I_n183), 
        .B2(CU_I_n49), .ZN(CU_I_n245) );
  OAI22_X1 CU_I_U160 ( .A1(pipe_if_id_en_i), .A2(CU_I_n23), .B1(CU_I_n50), 
        .B2(CU_I_n13), .ZN(CU_I_n236) );
  OAI211_X1 CU_I_U159 ( .C1(CU_I_n271), .C2(CU_I_n88), .A(CU_I_n89), .B(
        CU_I_n90), .ZN(CU_I_n86) );
  AOI211_X1 CU_I_U158 ( .C1(CU_I_n85), .C2(CU_I_n291), .A(CU_I_n86), .B(
        CU_I_n261), .ZN(CU_I_n84) );
  OAI22_X1 CU_I_U157 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n37), .B1(CU_I_n84), 
        .B2(CU_I_n49), .ZN(CU_I_n216) );
  OAI22_X1 CU_I_U156 ( .A1(pipe_if_id_en_i), .A2(CU_I_n11), .B1(CU_I_n268), 
        .B2(CU_I_n49), .ZN(CU_I_n238) );
  OAI22_X1 CU_I_U155 ( .A1(pipe_if_id_en_i), .A2(CU_I_n12), .B1(CU_I_n26), 
        .B2(CU_I_n49), .ZN(CU_I_n237) );
  INV_X1 CU_I_U154 ( .A(CU_I_n181), .ZN(CU_I_n258) );
  OAI22_X1 CU_I_U153 ( .A1(pipe_if_id_en_i), .A2(CU_I_n7), .B1(CU_I_n258), 
        .B2(CU_I_n49), .ZN(CU_I_n242) );
  NOR4_X1 CU_I_U152 ( .A1(CU_I_n263), .A2(CU_I_n149), .A3(CU_I_n150), .A4(
        CU_I_n265), .ZN(CU_I_n148) );
  OAI21_X1 CU_I_U151 ( .B1(CU_I_n162), .B2(CU_I_n163), .A(IRAM_DATA[31]), .ZN(
        CU_I_n146) );
  NAND4_X1 CU_I_U150 ( .A1(CU_I_n145), .A2(CU_I_n146), .A3(CU_I_n147), .A4(
        CU_I_n148), .ZN(CU_I_n112) );
  OAI22_X1 CU_I_U149 ( .A1(pipe_if_id_en_i), .A2(CU_I_n27), .B1(CU_I_n50), 
        .B2(CU_I_n15), .ZN(CU_I_n254) );
  OAI22_X1 CU_I_U148 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n22), .B1(CU_I_n50), 
        .B2(CU_I_n12), .ZN(CU_I_n235) );
  OAI22_X1 CU_I_U147 ( .A1(pipe_if_id_en_i), .A2(CU_I_n21), .B1(CU_I_n50), 
        .B2(CU_I_n11), .ZN(CU_I_n234) );
  OAI22_X1 CU_I_U146 ( .A1(pipe_if_id_en_i), .A2(CU_I_n19), .B1(CU_I_n50), 
        .B2(CU_I_n10), .ZN(CU_I_n233) );
  OAI22_X1 CU_I_U145 ( .A1(pipe_if_id_en_i), .A2(CU_I_n17), .B1(CU_I_n50), 
        .B2(CU_I_n9), .ZN(CU_I_n232) );
  OAI22_X1 CU_I_U144 ( .A1(pipe_if_id_en_i), .A2(CU_I_n15), .B1(CU_I_n50), 
        .B2(CU_I_n7), .ZN(CU_I_n230) );
  OAI22_X1 CU_I_U143 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n30), .B1(CU_I_n50), 
        .B2(CU_I_n21), .ZN(CU_I_n225) );
  OAI22_X1 CU_I_U142 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n31), .B1(CU_I_n50), 
        .B2(CU_I_n22), .ZN(CU_I_n224) );
  OAI22_X1 CU_I_U141 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n32), .B1(CU_I_n50), 
        .B2(CU_I_n23), .ZN(CU_I_n223) );
  INV_X1 CU_I_U140 ( .A(CU_I_n99), .ZN(CU_I_n262) );
  OAI211_X1 CU_I_U139 ( .C1(CU_I_n113), .C2(CU_I_n114), .A(CU_I_n115), .B(
        CU_I_n262), .ZN(CU_I_n110) );
  OAI22_X1 CU_I_U138 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n35), .B1(CU_I_n109), 
        .B2(CU_I_n68), .ZN(CU_I_n218) );
  OAI21_X1 CU_I_U137 ( .B1(CU_I_n139), .B2(CU_I_n114), .A(CU_I_n140), .ZN(
        CU_I_n138) );
  OAI211_X1 CU_I_U136 ( .C1(CU_I_n278), .C2(CU_I_n116), .A(CU_I_n101), .B(
        CU_I_n269), .ZN(CU_I_n137) );
  NOR3_X1 CU_I_U135 ( .A1(CU_I_n137), .A2(CU_I_n112), .A3(CU_I_n138), .ZN(
        CU_I_n136) );
  OAI22_X1 CU_I_U134 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n33), .B1(CU_I_n136), 
        .B2(CU_I_n67), .ZN(CU_I_n220) );
  NOR3_X1 CU_I_U133 ( .A1(CU_I_n124), .A2(CU_I_n105), .A3(CU_I_n125), .ZN(
        CU_I_n123) );
  OAI22_X1 CU_I_U132 ( .A1(pipe_ex_mem_en_i), .A2(CU_I_n34), .B1(CU_I_n123), 
        .B2(CU_I_n49), .ZN(CU_I_n219) );
  AOI22_X1 CU_I_U131 ( .A1(CU_I_n69), .A2(CU_I_cw3_4_), .B1(CU_I_n172), .B2(
        CU_I_cw2[4]), .ZN(CU_I_n210) );
  INV_X1 CU_I_U130 ( .A(CU_I_n210), .ZN(CU_I_n72) );
  AOI22_X1 CU_I_U129 ( .A1(CU_I_n68), .A2(CU_I_cw3_5_), .B1(CU_I_n172), .B2(
        CU_I_cw2[5]), .ZN(CU_I_n208) );
  INV_X1 CU_I_U128 ( .A(CU_I_n208), .ZN(CU_I_n73) );
  NOR2_X1 CU_I_U127 ( .A1(CU_I_n266), .A2(IRAM_DATA[30]), .ZN(CU_I_n161) );
  OAI22_X1 CU_I_U126 ( .A1(pipe_if_id_en_i), .A2(CU_I_n9), .B1(CU_I_n50), .B2(
        CU_I_n174), .ZN(CU_I_n240) );
  OAI22_X1 CU_I_U125 ( .A1(pipe_if_id_en_i), .A2(CU_I_n10), .B1(CU_I_n50), 
        .B2(CU_I_n173), .ZN(CU_I_n239) );
  OAI22_X1 CU_I_U124 ( .A1(pipe_if_id_en_i), .A2(CU_I_n5), .B1(CU_I_n50), .B2(
        CU_I_n178), .ZN(CU_I_n244) );
  INV_X1 CU_I_U123 ( .A(CU_I_n145), .ZN(CU_I_n70) );
  INV_X1 CU_I_U122 ( .A(CU_I_n189), .ZN(CU_I_n273) );
  NOR2_X1 CU_I_U121 ( .A1(CU_I_n273), .A2(CU_I_n184), .ZN(CU_I_n188) );
  NOR2_X1 CU_I_U120 ( .A1(CU_I_n114), .A2(IRAM_DATA[4]), .ZN(CU_I_n107) );
  NOR3_X1 CU_I_U119 ( .A1(IRAM_DATA[30]), .A2(IRAM_DATA[31]), .A3(
        IRAM_DATA[29]), .ZN(CU_I_n202) );
  NOR3_X1 CU_I_U118 ( .A1(CU_I_n274), .A2(IRAM_DATA[31]), .A3(CU_I_n275), .ZN(
        CU_I_n153) );
  OAI22_X1 CU_I_U117 ( .A1(IRAM_DATA[3]), .A2(CU_I_n291), .B1(CU_I_n144), .B2(
        CU_I_n283), .ZN(CU_I_n142) );
  AOI21_X1 CU_I_U116 ( .B1(CU_I_n106), .B2(CU_I_n119), .A(CU_I_n286), .ZN(
        CU_I_n143) );
  OAI211_X1 CU_I_U115 ( .C1(IRAM_DATA[1]), .C2(CU_I_n288), .A(CU_I_n291), .B(
        IRAM_DATA[2]), .ZN(CU_I_n141) );
  AOI221_X1 CU_I_U114 ( .B1(CU_I_n141), .B2(CU_I_n284), .C1(IRAM_DATA[1]), 
        .C2(CU_I_n142), .A(CU_I_n143), .ZN(CU_I_n139) );
  AOI211_X1 CU_I_U113 ( .C1(CU_I_n122), .C2(CU_I_n291), .A(IRAM_DATA[4]), .B(
        CU_I_n94), .ZN(CU_I_n121) );
  AOI21_X1 CU_I_U112 ( .B1(CU_I_n291), .B2(CU_I_n288), .A(CU_I_n108), .ZN(
        CU_I_n120) );
  OAI222_X1 CU_I_U111 ( .A1(CU_I_n288), .A2(CU_I_n119), .B1(IRAM_DATA[5]), 
        .B2(CU_I_n120), .C1(CU_I_n121), .C2(CU_I_n289), .ZN(CU_I_n118) );
  AOI221_X1 CU_I_U110 ( .B1(CU_I_n106), .B2(IRAM_DATA[1]), .C1(IRAM_DATA[4]), 
        .C2(CU_I_n288), .A(CU_I_n118), .ZN(CU_I_n113) );
  NOR2_X1 CU_I_U109 ( .A1(IRAM_DATA[27]), .A2(IRAM_DATA[26]), .ZN(CU_I_n160)
         );
  NOR3_X1 CU_I_U108 ( .A1(CU_I_n271), .A2(IRAM_DATA[5]), .A3(CU_I_n108), .ZN(
        CU_I_n85) );
  NOR2_X1 CU_I_U107 ( .A1(CU_I_n279), .A2(IRAM_DATA[26]), .ZN(CU_I_n132) );
  NOR2_X1 CU_I_U106 ( .A1(CU_I_n282), .A2(IRAM_DATA[27]), .ZN(CU_I_n117) );
  INV_X1 CU_I_U105 ( .A(is_zero_i), .ZN(CU_I_n76) );
  AOI22_X1 CU_I_U104 ( .A1(is_zero_i), .A2(CU_I_cw3_4_), .B1(CU_I_n76), .B2(
        CU_I_cw3_5_), .ZN(pipe_clear_n_i) );
  BUF_X1 CU_I_U103 ( .A(CU_I_n256), .Z(CU_I_n57) );
  BUF_X1 CU_I_U102 ( .A(CU_I_n256), .Z(CU_I_n56) );
  BUF_X1 CU_I_U101 ( .A(CU_I_n78), .Z(CU_I_n60) );
  AOI22_X1 CU_I_U100 ( .A1(CU_I_n157), .A2(CU_I_n117), .B1(CU_I_n160), .B2(
        CU_I_n161), .ZN(CU_I_n159) );
  INV_X1 CU_I_U99 ( .A(CU_I_n159), .ZN(CU_I_n259) );
  INV_X1 CU_I_U98 ( .A(CU_I_n201), .ZN(CU_I_n275) );
  INV_X1 CU_I_U97 ( .A(CU_I_n85), .ZN(CU_I_n270) );
  OAI21_X1 CU_I_U96 ( .B1(CU_I_n152), .B2(CU_I_n153), .A(CU_I_n154), .ZN(
        CU_I_n151) );
  INV_X1 CU_I_U95 ( .A(CU_I_n151), .ZN(CU_I_n265) );
  INV_X1 CU_I_U94 ( .A(CU_I_n107), .ZN(CU_I_n271) );
  INV_X1 CU_I_U93 ( .A(DRAM_ISSUE), .ZN(IRAM_ISSUE) );
  INV_X1 CU_I_U92 ( .A(CU_I_n132), .ZN(CU_I_n278) );
  NAND2_X1 CU_I_U91 ( .A1(CU_I_n176), .A2(CU_I_n132), .ZN(CU_I_n189) );
  INV_X1 CU_I_U90 ( .A(CU_I_n160), .ZN(CU_I_n281) );
  NOR2_X1 CU_I_U89 ( .A1(CU_I_n281), .A2(CU_I_n116), .ZN(CU_I_n149) );
  NAND2_X1 CU_I_U88 ( .A1(CU_I_n153), .A2(CU_I_n132), .ZN(CU_I_n196) );
  NAND2_X1 CU_I_U87 ( .A1(CU_I_n160), .A2(CU_I_n207), .ZN(CU_I_n115) );
  NAND2_X1 CU_I_U86 ( .A1(CU_I_n290), .A2(CU_I_n289), .ZN(CU_I_n119) );
  INV_X1 CU_I_U85 ( .A(CU_I_n106), .ZN(CU_I_n287) );
  AOI21_X1 CU_I_U84 ( .B1(CU_I_n85), .B2(CU_I_n287), .A(CU_I_n105), .ZN(
        CU_I_n104) );
  INV_X1 CU_I_U83 ( .A(pipe_clear_n_i), .ZN(CU_I_n75) );
  NAND2_X1 CU_I_U82 ( .A1(CU_I_n178), .A2(CU_I_n187), .ZN(CU_I_n181) );
  NAND2_X1 CU_I_U81 ( .A1(CU_I_n132), .A2(CU_I_n152), .ZN(CU_I_n134) );
  NAND2_X1 CU_I_U80 ( .A1(CU_I_n174), .A2(CU_I_n173), .ZN(CU_I_n184) );
  NAND2_X1 CU_I_U79 ( .A1(CU_I_n207), .A2(CU_I_n117), .ZN(CU_I_n89) );
  INV_X1 CU_I_U78 ( .A(CU_I_n134), .ZN(CU_I_n264) );
  NOR2_X1 CU_I_U77 ( .A1(CU_I_n288), .A2(CU_I_n284), .ZN(CU_I_n122) );
  NAND2_X1 CU_I_U76 ( .A1(CU_I_n152), .A2(CU_I_n117), .ZN(CU_I_n100) );
  INV_X1 CU_I_U75 ( .A(CU_I_n117), .ZN(CU_I_n280) );
  NOR2_X1 CU_I_U74 ( .A1(CU_I_n116), .A2(CU_I_n280), .ZN(CU_I_n99) );
  NAND2_X1 CU_I_U73 ( .A1(CU_I_n176), .A2(CU_I_n160), .ZN(CU_I_n114) );
  NOR2_X1 CU_I_U72 ( .A1(CU_I_n288), .A2(CU_I_n291), .ZN(CU_I_n106) );
  NOR3_X1 CU_I_U71 ( .A1(CU_I_n290), .A2(CU_I_n291), .A3(CU_I_n284), .ZN(
        CU_I_n94) );
  BUF_X1 CU_I_U70 ( .A(CU_I_n56), .Z(CU_I_n55) );
  BUF_X1 CU_I_U69 ( .A(CU_I_n57), .Z(CU_I_n52) );
  BUF_X1 CU_I_U68 ( .A(CU_I_n56), .Z(CU_I_n54) );
  BUF_X1 CU_I_U67 ( .A(CU_I_n57), .Z(CU_I_n53) );
  INV_X1 CU_I_U66 ( .A(CU_I_n155), .ZN(CU_I_n263) );
  INV_X1 CU_I_U65 ( .A(CU_I_n122), .ZN(CU_I_n283) );
  BUF_X1 CU_I_U64 ( .A(CU_I_n58), .Z(CU_I_n63) );
  INV_X1 CU_I_U63 ( .A(CU_I_n196), .ZN(CU_I_n267) );
  NAND2_X1 CU_I_U62 ( .A1(CU_I_n176), .A2(CU_I_n154), .ZN(CU_I_n177) );
  BUF_X1 CU_I_U61 ( .A(CU_I_n59), .Z(CU_I_n67) );
  BUF_X1 CU_I_U60 ( .A(CU_I_n59), .Z(CU_I_n64) );
  BUF_X1 CU_I_U59 ( .A(CU_I_n59), .Z(CU_I_n66) );
  INV_X1 CU_I_U58 ( .A(CU_I_n154), .ZN(CU_I_n277) );
  BUF_X1 CU_I_U57 ( .A(CU_I_n58), .Z(CU_I_n68) );
  BUF_X1 CU_I_U56 ( .A(CU_I_n58), .Z(CU_I_n65) );
  NAND2_X1 CU_I_U55 ( .A1(CU_I_n191), .A2(CU_I_n114), .ZN(CU_I_n179) );
  NAND2_X1 CU_I_U54 ( .A1(CU_I_n191), .A2(CU_I_n178), .ZN(CU_I_n185) );
  NAND2_X1 CU_I_U53 ( .A1(pipe_if_id_en_i), .A2(CU_I_n75), .ZN(CU_I_n80) );
  NOR2_X1 CU_I_U52 ( .A1(CU_I_n48), .A2(CU_I_n277), .ZN(CU_I_n98) );
  NOR2_X1 CU_I_U51 ( .A1(CU_I_n283), .A2(CU_I_n114), .ZN(CU_I_n91) );
  NOR2_X1 CU_I_U50 ( .A1(CU_I_n68), .A2(CU_I_n75), .ZN(CU_I_n172) );
  INV_X1 CU_I_U49 ( .A(CU_I_n91), .ZN(CU_I_n272) );
  INV_X1 CU_I_U48 ( .A(CU_I_n98), .ZN(CU_I_n269) );
  INV_X1 CU_I_U47 ( .A(CU_I_n186), .ZN(CU_I_n268) );
  INV_X1 CU_I_U46 ( .A(CU_I_n172), .ZN(CU_I_n71) );
  OR2_X1 CU_I_U45 ( .A1(CU_I_n177), .A2(CU_I_n51), .ZN(CU_I_n182) );
  BUF_X1 CU_I_U44 ( .A(CU_I_n71), .Z(CU_I_n49) );
  BUF_X1 CU_I_U43 ( .A(CU_I_n71), .Z(CU_I_n50) );
  BUF_X1 CU_I_U42 ( .A(CU_I_n71), .Z(CU_I_n51) );
  CLKBUF_X1 CU_I_U41 ( .A(CU_I_n78), .Z(CU_I_n59) );
  BUF_X2 CU_I_U40 ( .A(CU_I_n60), .Z(CU_I_n69) );
  INV_X2 CU_I_U39 ( .A(CU_I_n58), .ZN(pipe_if_id_en_i) );
  INV_X2 CU_I_U38 ( .A(IRAM_DATA[28]), .ZN(CU_I_n276) );
  OR4_X1 CU_I_U37 ( .A1(CU_I_n274), .A2(CU_I_n276), .A3(IRAM_DATA[29]), .A4(
        IRAM_DATA[31]), .ZN(CU_I_n48) );
  AOI211_X1 CU_I_U36 ( .C1(CU_I_n152), .C2(CU_I_n160), .A(CU_I_n41), .B(
        CU_I_n204), .ZN(CU_I_n47) );
  INV_X1 CU_I_U35 ( .A(IRAM_DATA[30]), .ZN(CU_I_n274) );
  AND3_X1 CU_I_U34 ( .A1(IRAM_DATA[30]), .A2(IRAM_DATA[29]), .A3(IRAM_DATA[31]), .ZN(CU_I_n205) );
  NOR2_X1 CU_I_U33 ( .A1(CU_I_n171), .A2(CU_I_n1), .ZN(CU_I_n175) );
  INV_X1 CU_I_U32 ( .A(CU_I_n43), .ZN(muxA_sel_i) );
  NOR2_X1 CU_I_U31 ( .A1(IRAM_DATA[29]), .A2(IRAM_DATA[31]), .ZN(CU_I_n42) );
  CLKBUF_X1 CU_I_U30 ( .A(CU_I_n111), .Z(CU_I_n41) );
  AND3_X1 CU_I_U29 ( .A1(IRAM_DATA[28]), .A2(IRAM_DATA[30]), .A3(CU_I_n42), 
        .ZN(CU_I_n180) );
  NAND2_X2 CU_I_U28 ( .A1(IRAM_DATA[29]), .A2(CU_I_n266), .ZN(CU_I_n157) );
  NAND2_X1 CU_I_U27 ( .A1(CU_I_n26), .A2(CU_I_n14), .ZN(CU_I_n171) );
  INV_X1 CU_I_U26 ( .A(CU_I_n39), .ZN(alu_op_i[0]) );
  INV_X2 CU_I_U25 ( .A(CU_I_n69), .ZN(pipe_ex_mem_en_i) );
  NOR3_X1 CU_I_U24 ( .A1(IRAM_DATA[28]), .A2(IRAM_DATA[30]), .A3(CU_I_n157), 
        .ZN(CU_I_n38) );
  INV_X1 CU_I_U23 ( .A(CU_I_n28), .ZN(CU_I_n29) );
  NAND2_X1 CU_I_U22 ( .A1(CU_I_n87), .A2(CU_I_n29), .ZN(CU_I_n194) );
  NAND3_X1 CU_I_U21 ( .A1(CU_I_n100), .A2(CU_I_n155), .A3(CU_I_n269), .ZN(
        CU_I_n28) );
  OAI221_X4 CU_I_U20 ( .B1(CU_I_n63), .B2(CU_I_n8), .C1(pipe_if_id_en_i), .C2(
        CU_I_n16), .A(CU_I_n80), .ZN(CU_I_n231) );
  AND2_X2 CU_I_U19 ( .A1(IRAM_DATA[27]), .A2(IRAM_DATA[26]), .ZN(CU_I_n154) );
  INV_X1 CU_I_U18 ( .A(CU_I_n45), .ZN(muxB_sel_i) );
  NOR3_X1 CU_I_U17 ( .A1(CU_I_n185), .A2(CU_I_n186), .A3(CU_I_n18), .ZN(
        CU_I_n183) );
  INV_X1 CU_I_U16 ( .A(CU_I_n24), .ZN(CU_I_n25) );
  NOR2_X1 CU_I_U15 ( .A1(CU_I_n133), .A2(CU_I_n28), .ZN(CU_I_n20) );
  AND2_X1 CU_I_U14 ( .A1(CU_I_n20), .A2(CU_I_n87), .ZN(CU_I_n203) );
  INV_X2 CU_I_U13 ( .A(RST), .ZN(CU_I_n256) );
  OR2_X1 CU_I_U12 ( .A1(CU_I_n184), .A2(CU_I_n257), .ZN(CU_I_n18) );
  AND2_X1 CU_I_U11 ( .A1(CU_I_n178), .A2(CU_I_n177), .ZN(CU_I_n14) );
  OR3_X1 CU_I_U10 ( .A1(CU_I_n267), .A2(CU_I_n70), .A3(CU_I_n176), .ZN(CU_I_n1) );
  BUF_X1 CU_I_U9 ( .A(CU_I_n78), .Z(CU_I_n58) );
  OAI221_X1 CU_I_U8 ( .B1(CU_I_n188), .B2(CU_I_n51), .C1(pipe_if_id_en_i), 
        .C2(CU_I_n3), .A(CU_I_n182), .ZN(CU_I_n246) );
  NOR2_X1 CU_I_U7 ( .A1(DRAM_READY), .A2(CU_I_n27), .ZN(DRAM_ISSUE) );
  INV_X1 CU_I_U6 ( .A(IRAM_DATA[3]), .ZN(CU_I_n288) );
  AND2_X1 CU_I_U5 ( .A1(CU_I_n191), .A2(CU_I_n114), .ZN(CU_I_n26) );
  AND4_X1 CU_I_U4 ( .A1(CU_I_n89), .A2(CU_I_n115), .A3(CU_I_n116), .A4(
        CU_I_n203), .ZN(CU_I_n191) );
  OAI221_X1 CU_I_U3 ( .B1(IRAM_DATA[27]), .B2(CU_I_n275), .C1(CU_I_n157), .C2(
        CU_I_n277), .A(CU_I_n158), .ZN(CU_I_n156) );
  DFFR_X1 CU_I_cw1_reg_17_ ( .D(CU_I_n252), .CK(CLK), .RN(CU_I_n256), .Q(
        rf_rs1_en_i) );
  DFFR_X1 CU_I_cw1_reg_12_ ( .D(CU_I_n247), .CK(CLK), .RN(CU_I_n256), .Q(
        regrd_sel_i) );
  DFFR_X1 CU_I_cw1_reg_14_ ( .D(CU_I_n249), .CK(CLK), .RN(CU_I_n256), .Q(
        imm_uns_i) );
  DFFR_X1 CU_I_cw1_reg_15_ ( .D(CU_I_n250), .CK(CLK), .RN(CU_I_n256), .Q(
        imm_isoff_i) );
  DFFR_X1 CU_I_cw1_reg_16_ ( .D(CU_I_n251), .CK(CLK), .RN(CU_I_n256), .Q(
        rf_rs2_en_i) );
  DFFR_X1 CU_I_aluOpcode2_reg_1_ ( .D(CU_I_n212), .CK(CLK), .RN(CU_I_n256), 
        .Q(alu_op_i[1]) );
  DFFR_X1 CU_I_cw2_reg_8_ ( .D(CU_I_n229), .CK(CLK), .RN(CU_I_n256), .Q(
        npc_wb_en_i) );
  DFFR_X1 CU_I_cw2_reg_9_ ( .D(CU_I_n228), .CK(CLK), .RN(CU_I_n256), .Q(
        mem_in_en_i) );
  DFFR_X1 CU_I_cw4_reg_1_ ( .D(CU_I_n221), .CK(CLK), .RN(CU_I_n256), .Q(
        rf_we_i) );
  DFFR_X1 CU_I_cw4_reg_2_ ( .D(CU_I_n222), .CK(CLK), .RN(CU_I_n256), .Q(
        wb_mux_sel_i) );
  DFFR_X1 CU_I_cw3_reg_4_ ( .D(CU_I_n72), .CK(CLK), .RN(CU_I_n256), .Q(
        CU_I_cw3_4_) );
  DFFR_X1 CU_I_cw3_reg_5_ ( .D(CU_I_n73), .CK(CLK), .RN(CU_I_n256), .Q(
        CU_I_cw3_5_) );
  DFFR_X1 CU_I_cw1_reg_2_ ( .D(CU_I_n237), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n12) );
  DFFR_X1 CU_I_cw1_reg_11_ ( .D(CU_I_n246), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n3) );
  DFFR_X1 CU_I_aluOpcode1_reg_0_ ( .D(CU_I_n216), .CK(CLK), .RN(CU_I_n256), 
        .QN(CU_I_n37) );
  DFFR_X1 CU_I_cw1_reg_8_ ( .D(CU_I_n243), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n6) );
  DFFR_X1 CU_I_cw1_reg_4_ ( .D(CU_I_n239), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n10) );
  DFFR_X1 CU_I_cw1_reg_5_ ( .D(CU_I_n240), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n9) );
  DFFR_X1 CU_I_cw1_reg_9_ ( .D(CU_I_n244), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n5) );
  DFFR_X1 CU_I_cw2_reg_1_ ( .D(CU_I_n236), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n23) );
  DFFR_X1 CU_I_cw2_reg_2_ ( .D(CU_I_n235), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n22) );
  DFFR_X1 CU_I_cw2_reg_3_ ( .D(CU_I_n234), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n21) );
  DFFR_X1 CU_I_cw2_reg_7_ ( .D(CU_I_n230), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n15) );
  DFFR_X1 CU_I_cw3_reg_1_ ( .D(CU_I_n223), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n32) );
  DFFR_X1 CU_I_cw3_reg_2_ ( .D(CU_I_n224), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n31) );
  DFFR_X1 CU_I_cw3_reg_3_ ( .D(CU_I_n225), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n30) );
  DFFR_X1 CU_I_cw3_reg_7_ ( .D(CU_I_n254), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n27) );
  DFFR_X1 CU_I_cw1_reg_3_ ( .D(CU_I_n238), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n11) );
  DFFR_X1 CU_I_cw1_reg_7_ ( .D(CU_I_n242), .CK(CLK), .RN(CU_I_n256), .QN(
        CU_I_n7) );
  DFFS_X1 CU_I_aluOpcode2_reg_2_ ( .D(CU_I_n213), .CK(CLK), .SN(CU_I_n256), 
        .Q(alu_op_i[2]) );
  DFFS_X2 CU_I_aluOpcode2_reg_4_ ( .D(CU_I_n215), .CK(CLK), .SN(CU_I_n55), .Q(
        alu_op_i[4]), .QN(CU_I_n24) );
  NAND3_X1 CU_I_U231 ( .A1(CU_I_n117), .A2(IRAM_DATA[28]), .A3(CU_I_n205), 
        .ZN(CU_I_n130) );
  NAND3_X1 CU_I_U230 ( .A1(CU_I_n154), .A2(CU_I_n276), .A3(CU_I_n205), .ZN(
        CU_I_n127) );
  NAND3_X1 CU_I_U229 ( .A1(CU_I_n132), .A2(CU_I_n276), .A3(CU_I_n205), .ZN(
        CU_I_n140) );
  NAND3_X1 CU_I_U228 ( .A1(CU_I_n134), .A2(CU_I_n101), .A3(CU_I_n140), .ZN(
        CU_I_n204) );
  NAND3_X1 CU_I_U227 ( .A1(CU_I_n160), .A2(IRAM_DATA[28]), .A3(CU_I_n202), 
        .ZN(CU_I_n174) );
  NAND3_X1 CU_I_U226 ( .A1(CU_I_n117), .A2(IRAM_DATA[28]), .A3(CU_I_n202), 
        .ZN(CU_I_n173) );
  NAND3_X1 CU_I_U225 ( .A1(CU_I_n201), .A2(CU_I_n154), .A3(CU_I_n161), .ZN(
        CU_I_n178) );
  NAND3_X1 CU_I_U224 ( .A1(CU_I_n189), .A2(CU_I_n196), .A3(CU_I_n177), .ZN(
        CU_I_n186) );
  NAND3_X1 CU_I_U222 ( .A1(IRAM_DATA[28]), .A2(IRAM_DATA[29]), .A3(
        IRAM_DATA[27]), .ZN(CU_I_n158) );
  NAND3_X1 CU_I_U221 ( .A1(CU_I_n129), .A2(CU_I_n130), .A3(CU_I_n131), .ZN(
        CU_I_n124) );
  OAI33_X1 CU_I_U220 ( .A1(CU_I_n286), .A2(CU_I_n291), .A3(CU_I_n289), .B1(
        IRAM_DATA[0]), .B2(IRAM_DATA[4]), .B3(IRAM_DATA[2]), .ZN(CU_I_n126) );
  OAI33_X1 CU_I_U219 ( .A1(CU_I_n270), .A2(IRAM_DATA[0]), .A3(CU_I_n288), .B1(
        CU_I_n272), .B2(IRAM_DATA[1]), .B3(CU_I_n285), .ZN(CU_I_n125) );
  NAND3_X1 CU_I_U218 ( .A1(CU_I_n103), .A2(CU_I_n89), .A3(CU_I_n104), .ZN(
        CU_I_n96) );
  NAND3_X1 CU_I_U217 ( .A1(CU_I_n100), .A2(CU_I_n101), .A3(CU_I_n102), .ZN(
        CU_I_n97) );
  OAI33_X1 CU_I_U216 ( .A1(CU_I_n286), .A2(IRAM_DATA[2]), .A3(CU_I_n290), .B1(
        CU_I_n289), .B2(IRAM_DATA[1]), .B3(CU_I_n291), .ZN(CU_I_n92) );
  DFFR_X1 CU_I_aluOpcode2_reg_0_ ( .D(CU_I_n211), .CK(CLK), .RN(CU_I_n53), .Q(
        CU_I_n294), .QN(CU_I_n39) );
  DFFR_X1 CU_I_aluOpcode2_reg_3_ ( .D(CU_I_n214), .CK(CLK), .RN(CU_I_n52), .Q(
        alu_op_i[3]) );
  DFFR_X1 CU_I_aluOpcode1_reg_1_ ( .D(CU_I_n217), .CK(CLK), .RN(CU_I_n52), 
        .QN(CU_I_n36) );
  DFFS_X1 CU_I_aluOpcode1_reg_2_ ( .D(CU_I_n218), .CK(CLK), .SN(CU_I_n55), 
        .QN(CU_I_n35) );
  DFFR_X1 CU_I_aluOpcode1_reg_3_ ( .D(CU_I_n219), .CK(CLK), .RN(CU_I_n52), 
        .QN(CU_I_n34) );
  DFFS_X1 CU_I_aluOpcode1_reg_4_ ( .D(CU_I_n220), .CK(CLK), .SN(CU_I_n55), 
        .QN(CU_I_n33) );
  DFFR_X1 CU_I_cw1_reg_1_ ( .D(CU_I_n74), .CK(CLK), .RN(CU_I_n53), .Q(
        CU_I_cw1_1_), .QN(CU_I_n13) );
  DFFS_X1 CU_I_cw3_reg_6_ ( .D(CU_I_n253), .CK(CLK), .SN(CU_I_n55), .Q(
        DRAM_READNOTWRITE) );
  DFFS_X1 CU_I_cw2_reg_6_ ( .D(CU_I_n231), .CK(CLK), .SN(CU_I_n55), .QN(
        CU_I_n16) );
  DFFS_X1 CU_I_cw1_reg_6_ ( .D(CU_I_n241), .CK(CLK), .SN(CU_I_n55), .QN(
        CU_I_n8) );
  DFFR_X1 CU_I_cw2_reg_10_ ( .D(CU_I_n227), .CK(CLK), .RN(CU_I_n53), .Q(
        CU_I_n293), .QN(CU_I_n45) );
  DFFR_X1 CU_I_cw2_reg_11_ ( .D(CU_I_n226), .CK(CLK), .RN(CU_I_n54), .Q(
        CU_I_n292), .QN(CU_I_n43) );
  DFFR_X1 CU_I_cw1_reg_13_ ( .D(CU_I_n248), .CK(CLK), .RN(CU_I_n53), .Q(
        reg31_sel_i), .QN(CU_I_n2) );
  DFFR_X1 CU_I_cw1_reg_10_ ( .D(CU_I_n245), .CK(CLK), .RN(CU_I_n54), .QN(
        CU_I_n4) );
  DFFR_X1 CU_I_cw2_reg_5_ ( .D(CU_I_n232), .CK(CLK), .RN(CU_I_n54), .Q(
        CU_I_cw2[5]), .QN(CU_I_n17) );
  DFFR_X1 CU_I_cw2_reg_4_ ( .D(CU_I_n233), .CK(CLK), .RN(CU_I_n54), .Q(
        CU_I_cw2[4]), .QN(CU_I_n19) );
  INV_X1 dp_U792 ( .A(dp_n141), .ZN(dp_n941) );
  AOI22_X1 dp_U791 ( .A1(dp_alu_out_ex_o[0]), .A2(dp_n15), .B1(dp_n17), .B2(
        DRAM_ADDRESS[0]), .ZN(dp_n141) );
  OAI21_X1 dp_U790 ( .B1(dp_n558), .B2(dp_n110), .A(dp_n140), .ZN(dp_n691) );
  NAND2_X1 dp_U789 ( .A1(dp_npc_if_o[16]), .A2(dp_n104), .ZN(dp_n140) );
  OAI21_X1 dp_U788 ( .B1(dp_n559), .B2(dp_n110), .A(dp_n139), .ZN(dp_n692) );
  NAND2_X1 dp_U787 ( .A1(dp_npc_if_o[17]), .A2(dp_n104), .ZN(dp_n139) );
  OAI21_X1 dp_U786 ( .B1(dp_n560), .B2(dp_n110), .A(dp_n138), .ZN(dp_n693) );
  NAND2_X1 dp_U785 ( .A1(dp_npc_if_o[18]), .A2(dp_n104), .ZN(dp_n138) );
  OAI21_X1 dp_U784 ( .B1(dp_n561), .B2(dp_n110), .A(dp_n137), .ZN(dp_n694) );
  NAND2_X1 dp_U783 ( .A1(dp_npc_if_o[19]), .A2(dp_n104), .ZN(dp_n137) );
  OAI21_X1 dp_U782 ( .B1(dp_n562), .B2(dp_n110), .A(dp_n136), .ZN(dp_n695) );
  NAND2_X1 dp_U781 ( .A1(dp_npc_if_o[20]), .A2(dp_n104), .ZN(dp_n136) );
  OAI21_X1 dp_U780 ( .B1(dp_n563), .B2(dp_n110), .A(dp_n135), .ZN(dp_n696) );
  NAND2_X1 dp_U779 ( .A1(dp_npc_if_o[21]), .A2(dp_n104), .ZN(dp_n135) );
  OAI21_X1 dp_U778 ( .B1(dp_n564), .B2(dp_n110), .A(dp_n134), .ZN(dp_n697) );
  NAND2_X1 dp_U777 ( .A1(dp_npc_if_o[22]), .A2(dp_n104), .ZN(dp_n134) );
  OAI21_X1 dp_U776 ( .B1(dp_n565), .B2(dp_n110), .A(dp_n133), .ZN(dp_n698) );
  NAND2_X1 dp_U775 ( .A1(dp_npc_if_o[23]), .A2(dp_n104), .ZN(dp_n133) );
  OAI21_X1 dp_U774 ( .B1(dp_n566), .B2(dp_n110), .A(dp_n130), .ZN(dp_n699) );
  NAND2_X1 dp_U773 ( .A1(dp_npc_if_o[24]), .A2(dp_n104), .ZN(dp_n130) );
  OAI21_X1 dp_U772 ( .B1(dp_n567), .B2(dp_n111), .A(dp_n129), .ZN(dp_n700) );
  NAND2_X1 dp_U771 ( .A1(dp_npc_if_o[25]), .A2(dp_n104), .ZN(dp_n129) );
  OAI21_X1 dp_U770 ( .B1(dp_n568), .B2(dp_n110), .A(dp_n128), .ZN(dp_n701) );
  NAND2_X1 dp_U769 ( .A1(dp_npc_if_o[26]), .A2(dp_n104), .ZN(dp_n128) );
  OAI21_X1 dp_U768 ( .B1(dp_n569), .B2(dp_n110), .A(dp_n127), .ZN(dp_n702) );
  NAND2_X1 dp_U767 ( .A1(dp_npc_if_o[27]), .A2(dp_n104), .ZN(dp_n127) );
  OAI21_X1 dp_U766 ( .B1(dp_n570), .B2(dp_n111), .A(dp_n126), .ZN(dp_n703) );
  NAND2_X1 dp_U765 ( .A1(dp_npc_if_o[28]), .A2(dp_n104), .ZN(dp_n126) );
  OAI21_X1 dp_U764 ( .B1(dp_n571), .B2(dp_n111), .A(dp_n125), .ZN(dp_n704) );
  NAND2_X1 dp_U763 ( .A1(dp_npc_if_o[29]), .A2(dp_n104), .ZN(dp_n125) );
  OAI21_X1 dp_U762 ( .B1(dp_n572), .B2(dp_n111), .A(dp_n124), .ZN(dp_n705) );
  NAND2_X1 dp_U761 ( .A1(dp_npc_if_o[30]), .A2(dp_n104), .ZN(dp_n124) );
  OAI21_X1 dp_U760 ( .B1(dp_n573), .B2(dp_n111), .A(dp_n123), .ZN(dp_n706) );
  NAND2_X1 dp_U759 ( .A1(dp_npc_if_o[31]), .A2(dp_n103), .ZN(dp_n123) );
  OR2_X1 dp_U758 ( .A1(pipe_if_id_en_i), .A2(dp_n142), .ZN(dp_n68) );
  INV_X1 dp_U757 ( .A(pipe_clear_n_i), .ZN(dp_n142) );
  INV_X1 dp_U756 ( .A(dp_n121), .ZN(dp_n114) );
  INV_X1 dp_U755 ( .A(pipe_ex_mem_en_i), .ZN(dp_n112) );
  INV_X1 dp_U754 ( .A(dp_n103), .ZN(dp_n102) );
  CLKBUF_X1 dp_U751 ( .A(dp_n89), .Z(dp_n99) );
  CLKBUF_X1 dp_U750 ( .A(dp_n22), .Z(dp_n45) );
  CLKBUF_X1 dp_U749 ( .A(dp_n22), .Z(dp_n44) );
  CLKBUF_X1 dp_U748 ( .A(dp_n21), .Z(dp_n43) );
  CLKBUF_X1 dp_U747 ( .A(dp_n21), .Z(dp_n42) );
  CLKBUF_X1 dp_U746 ( .A(dp_n21), .Z(dp_n41) );
  CLKBUF_X1 dp_U745 ( .A(dp_n21), .Z(dp_n40) );
  CLKBUF_X1 dp_U744 ( .A(dp_n21), .Z(dp_n39) );
  CLKBUF_X1 dp_U743 ( .A(dp_n21), .Z(dp_n38) );
  CLKBUF_X1 dp_U742 ( .A(dp_n20), .Z(dp_n37) );
  CLKBUF_X1 dp_U741 ( .A(dp_n20), .Z(dp_n36) );
  CLKBUF_X1 dp_U740 ( .A(dp_n20), .Z(dp_n35) );
  CLKBUF_X1 dp_U739 ( .A(dp_n19), .Z(dp_n34) );
  CLKBUF_X1 dp_U738 ( .A(dp_n19), .Z(dp_n33) );
  CLKBUF_X1 dp_U737 ( .A(dp_n19), .Z(dp_n32) );
  CLKBUF_X1 dp_U736 ( .A(dp_n19), .Z(dp_n31) );
  CLKBUF_X1 dp_U735 ( .A(dp_n18), .Z(dp_n30) );
  CLKBUF_X1 dp_U734 ( .A(dp_n18), .Z(dp_n29) );
  CLKBUF_X1 dp_U733 ( .A(dp_n18), .Z(dp_n28) );
  CLKBUF_X1 dp_U732 ( .A(dp_n18), .Z(dp_n27) );
  CLKBUF_X1 dp_U731 ( .A(dp_n18), .Z(dp_n26) );
  CLKBUF_X1 dp_U730 ( .A(dp_n18), .Z(dp_n25) );
  OAI22_X1 dp_U729 ( .A1(dp_n857), .A2(dp_n72), .B1(dp_n67), .B2(dp_n169), 
        .ZN(dp_n921) );
  OAI22_X1 dp_U728 ( .A1(dp_n851), .A2(dp_n71), .B1(dp_n163), .B2(dp_n67), 
        .ZN(dp_n915) );
  INV_X1 dp_U727 ( .A(dp_alu_out_ex_o[25]), .ZN(dp_n164) );
  OAI22_X1 dp_U726 ( .A1(dp_n852), .A2(dp_n71), .B1(dp_n164), .B2(dp_n67), 
        .ZN(dp_n916) );
  INV_X1 dp_U725 ( .A(dp_alu_out_ex_o[30]), .ZN(dp_n159) );
  OAI22_X1 dp_U724 ( .A1(dp_n853), .A2(dp_n71), .B1(dp_n67), .B2(dp_n165), 
        .ZN(dp_n917) );
  INV_X1 dp_U723 ( .A(dp_alu_out_ex_o[21]), .ZN(dp_n168) );
  INV_X1 dp_U722 ( .A(dp_alu_out_ex_o[29]), .ZN(dp_n160) );
  OAI22_X1 dp_U721 ( .A1(dp_n848), .A2(dp_n71), .B1(dp_n160), .B2(dp_n67), 
        .ZN(dp_n912) );
  INV_X1 dp_U720 ( .A(dp_alu_out_ex_o[28]), .ZN(dp_n161) );
  INV_X1 dp_U719 ( .A(dp_alu_out_ex_o[22]), .ZN(dp_n167) );
  INV_X1 dp_U718 ( .A(dp_alu_out_ex_o[24]), .ZN(dp_n165) );
  INV_X1 dp_U717 ( .A(dp_alu_out_ex_o[27]), .ZN(dp_n162) );
  OAI22_X1 dp_U716 ( .A1(dp_n850), .A2(dp_n71), .B1(dp_n67), .B2(dp_n162), 
        .ZN(dp_n914) );
  INV_X1 dp_U715 ( .A(dp_alu_out_ex_o[26]), .ZN(dp_n163) );
  OAI22_X1 dp_U714 ( .A1(dp_n847), .A2(dp_n71), .B1(dp_n159), .B2(dp_n67), 
        .ZN(dp_n911) );
  OAI22_X1 dp_U713 ( .A1(dp_n856), .A2(dp_n71), .B1(dp_n67), .B2(dp_n168), 
        .ZN(dp_n920) );
  INV_X1 dp_U712 ( .A(dp_alu_out_ex_o[20]), .ZN(dp_n169) );
  INV_X1 dp_U711 ( .A(dp_alu_out_ex_o[31]), .ZN(dp_n158) );
  INV_X1 dp_U710 ( .A(dp_alu_out_ex_o[23]), .ZN(dp_n166) );
  OAI22_X1 dp_U709 ( .A1(dp_n854), .A2(dp_n71), .B1(dp_n67), .B2(dp_n166), 
        .ZN(dp_n918) );
  OAI22_X1 dp_U708 ( .A1(dp_n849), .A2(dp_n71), .B1(dp_n161), .B2(dp_n67), 
        .ZN(dp_n913) );
  OAI22_X1 dp_U707 ( .A1(dp_n855), .A2(dp_n71), .B1(dp_n167), .B2(dp_n67), 
        .ZN(dp_n919) );
  OAI22_X1 dp_U706 ( .A1(dp_n846), .A2(dp_n71), .B1(dp_n158), .B2(dp_n67), 
        .ZN(dp_n910) );
  INV_X1 dp_U705 ( .A(dp_alu_out_ex_o[5]), .ZN(dp_n184) );
  INV_X1 dp_U704 ( .A(dp_alu_out_ex_o[4]), .ZN(dp_n185) );
  INV_X1 dp_U703 ( .A(wb_mux_sel_i), .ZN(dp_n122) );
  INV_X1 dp_U702 ( .A(mem_in_en_i), .ZN(dp_n1027) );
  INV_X1 dp_U701 ( .A(DRAM_DATA[0]), .ZN(dp_n400) );
  INV_X1 dp_U700 ( .A(DRAM_DATA[1]), .ZN(dp_n365) );
  INV_X1 dp_U699 ( .A(DRAM_DATA[2]), .ZN(dp_n364) );
  INV_X1 dp_U698 ( .A(DRAM_DATA[3]), .ZN(dp_n363) );
  INV_X1 dp_U697 ( .A(DRAM_DATA[4]), .ZN(dp_n362) );
  INV_X1 dp_U696 ( .A(DRAM_DATA[5]), .ZN(dp_n361) );
  INV_X1 dp_U695 ( .A(DRAM_DATA[6]), .ZN(dp_n360) );
  INV_X1 dp_U694 ( .A(DRAM_DATA[7]), .ZN(dp_n359) );
  INV_X1 dp_U693 ( .A(DRAM_DATA[8]), .ZN(dp_n358) );
  INV_X1 dp_U692 ( .A(DRAM_DATA[9]), .ZN(dp_n357) );
  INV_X1 dp_U691 ( .A(DRAM_DATA[10]), .ZN(dp_n356) );
  INV_X1 dp_U690 ( .A(DRAM_DATA[11]), .ZN(dp_n355) );
  INV_X1 dp_U689 ( .A(DRAM_DATA[12]), .ZN(dp_n354) );
  INV_X1 dp_U688 ( .A(DRAM_DATA[13]), .ZN(dp_n353) );
  INV_X1 dp_U687 ( .A(DRAM_DATA[14]), .ZN(dp_n352) );
  INV_X1 dp_U686 ( .A(DRAM_DATA[15]), .ZN(dp_n351) );
  INV_X1 dp_U685 ( .A(DRAM_DATA[16]), .ZN(dp_n350) );
  INV_X1 dp_U684 ( .A(DRAM_DATA[17]), .ZN(dp_n349) );
  INV_X1 dp_U683 ( .A(DRAM_DATA[18]), .ZN(dp_n348) );
  INV_X1 dp_U682 ( .A(DRAM_DATA[19]), .ZN(dp_n347) );
  INV_X1 dp_U681 ( .A(DRAM_DATA[20]), .ZN(dp_n346) );
  INV_X1 dp_U680 ( .A(DRAM_DATA[21]), .ZN(dp_n345) );
  INV_X1 dp_U679 ( .A(DRAM_DATA[22]), .ZN(dp_n344) );
  INV_X1 dp_U678 ( .A(DRAM_DATA[23]), .ZN(dp_n343) );
  INV_X1 dp_U677 ( .A(DRAM_DATA[24]), .ZN(dp_n342) );
  INV_X1 dp_U676 ( .A(DRAM_DATA[25]), .ZN(dp_n341) );
  INV_X1 dp_U675 ( .A(DRAM_DATA[26]), .ZN(dp_n340) );
  INV_X1 dp_U674 ( .A(DRAM_DATA[27]), .ZN(dp_n339) );
  INV_X1 dp_U673 ( .A(DRAM_DATA[28]), .ZN(dp_n338) );
  INV_X1 dp_U672 ( .A(DRAM_DATA[29]), .ZN(dp_n337) );
  INV_X1 dp_U671 ( .A(DRAM_DATA[30]), .ZN(dp_n336) );
  INV_X1 dp_U670 ( .A(DRAM_DATA[31]), .ZN(dp_n335) );
  OAI22_X1 dp_U669 ( .A1(dp_n331), .A2(dp_n63), .B1(dp_n877), .B2(dp_n57), 
        .ZN(dp_n909) );
  OAI22_X1 dp_U668 ( .A1(dp_n525), .A2(dp_n65), .B1(dp_n857), .B2(dp_n55), 
        .ZN(dp_n889) );
  OAI22_X1 dp_U667 ( .A1(dp_n584), .A2(dp_n65), .B1(dp_n856), .B2(dp_n55), 
        .ZN(dp_n888) );
  OAI22_X1 dp_U666 ( .A1(dp_n585), .A2(dp_n65), .B1(dp_n855), .B2(dp_n55), 
        .ZN(dp_n887) );
  OAI22_X1 dp_U665 ( .A1(dp_n586), .A2(dp_n65), .B1(dp_n854), .B2(dp_n55), 
        .ZN(dp_n886) );
  OAI22_X1 dp_U664 ( .A1(dp_n587), .A2(dp_n65), .B1(dp_n853), .B2(dp_n55), 
        .ZN(dp_n885) );
  OAI22_X1 dp_U663 ( .A1(dp_n588), .A2(dp_n65), .B1(dp_n852), .B2(dp_n55), 
        .ZN(dp_n884) );
  OAI22_X1 dp_U662 ( .A1(dp_n589), .A2(dp_n66), .B1(dp_n851), .B2(dp_n55), 
        .ZN(dp_n883) );
  OAI22_X1 dp_U661 ( .A1(dp_n590), .A2(dp_n66), .B1(dp_n850), .B2(dp_n55), 
        .ZN(dp_n882) );
  OAI22_X1 dp_U660 ( .A1(dp_n591), .A2(dp_n66), .B1(dp_n849), .B2(dp_n55), 
        .ZN(dp_n881) );
  OAI22_X1 dp_U659 ( .A1(dp_n592), .A2(dp_n66), .B1(dp_n848), .B2(dp_n55), 
        .ZN(dp_n880) );
  OAI22_X1 dp_U658 ( .A1(dp_n593), .A2(dp_n66), .B1(dp_n847), .B2(dp_n55), 
        .ZN(dp_n879) );
  OAI22_X1 dp_U657 ( .A1(dp_n1025), .A2(dp_n61), .B1(dp_n846), .B2(dp_n55), 
        .ZN(dp_n878) );
  OAI22_X1 dp_U656 ( .A1(dp_n444), .A2(dp_n91), .B1(dp_n76), .B2(dp_n624), 
        .ZN(dp_n774) );
  OAI22_X1 dp_U655 ( .A1(dp_n445), .A2(dp_n90), .B1(dp_n78), .B2(dp_n625), 
        .ZN(dp_n775) );
  OAI22_X1 dp_U654 ( .A1(dp_n447), .A2(dp_n90), .B1(dp_n81), .B2(dp_n625), 
        .ZN(dp_n777) );
  OAI22_X1 dp_U653 ( .A1(dp_n446), .A2(dp_n90), .B1(dp_n81), .B2(dp_n624), 
        .ZN(dp_n776) );
  OAI22_X1 dp_U652 ( .A1(dp_n449), .A2(dp_n94), .B1(dp_n81), .B2(dp_n625), 
        .ZN(dp_n779) );
  INV_X1 dp_U651 ( .A(dp_imm_id_o[31]), .ZN(dp_n625) );
  OAI22_X1 dp_U650 ( .A1(dp_n450), .A2(dp_n93), .B1(dp_n79), .B2(dp_n625), 
        .ZN(dp_n780) );
  INV_X1 dp_U649 ( .A(dp_imm_id_o[31]), .ZN(dp_n624) );
  OAI22_X1 dp_U648 ( .A1(dp_n448), .A2(dp_n94), .B1(dp_n80), .B2(dp_n624), 
        .ZN(dp_n778) );
  OAI221_X1 dp_U647 ( .B1(dp_n575), .B2(regrd_sel_i), .C1(dp_n574), .C2(
        dp_n1028), .A(dp_n1026), .ZN(dp_rd_fwd_id_o[0]) );
  INV_X1 dp_U646 ( .A(dp_rd_fwd_id_o[0]), .ZN(dp_n605) );
  OAI22_X1 dp_U645 ( .A1(dp_n93), .A2(dp_n414), .B1(dp_n80), .B2(dp_n605), 
        .ZN(dp_n712) );
  INV_X1 dp_U644 ( .A(dp_imm_id_o[22]), .ZN(dp_n621) );
  OAI22_X1 dp_U643 ( .A1(dp_n441), .A2(dp_n90), .B1(dp_n79), .B2(dp_n621), 
        .ZN(dp_n771) );
  INV_X1 dp_U642 ( .A(dp_alu_out_ex_o[19]), .ZN(dp_n170) );
  OAI22_X1 dp_U641 ( .A1(dp_n858), .A2(dp_n72), .B1(dp_n170), .B2(dp_n67), 
        .ZN(dp_n922) );
  INV_X1 dp_U640 ( .A(dp_rf_out2_id_o[3]), .ZN(dp_n245) );
  OAI22_X1 dp_U639 ( .A1(dp_n96), .A2(dp_n454), .B1(dp_n83), .B2(dp_n245), 
        .ZN(dp_n784) );
  INV_X1 dp_U638 ( .A(dp_rf_out2_id_o[4]), .ZN(dp_n243) );
  OAI22_X1 dp_U637 ( .A1(dp_n96), .A2(dp_n455), .B1(dp_n82), .B2(dp_n243), 
        .ZN(dp_n785) );
  INV_X1 dp_U636 ( .A(dp_rf_out2_id_o[5]), .ZN(dp_n241) );
  OAI22_X1 dp_U635 ( .A1(dp_n96), .A2(dp_n456), .B1(dp_n86), .B2(dp_n241), 
        .ZN(dp_n786) );
  INV_X1 dp_U634 ( .A(dp_rf_out2_id_o[6]), .ZN(dp_n239) );
  OAI22_X1 dp_U633 ( .A1(dp_n96), .A2(dp_n457), .B1(dp_n86), .B2(dp_n239), 
        .ZN(dp_n787) );
  INV_X1 dp_U632 ( .A(dp_rf_out2_id_o[7]), .ZN(dp_n237) );
  OAI22_X1 dp_U631 ( .A1(dp_n96), .A2(dp_n458), .B1(dp_n86), .B2(dp_n237), 
        .ZN(dp_n788) );
  INV_X1 dp_U630 ( .A(dp_rf_out2_id_o[8]), .ZN(dp_n235) );
  OAI22_X1 dp_U629 ( .A1(dp_n96), .A2(dp_n459), .B1(dp_n86), .B2(dp_n235), 
        .ZN(dp_n789) );
  INV_X1 dp_U628 ( .A(dp_rf_out2_id_o[9]), .ZN(dp_n233) );
  OAI22_X1 dp_U627 ( .A1(dp_n96), .A2(dp_n460), .B1(dp_n86), .B2(dp_n233), 
        .ZN(dp_n790) );
  INV_X1 dp_U626 ( .A(dp_rf_out2_id_o[10]), .ZN(dp_n231) );
  OAI22_X1 dp_U625 ( .A1(dp_n95), .A2(dp_n461), .B1(dp_n86), .B2(dp_n231), 
        .ZN(dp_n791) );
  INV_X1 dp_U624 ( .A(dp_rf_out2_id_o[11]), .ZN(dp_n229) );
  OAI22_X1 dp_U623 ( .A1(dp_n95), .A2(dp_n462), .B1(dp_n86), .B2(dp_n229), 
        .ZN(dp_n792) );
  INV_X1 dp_U622 ( .A(dp_rf_out2_id_o[12]), .ZN(dp_n227) );
  OAI22_X1 dp_U621 ( .A1(dp_n95), .A2(dp_n463), .B1(dp_n86), .B2(dp_n227), 
        .ZN(dp_n793) );
  INV_X1 dp_U620 ( .A(dp_rf_out2_id_o[13]), .ZN(dp_n225) );
  OAI22_X1 dp_U619 ( .A1(dp_n95), .A2(dp_n464), .B1(dp_n86), .B2(dp_n225), 
        .ZN(dp_n794) );
  INV_X1 dp_U618 ( .A(dp_rf_out2_id_o[14]), .ZN(dp_n223) );
  OAI22_X1 dp_U617 ( .A1(dp_n95), .A2(dp_n465), .B1(dp_n86), .B2(dp_n223), 
        .ZN(dp_n795) );
  INV_X1 dp_U616 ( .A(dp_rf_out2_id_o[15]), .ZN(dp_n221) );
  OAI22_X1 dp_U615 ( .A1(dp_n95), .A2(dp_n466), .B1(dp_n83), .B2(dp_n221), 
        .ZN(dp_n796) );
  INV_X1 dp_U614 ( .A(dp_rf_out2_id_o[16]), .ZN(dp_n219) );
  OAI22_X1 dp_U613 ( .A1(dp_n95), .A2(dp_n467), .B1(dp_n82), .B2(dp_n219), 
        .ZN(dp_n797) );
  INV_X1 dp_U612 ( .A(dp_rf_out2_id_o[17]), .ZN(dp_n217) );
  OAI22_X1 dp_U611 ( .A1(dp_n95), .A2(dp_n468), .B1(dp_n84), .B2(dp_n217), 
        .ZN(dp_n798) );
  INV_X1 dp_U610 ( .A(dp_rf_out2_id_o[18]), .ZN(dp_n215) );
  OAI22_X1 dp_U609 ( .A1(dp_n95), .A2(dp_n469), .B1(dp_n83), .B2(dp_n215), 
        .ZN(dp_n799) );
  INV_X1 dp_U608 ( .A(dp_rf_out2_id_o[19]), .ZN(dp_n213) );
  OAI22_X1 dp_U607 ( .A1(dp_n95), .A2(dp_n470), .B1(dp_n82), .B2(dp_n213), 
        .ZN(dp_n800) );
  INV_X1 dp_U606 ( .A(dp_rf_out2_id_o[20]), .ZN(dp_n211) );
  OAI22_X1 dp_U605 ( .A1(dp_n95), .A2(dp_n471), .B1(dp_n85), .B2(dp_n211), 
        .ZN(dp_n801) );
  INV_X1 dp_U604 ( .A(dp_rf_out2_id_o[21]), .ZN(dp_n209) );
  OAI22_X1 dp_U603 ( .A1(dp_n95), .A2(dp_n472), .B1(dp_n87), .B2(dp_n209), 
        .ZN(dp_n802) );
  INV_X1 dp_U602 ( .A(dp_rf_out1_id_o[0]), .ZN(dp_n252) );
  OAI22_X1 dp_U601 ( .A1(dp_n95), .A2(dp_n483), .B1(dp_n83), .B2(dp_n252), 
        .ZN(dp_n813) );
  INV_X1 dp_U600 ( .A(dp_rf_out2_id_o[22]), .ZN(dp_n207) );
  OAI22_X1 dp_U599 ( .A1(dp_n92), .A2(dp_n473), .B1(dp_n84), .B2(dp_n207), 
        .ZN(dp_n803) );
  INV_X1 dp_U598 ( .A(dp_rf_out2_id_o[23]), .ZN(dp_n205) );
  OAI22_X1 dp_U597 ( .A1(dp_n91), .A2(dp_n474), .B1(dp_n83), .B2(dp_n205), 
        .ZN(dp_n804) );
  INV_X1 dp_U596 ( .A(dp_rf_out2_id_o[24]), .ZN(dp_n203) );
  OAI22_X1 dp_U595 ( .A1(dp_n90), .A2(dp_n475), .B1(dp_n82), .B2(dp_n203), 
        .ZN(dp_n805) );
  INV_X1 dp_U594 ( .A(dp_rf_out2_id_o[25]), .ZN(dp_n201) );
  OAI22_X1 dp_U593 ( .A1(dp_n94), .A2(dp_n476), .B1(dp_n85), .B2(dp_n201), 
        .ZN(dp_n806) );
  INV_X1 dp_U592 ( .A(dp_rf_out2_id_o[26]), .ZN(dp_n199) );
  OAI22_X1 dp_U591 ( .A1(dp_n93), .A2(dp_n477), .B1(dp_n87), .B2(dp_n199), 
        .ZN(dp_n807) );
  INV_X1 dp_U590 ( .A(dp_rf_out2_id_o[27]), .ZN(dp_n197) );
  OAI22_X1 dp_U589 ( .A1(dp_n92), .A2(dp_n478), .B1(dp_n82), .B2(dp_n197), 
        .ZN(dp_n808) );
  INV_X1 dp_U588 ( .A(dp_rf_out2_id_o[28]), .ZN(dp_n195) );
  OAI22_X1 dp_U587 ( .A1(dp_n94), .A2(dp_n479), .B1(dp_n84), .B2(dp_n195), 
        .ZN(dp_n809) );
  INV_X1 dp_U586 ( .A(dp_rf_out2_id_o[29]), .ZN(dp_n193) );
  OAI22_X1 dp_U585 ( .A1(dp_n93), .A2(dp_n480), .B1(dp_n87), .B2(dp_n193), 
        .ZN(dp_n810) );
  INV_X1 dp_U584 ( .A(dp_rf_out2_id_o[30]), .ZN(dp_n191) );
  OAI22_X1 dp_U583 ( .A1(dp_n91), .A2(dp_n481), .B1(dp_n85), .B2(dp_n191), 
        .ZN(dp_n811) );
  INV_X1 dp_U582 ( .A(dp_rf_out2_id_o[31]), .ZN(dp_n189) );
  OAI22_X1 dp_U581 ( .A1(dp_n94), .A2(dp_n482), .B1(dp_n83), .B2(dp_n189), 
        .ZN(dp_n812) );
  INV_X1 dp_U580 ( .A(dp_rf_out1_id_o[1]), .ZN(dp_n250) );
  OAI22_X1 dp_U579 ( .A1(dp_n93), .A2(dp_n484), .B1(dp_n82), .B2(dp_n250), 
        .ZN(dp_n814) );
  INV_X1 dp_U578 ( .A(dp_rf_out1_id_o[2]), .ZN(dp_n248) );
  OAI22_X1 dp_U577 ( .A1(dp_n90), .A2(dp_n485), .B1(dp_n84), .B2(dp_n248), 
        .ZN(dp_n815) );
  INV_X1 dp_U576 ( .A(dp_rf_out1_id_o[3]), .ZN(dp_n246) );
  OAI22_X1 dp_U575 ( .A1(dp_n90), .A2(dp_n486), .B1(dp_n84), .B2(dp_n246), 
        .ZN(dp_n816) );
  INV_X1 dp_U574 ( .A(dp_rf_out1_id_o[4]), .ZN(dp_n244) );
  OAI22_X1 dp_U573 ( .A1(dp_n92), .A2(dp_n487), .B1(dp_n87), .B2(dp_n244), 
        .ZN(dp_n817) );
  INV_X1 dp_U572 ( .A(dp_rf_out1_id_o[5]), .ZN(dp_n242) );
  OAI22_X1 dp_U571 ( .A1(dp_n90), .A2(dp_n488), .B1(dp_n85), .B2(dp_n242), 
        .ZN(dp_n818) );
  INV_X1 dp_U570 ( .A(dp_rf_out1_id_o[6]), .ZN(dp_n240) );
  OAI22_X1 dp_U569 ( .A1(dp_n91), .A2(dp_n489), .B1(dp_n82), .B2(dp_n240), 
        .ZN(dp_n819) );
  INV_X1 dp_U568 ( .A(dp_rf_out1_id_o[7]), .ZN(dp_n238) );
  OAI22_X1 dp_U567 ( .A1(dp_n90), .A2(dp_n490), .B1(dp_n83), .B2(dp_n238), 
        .ZN(dp_n820) );
  INV_X1 dp_U566 ( .A(dp_rf_out1_id_o[8]), .ZN(dp_n236) );
  OAI22_X1 dp_U565 ( .A1(dp_n93), .A2(dp_n491), .B1(dp_n84), .B2(dp_n236), 
        .ZN(dp_n821) );
  INV_X1 dp_U564 ( .A(dp_rf_out1_id_o[9]), .ZN(dp_n234) );
  OAI22_X1 dp_U563 ( .A1(dp_n92), .A2(dp_n492), .B1(dp_n87), .B2(dp_n234), 
        .ZN(dp_n822) );
  INV_X1 dp_U562 ( .A(dp_rf_out1_id_o[10]), .ZN(dp_n232) );
  OAI22_X1 dp_U561 ( .A1(dp_n90), .A2(dp_n493), .B1(dp_n85), .B2(dp_n232), 
        .ZN(dp_n823) );
  INV_X1 dp_U560 ( .A(dp_rf_out1_id_o[11]), .ZN(dp_n230) );
  OAI22_X1 dp_U559 ( .A1(dp_n91), .A2(dp_n494), .B1(dp_n84), .B2(dp_n230), 
        .ZN(dp_n824) );
  INV_X1 dp_U558 ( .A(dp_rf_out1_id_o[12]), .ZN(dp_n228) );
  OAI22_X1 dp_U557 ( .A1(dp_n90), .A2(dp_n495), .B1(dp_n83), .B2(dp_n228), 
        .ZN(dp_n825) );
  INV_X1 dp_U556 ( .A(dp_rf_out1_id_o[13]), .ZN(dp_n226) );
  OAI22_X1 dp_U555 ( .A1(dp_n90), .A2(dp_n496), .B1(dp_n82), .B2(dp_n226), 
        .ZN(dp_n826) );
  INV_X1 dp_U554 ( .A(dp_rf_out1_id_o[14]), .ZN(dp_n224) );
  OAI22_X1 dp_U553 ( .A1(dp_n94), .A2(dp_n497), .B1(dp_n84), .B2(dp_n224), 
        .ZN(dp_n827) );
  INV_X1 dp_U552 ( .A(dp_rf_out1_id_o[15]), .ZN(dp_n222) );
  OAI22_X1 dp_U551 ( .A1(dp_n94), .A2(dp_n498), .B1(dp_n85), .B2(dp_n222), 
        .ZN(dp_n828) );
  INV_X1 dp_U550 ( .A(dp_rf_out1_id_o[16]), .ZN(dp_n220) );
  OAI22_X1 dp_U549 ( .A1(dp_n93), .A2(dp_n499), .B1(dp_n83), .B2(dp_n220), 
        .ZN(dp_n829) );
  INV_X1 dp_U548 ( .A(dp_rf_out1_id_o[17]), .ZN(dp_n218) );
  OAI22_X1 dp_U547 ( .A1(dp_n93), .A2(dp_n500), .B1(dp_n82), .B2(dp_n218), 
        .ZN(dp_n830) );
  INV_X1 dp_U546 ( .A(dp_rf_out1_id_o[18]), .ZN(dp_n216) );
  OAI22_X1 dp_U545 ( .A1(dp_n92), .A2(dp_n501), .B1(dp_n87), .B2(dp_n216), 
        .ZN(dp_n831) );
  INV_X1 dp_U544 ( .A(dp_rf_out1_id_o[19]), .ZN(dp_n214) );
  OAI22_X1 dp_U543 ( .A1(dp_n92), .A2(dp_n502), .B1(dp_n84), .B2(dp_n214), 
        .ZN(dp_n832) );
  INV_X1 dp_U542 ( .A(dp_rf_out1_id_o[20]), .ZN(dp_n212) );
  OAI22_X1 dp_U541 ( .A1(dp_n91), .A2(dp_n503), .B1(dp_n84), .B2(dp_n212), 
        .ZN(dp_n833) );
  INV_X1 dp_U540 ( .A(dp_rf_out1_id_o[21]), .ZN(dp_n210) );
  OAI22_X1 dp_U539 ( .A1(dp_n91), .A2(dp_n504), .B1(dp_n84), .B2(dp_n210), 
        .ZN(dp_n834) );
  INV_X1 dp_U538 ( .A(dp_rf_out1_id_o[22]), .ZN(dp_n208) );
  OAI22_X1 dp_U537 ( .A1(dp_n90), .A2(dp_n505), .B1(dp_n84), .B2(dp_n208), 
        .ZN(dp_n835) );
  INV_X1 dp_U536 ( .A(dp_rf_out1_id_o[23]), .ZN(dp_n206) );
  OAI22_X1 dp_U535 ( .A1(dp_n90), .A2(dp_n506), .B1(dp_n87), .B2(dp_n206), 
        .ZN(dp_n836) );
  INV_X1 dp_U534 ( .A(dp_rf_out1_id_o[24]), .ZN(dp_n204) );
  OAI22_X1 dp_U533 ( .A1(dp_n90), .A2(dp_n507), .B1(dp_n83), .B2(dp_n204), 
        .ZN(dp_n837) );
  INV_X1 dp_U532 ( .A(dp_npc_id_o[3]), .ZN(dp_n629) );
  OAI22_X1 dp_U531 ( .A1(dp_n98), .A2(dp_n263), .B1(dp_n81), .B2(dp_n629), 
        .ZN(dp_n720) );
  INV_X1 dp_U530 ( .A(dp_npc_id_o[4]), .ZN(dp_n630) );
  OAI22_X1 dp_U529 ( .A1(dp_n98), .A2(dp_n264), .B1(dp_n81), .B2(dp_n630), 
        .ZN(dp_n721) );
  INV_X1 dp_U528 ( .A(dp_npc_id_o[5]), .ZN(dp_n631) );
  OAI22_X1 dp_U527 ( .A1(dp_n98), .A2(dp_n265), .B1(dp_n76), .B2(dp_n631), 
        .ZN(dp_n722) );
  INV_X1 dp_U526 ( .A(dp_npc_id_o[6]), .ZN(dp_n632) );
  OAI22_X1 dp_U525 ( .A1(dp_n98), .A2(dp_n266), .B1(dp_n81), .B2(dp_n632), 
        .ZN(dp_n723) );
  INV_X1 dp_U524 ( .A(dp_npc_id_o[7]), .ZN(dp_n633) );
  OAI22_X1 dp_U523 ( .A1(dp_n98), .A2(dp_n267), .B1(dp_n80), .B2(dp_n633), 
        .ZN(dp_n724) );
  INV_X1 dp_U522 ( .A(dp_npc_id_o[8]), .ZN(dp_n634) );
  OAI22_X1 dp_U521 ( .A1(dp_n98), .A2(dp_n268), .B1(dp_n76), .B2(dp_n634), 
        .ZN(dp_n725) );
  INV_X1 dp_U520 ( .A(dp_npc_id_o[9]), .ZN(dp_n635) );
  OAI22_X1 dp_U519 ( .A1(dp_n98), .A2(dp_n269), .B1(dp_n76), .B2(dp_n635), 
        .ZN(dp_n726) );
  INV_X1 dp_U518 ( .A(dp_npc_id_o[10]), .ZN(dp_n636) );
  OAI22_X1 dp_U517 ( .A1(dp_n98), .A2(dp_n270), .B1(dp_n79), .B2(dp_n636), 
        .ZN(dp_n727) );
  INV_X1 dp_U516 ( .A(dp_npc_id_o[11]), .ZN(dp_n637) );
  OAI22_X1 dp_U515 ( .A1(dp_n98), .A2(dp_n271), .B1(dp_n81), .B2(dp_n637), 
        .ZN(dp_n728) );
  INV_X1 dp_U514 ( .A(dp_npc_id_o[12]), .ZN(dp_n638) );
  OAI22_X1 dp_U513 ( .A1(dp_n98), .A2(dp_n272), .B1(dp_n80), .B2(dp_n638), 
        .ZN(dp_n729) );
  INV_X1 dp_U512 ( .A(dp_npc_id_o[13]), .ZN(dp_n639) );
  OAI22_X1 dp_U511 ( .A1(dp_n98), .A2(dp_n273), .B1(dp_n79), .B2(dp_n639), 
        .ZN(dp_n730) );
  INV_X1 dp_U510 ( .A(dp_npc_id_o[14]), .ZN(dp_n640) );
  OAI22_X1 dp_U509 ( .A1(dp_n98), .A2(dp_n274), .B1(dp_n78), .B2(dp_n640), 
        .ZN(dp_n731) );
  INV_X1 dp_U508 ( .A(dp_npc_id_o[15]), .ZN(dp_n641) );
  OAI22_X1 dp_U507 ( .A1(dp_n98), .A2(dp_n275), .B1(dp_n80), .B2(dp_n641), 
        .ZN(dp_n732) );
  INV_X1 dp_U506 ( .A(dp_npc_id_o[16]), .ZN(dp_n642) );
  OAI22_X1 dp_U505 ( .A1(dp_n97), .A2(dp_n276), .B1(dp_n76), .B2(dp_n642), 
        .ZN(dp_n733) );
  INV_X1 dp_U504 ( .A(dp_npc_id_o[17]), .ZN(dp_n643) );
  OAI22_X1 dp_U503 ( .A1(dp_n97), .A2(dp_n277), .B1(dp_n77), .B2(dp_n643), 
        .ZN(dp_n734) );
  INV_X1 dp_U502 ( .A(dp_npc_id_o[18]), .ZN(dp_n644) );
  OAI22_X1 dp_U501 ( .A1(dp_n97), .A2(dp_n278), .B1(dp_n81), .B2(dp_n644), 
        .ZN(dp_n735) );
  INV_X1 dp_U500 ( .A(dp_npc_id_o[19]), .ZN(dp_n645) );
  OAI22_X1 dp_U499 ( .A1(dp_n97), .A2(dp_n279), .B1(dp_n81), .B2(dp_n645), 
        .ZN(dp_n736) );
  INV_X1 dp_U498 ( .A(dp_npc_id_o[20]), .ZN(dp_n646) );
  OAI22_X1 dp_U497 ( .A1(dp_n97), .A2(dp_n280), .B1(dp_n81), .B2(dp_n646), 
        .ZN(dp_n737) );
  INV_X1 dp_U496 ( .A(dp_npc_id_o[21]), .ZN(dp_n647) );
  OAI22_X1 dp_U495 ( .A1(dp_n97), .A2(dp_n281), .B1(dp_n76), .B2(dp_n647), 
        .ZN(dp_n738) );
  INV_X1 dp_U494 ( .A(dp_npc_id_o[22]), .ZN(dp_n648) );
  OAI22_X1 dp_U493 ( .A1(dp_n97), .A2(dp_n282), .B1(dp_n76), .B2(dp_n648), 
        .ZN(dp_n739) );
  INV_X1 dp_U492 ( .A(dp_npc_id_o[23]), .ZN(dp_n1016) );
  OAI22_X1 dp_U491 ( .A1(dp_n97), .A2(dp_n283), .B1(dp_n76), .B2(dp_n1016), 
        .ZN(dp_n740) );
  INV_X1 dp_U490 ( .A(dp_npc_id_o[24]), .ZN(dp_n1017) );
  OAI22_X1 dp_U489 ( .A1(dp_n97), .A2(dp_n284), .B1(dp_n81), .B2(dp_n1017), 
        .ZN(dp_n741) );
  INV_X1 dp_U488 ( .A(dp_npc_id_o[25]), .ZN(dp_n1018) );
  OAI22_X1 dp_U487 ( .A1(dp_n97), .A2(dp_n285), .B1(dp_n77), .B2(dp_n1018), 
        .ZN(dp_n742) );
  INV_X1 dp_U486 ( .A(dp_npc_id_o[26]), .ZN(dp_n1019) );
  OAI22_X1 dp_U485 ( .A1(dp_n97), .A2(dp_n286), .B1(dp_n81), .B2(dp_n1019), 
        .ZN(dp_n743) );
  INV_X1 dp_U484 ( .A(dp_npc_id_o[27]), .ZN(dp_n1020) );
  OAI22_X1 dp_U483 ( .A1(dp_n97), .A2(dp_n287), .B1(dp_n78), .B2(dp_n1020), 
        .ZN(dp_n744) );
  INV_X1 dp_U482 ( .A(dp_npc_id_o[28]), .ZN(dp_n1021) );
  OAI22_X1 dp_U481 ( .A1(dp_n97), .A2(dp_n288), .B1(dp_n79), .B2(dp_n1021), 
        .ZN(dp_n745) );
  INV_X1 dp_U480 ( .A(dp_npc_id_o[29]), .ZN(dp_n1022) );
  OAI22_X1 dp_U479 ( .A1(dp_n96), .A2(dp_n289), .B1(dp_n77), .B2(dp_n1022), 
        .ZN(dp_n746) );
  INV_X1 dp_U478 ( .A(dp_npc_id_o[30]), .ZN(dp_n1023) );
  OAI22_X1 dp_U477 ( .A1(dp_n96), .A2(dp_n290), .B1(dp_n77), .B2(dp_n1023), 
        .ZN(dp_n747) );
  INV_X1 dp_U476 ( .A(dp_npc_id_o[31]), .ZN(dp_n1024) );
  OAI22_X1 dp_U475 ( .A1(dp_n96), .A2(dp_n291), .B1(dp_n77), .B2(dp_n1024), 
        .ZN(dp_n748) );
  INV_X1 dp_U474 ( .A(dp_imm_id_o[16]), .ZN(dp_n615) );
  OAI22_X1 dp_U473 ( .A1(dp_n435), .A2(dp_n94), .B1(dp_n81), .B2(dp_n615), 
        .ZN(dp_n765) );
  INV_X1 dp_U472 ( .A(dp_imm_id_o[19]), .ZN(dp_n618) );
  OAI22_X1 dp_U471 ( .A1(dp_n438), .A2(dp_n93), .B1(dp_n79), .B2(dp_n618), 
        .ZN(dp_n768) );
  INV_X1 dp_U470 ( .A(dp_imm_id_o[20]), .ZN(dp_n619) );
  OAI22_X1 dp_U469 ( .A1(dp_n439), .A2(dp_n92), .B1(dp_n80), .B2(dp_n619), 
        .ZN(dp_n769) );
  INV_X1 dp_U468 ( .A(dp_imm_id_o[23]), .ZN(dp_n622) );
  OAI22_X1 dp_U467 ( .A1(dp_n442), .A2(dp_n94), .B1(dp_n80), .B2(dp_n622), 
        .ZN(dp_n772) );
  INV_X1 dp_U466 ( .A(dp_imm_id_o[18]), .ZN(dp_n617) );
  OAI22_X1 dp_U465 ( .A1(dp_n437), .A2(dp_n93), .B1(dp_n80), .B2(dp_n617), 
        .ZN(dp_n767) );
  INV_X1 dp_U464 ( .A(dp_imm_id_o[21]), .ZN(dp_n620) );
  OAI22_X1 dp_U463 ( .A1(dp_n440), .A2(dp_n92), .B1(dp_n79), .B2(dp_n620), 
        .ZN(dp_n770) );
  INV_X1 dp_U462 ( .A(dp_imm_id_o[24]), .ZN(dp_n623) );
  OAI22_X1 dp_U461 ( .A1(dp_n443), .A2(dp_n92), .B1(dp_n81), .B2(dp_n623), 
        .ZN(dp_n773) );
  INV_X1 dp_U460 ( .A(dp_imm_id_o[17]), .ZN(dp_n616) );
  OAI22_X1 dp_U459 ( .A1(dp_n436), .A2(dp_n90), .B1(dp_n80), .B2(dp_n616), 
        .ZN(dp_n766) );
  INV_X1 dp_U458 ( .A(dp_rf_out1_id_o[31]), .ZN(dp_n190) );
  OAI22_X1 dp_U457 ( .A1(dp_n94), .A2(dp_n514), .B1(dp_n85), .B2(dp_n190), 
        .ZN(dp_n844) );
  INV_X1 dp_U456 ( .A(dp_rf_out1_id_o[26]), .ZN(dp_n200) );
  OAI22_X1 dp_U455 ( .A1(dp_n92), .A2(dp_n509), .B1(dp_n82), .B2(dp_n200), 
        .ZN(dp_n839) );
  INV_X1 dp_U454 ( .A(dp_rf_out1_id_o[29]), .ZN(dp_n194) );
  OAI22_X1 dp_U453 ( .A1(dp_n91), .A2(dp_n512), .B1(dp_n85), .B2(dp_n194), 
        .ZN(dp_n842) );
  INV_X1 dp_U452 ( .A(dp_rf_out1_id_o[25]), .ZN(dp_n202) );
  OAI22_X1 dp_U451 ( .A1(dp_n94), .A2(dp_n508), .B1(dp_n85), .B2(dp_n202), 
        .ZN(dp_n838) );
  INV_X1 dp_U450 ( .A(dp_rf_out1_id_o[27]), .ZN(dp_n198) );
  OAI22_X1 dp_U449 ( .A1(dp_n92), .A2(dp_n510), .B1(dp_n84), .B2(dp_n198), 
        .ZN(dp_n840) );
  INV_X1 dp_U448 ( .A(dp_rf_out1_id_o[28]), .ZN(dp_n196) );
  OAI22_X1 dp_U447 ( .A1(dp_n93), .A2(dp_n511), .B1(dp_n87), .B2(dp_n196), 
        .ZN(dp_n841) );
  INV_X1 dp_U446 ( .A(dp_rf_out1_id_o[30]), .ZN(dp_n192) );
  OAI22_X1 dp_U445 ( .A1(dp_n91), .A2(dp_n513), .B1(dp_n84), .B2(dp_n192), 
        .ZN(dp_n843) );
  INV_X1 dp_U444 ( .A(dp_rf_out2_id_o[0]), .ZN(dp_n251) );
  OAI22_X1 dp_U443 ( .A1(dp_n96), .A2(dp_n451), .B1(dp_n77), .B2(dp_n251), 
        .ZN(dp_n781) );
  INV_X1 dp_U442 ( .A(dp_rf_out2_id_o[1]), .ZN(dp_n249) );
  OAI22_X1 dp_U441 ( .A1(dp_n96), .A2(dp_n452), .B1(dp_n78), .B2(dp_n249), 
        .ZN(dp_n782) );
  INV_X1 dp_U440 ( .A(dp_rf_out2_id_o[2]), .ZN(dp_n247) );
  OAI22_X1 dp_U439 ( .A1(dp_n96), .A2(dp_n453), .B1(dp_n78), .B2(dp_n247), 
        .ZN(dp_n783) );
  INV_X1 dp_U438 ( .A(dp_imm_id_o[14]), .ZN(dp_n612) );
  OAI22_X1 dp_U437 ( .A1(dp_n433), .A2(dp_n91), .B1(dp_n78), .B2(dp_n612), 
        .ZN(dp_n763) );
  INV_X1 dp_U436 ( .A(dp_imm_id_o[1]), .ZN(dp_n595) );
  OAI22_X1 dp_U435 ( .A1(dp_n420), .A2(dp_n93), .B1(dp_n79), .B2(dp_n595), 
        .ZN(dp_n750) );
  INV_X1 dp_U434 ( .A(dp_imm_id_o[2]), .ZN(dp_n596) );
  OAI22_X1 dp_U433 ( .A1(dp_n421), .A2(dp_n92), .B1(dp_n80), .B2(dp_n596), 
        .ZN(dp_n751) );
  INV_X1 dp_U432 ( .A(dp_imm_id_o[4]), .ZN(dp_n598) );
  OAI22_X1 dp_U431 ( .A1(dp_n423), .A2(dp_n91), .B1(dp_n76), .B2(dp_n598), 
        .ZN(dp_n753) );
  INV_X1 dp_U430 ( .A(dp_imm_id_o[5]), .ZN(dp_n599) );
  OAI22_X1 dp_U429 ( .A1(dp_n424), .A2(dp_n90), .B1(dp_n76), .B2(dp_n599), 
        .ZN(dp_n754) );
  INV_X1 dp_U428 ( .A(dp_imm_id_o[7]), .ZN(dp_n601) );
  OAI22_X1 dp_U427 ( .A1(dp_n426), .A2(dp_n94), .B1(dp_n77), .B2(dp_n601), 
        .ZN(dp_n756) );
  INV_X1 dp_U426 ( .A(dp_imm_id_o[11]), .ZN(dp_n606) );
  OAI22_X1 dp_U425 ( .A1(dp_n430), .A2(dp_n91), .B1(dp_n81), .B2(dp_n606), 
        .ZN(dp_n760) );
  INV_X1 dp_U424 ( .A(dp_imm_id_o[0]), .ZN(dp_n594) );
  OAI22_X1 dp_U423 ( .A1(dp_n419), .A2(dp_n90), .B1(dp_n81), .B2(dp_n594), 
        .ZN(dp_n749) );
  INV_X1 dp_U422 ( .A(dp_imm_id_o[3]), .ZN(dp_n597) );
  OAI22_X1 dp_U421 ( .A1(dp_n422), .A2(dp_n93), .B1(dp_n79), .B2(dp_n597), 
        .ZN(dp_n752) );
  INV_X1 dp_U420 ( .A(dp_imm_id_o[6]), .ZN(dp_n600) );
  OAI22_X1 dp_U419 ( .A1(dp_n425), .A2(dp_n92), .B1(dp_n77), .B2(dp_n600), 
        .ZN(dp_n755) );
  INV_X1 dp_U418 ( .A(dp_imm_id_o[8]), .ZN(dp_n602) );
  OAI22_X1 dp_U417 ( .A1(dp_n427), .A2(dp_n91), .B1(dp_n79), .B2(dp_n602), 
        .ZN(dp_n757) );
  INV_X1 dp_U416 ( .A(dp_imm_id_o[9]), .ZN(dp_n603) );
  OAI22_X1 dp_U415 ( .A1(dp_n428), .A2(dp_n94), .B1(dp_n81), .B2(dp_n603), 
        .ZN(dp_n758) );
  INV_X1 dp_U414 ( .A(dp_imm_id_o[10]), .ZN(dp_n604) );
  OAI22_X1 dp_U413 ( .A1(dp_n429), .A2(dp_n90), .B1(dp_n79), .B2(dp_n604), 
        .ZN(dp_n759) );
  INV_X1 dp_U412 ( .A(dp_imm_id_o[12]), .ZN(dp_n608) );
  OAI22_X1 dp_U411 ( .A1(dp_n431), .A2(dp_n90), .B1(dp_n78), .B2(dp_n608), 
        .ZN(dp_n761) );
  INV_X1 dp_U410 ( .A(dp_imm_id_o[13]), .ZN(dp_n610) );
  OAI22_X1 dp_U409 ( .A1(dp_n432), .A2(dp_n90), .B1(dp_n78), .B2(dp_n610), 
        .ZN(dp_n762) );
  INV_X1 dp_U408 ( .A(dp_imm_id_o[15]), .ZN(dp_n614) );
  OAI22_X1 dp_U407 ( .A1(dp_n434), .A2(dp_n94), .B1(dp_n77), .B2(dp_n614), 
        .ZN(dp_n764) );
  OAI22_X1 dp_U406 ( .A1(dp_n332), .A2(dp_n63), .B1(dp_n876), .B2(dp_n57), 
        .ZN(dp_n908) );
  OAI22_X1 dp_U405 ( .A1(dp_n333), .A2(dp_n64), .B1(dp_n875), .B2(dp_n57), 
        .ZN(dp_n907) );
  OAI22_X1 dp_U404 ( .A1(dp_n334), .A2(dp_n64), .B1(dp_n874), .B2(dp_n57), 
        .ZN(dp_n906) );
  OAI22_X1 dp_U403 ( .A1(dp_n402), .A2(dp_n64), .B1(dp_n873), .B2(dp_n57), 
        .ZN(dp_n905) );
  OAI22_X1 dp_U402 ( .A1(dp_n403), .A2(dp_n64), .B1(dp_n872), .B2(dp_n57), 
        .ZN(dp_n904) );
  OAI22_X1 dp_U401 ( .A1(dp_n404), .A2(dp_n64), .B1(dp_n871), .B2(dp_n57), 
        .ZN(dp_n903) );
  OAI22_X1 dp_U400 ( .A1(dp_n405), .A2(dp_n64), .B1(dp_n870), .B2(dp_n57), 
        .ZN(dp_n902) );
  OAI22_X1 dp_U399 ( .A1(dp_n406), .A2(dp_n64), .B1(dp_n869), .B2(dp_n56), 
        .ZN(dp_n901) );
  OAI22_X1 dp_U398 ( .A1(dp_n407), .A2(dp_n64), .B1(dp_n868), .B2(dp_n56), 
        .ZN(dp_n900) );
  OAI22_X1 dp_U397 ( .A1(dp_n408), .A2(dp_n64), .B1(dp_n867), .B2(dp_n56), 
        .ZN(dp_n899) );
  OAI22_X1 dp_U396 ( .A1(dp_n409), .A2(dp_n64), .B1(dp_n866), .B2(dp_n56), 
        .ZN(dp_n898) );
  OAI22_X1 dp_U395 ( .A1(dp_n410), .A2(dp_n64), .B1(dp_n865), .B2(dp_n56), 
        .ZN(dp_n897) );
  OAI22_X1 dp_U394 ( .A1(dp_n411), .A2(dp_n64), .B1(dp_n864), .B2(dp_n56), 
        .ZN(dp_n896) );
  OAI22_X1 dp_U393 ( .A1(dp_n412), .A2(dp_n65), .B1(dp_n863), .B2(dp_n56), 
        .ZN(dp_n895) );
  OAI22_X1 dp_U392 ( .A1(dp_n413), .A2(dp_n65), .B1(dp_n862), .B2(dp_n56), 
        .ZN(dp_n894) );
  OAI22_X1 dp_U391 ( .A1(dp_n517), .A2(dp_n65), .B1(dp_n861), .B2(dp_n56), 
        .ZN(dp_n893) );
  OAI22_X1 dp_U390 ( .A1(dp_n519), .A2(dp_n65), .B1(dp_n860), .B2(dp_n56), 
        .ZN(dp_n892) );
  OAI22_X1 dp_U389 ( .A1(dp_n521), .A2(dp_n65), .B1(dp_n859), .B2(dp_n56), 
        .ZN(dp_n891) );
  OAI22_X1 dp_U388 ( .A1(dp_n523), .A2(dp_n65), .B1(dp_n858), .B2(dp_n56), 
        .ZN(dp_n890) );
  INV_X1 dp_U387 ( .A(reg31_sel_i), .ZN(dp_n1026) );
  INV_X1 dp_U386 ( .A(regrd_sel_i), .ZN(dp_n1028) );
  INV_X1 dp_U385 ( .A(dp_npc_if_o[10]), .ZN(dp_n148) );
  OAI22_X1 dp_U384 ( .A1(dp_n110), .A2(dp_n552), .B1(dp_n102), .B2(dp_n148), 
        .ZN(dp_n685) );
  INV_X1 dp_U383 ( .A(dp_npc_if_o[11]), .ZN(dp_n147) );
  OAI22_X1 dp_U382 ( .A1(dp_n109), .A2(dp_n553), .B1(dp_n4), .B2(dp_n147), 
        .ZN(dp_n686) );
  INV_X1 dp_U381 ( .A(dp_npc_if_o[12]), .ZN(dp_n146) );
  OAI22_X1 dp_U380 ( .A1(dp_n109), .A2(dp_n554), .B1(dp_n101), .B2(dp_n146), 
        .ZN(dp_n687) );
  INV_X1 dp_U379 ( .A(dp_npc_if_o[13]), .ZN(dp_n145) );
  OAI22_X1 dp_U378 ( .A1(dp_n109), .A2(dp_n555), .B1(dp_n4), .B2(dp_n145), 
        .ZN(dp_n688) );
  INV_X1 dp_U377 ( .A(dp_npc_if_o[14]), .ZN(dp_n144) );
  OAI22_X1 dp_U376 ( .A1(dp_n109), .A2(dp_n556), .B1(dp_n100), .B2(dp_n144), 
        .ZN(dp_n689) );
  INV_X1 dp_U375 ( .A(dp_npc_if_o[15]), .ZN(dp_n143) );
  OAI22_X1 dp_U374 ( .A1(dp_n110), .A2(dp_n557), .B1(dp_n102), .B2(dp_n143), 
        .ZN(dp_n690) );
  INV_X1 dp_U373 ( .A(dp_npc_if_o[0]), .ZN(dp_n253) );
  OAI22_X1 dp_U372 ( .A1(dp_n109), .A2(dp_n542), .B1(dp_n4), .B2(dp_n253), 
        .ZN(dp_n675) );
  INV_X1 dp_U371 ( .A(dp_npc_if_o[1]), .ZN(dp_n157) );
  OAI22_X1 dp_U370 ( .A1(dp_n110), .A2(dp_n543), .B1(dp_n3), .B2(dp_n157), 
        .ZN(dp_n676) );
  INV_X1 dp_U369 ( .A(dp_npc_if_o[2]), .ZN(dp_n156) );
  OAI22_X1 dp_U368 ( .A1(dp_n109), .A2(dp_n544), .B1(dp_n4), .B2(dp_n156), 
        .ZN(dp_n677) );
  INV_X1 dp_U367 ( .A(dp_npc_if_o[3]), .ZN(dp_n155) );
  OAI22_X1 dp_U366 ( .A1(dp_n109), .A2(dp_n545), .B1(dp_n101), .B2(dp_n155), 
        .ZN(dp_n678) );
  INV_X1 dp_U365 ( .A(dp_npc_if_o[4]), .ZN(dp_n154) );
  OAI22_X1 dp_U364 ( .A1(dp_n110), .A2(dp_n546), .B1(dp_n101), .B2(dp_n154), 
        .ZN(dp_n679) );
  INV_X1 dp_U363 ( .A(dp_npc_if_o[5]), .ZN(dp_n153) );
  OAI22_X1 dp_U362 ( .A1(dp_n109), .A2(dp_n547), .B1(dp_n100), .B2(dp_n153), 
        .ZN(dp_n680) );
  INV_X1 dp_U361 ( .A(dp_npc_if_o[6]), .ZN(dp_n152) );
  OAI22_X1 dp_U360 ( .A1(dp_n110), .A2(dp_n548), .B1(dp_n101), .B2(dp_n152), 
        .ZN(dp_n681) );
  INV_X1 dp_U359 ( .A(dp_npc_if_o[7]), .ZN(dp_n151) );
  OAI22_X1 dp_U358 ( .A1(dp_n109), .A2(dp_n549), .B1(dp_n3), .B2(dp_n151), 
        .ZN(dp_n682) );
  INV_X1 dp_U357 ( .A(dp_npc_if_o[8]), .ZN(dp_n150) );
  OAI22_X1 dp_U356 ( .A1(dp_n109), .A2(dp_n550), .B1(dp_n3), .B2(dp_n150), 
        .ZN(dp_n683) );
  INV_X1 dp_U355 ( .A(dp_npc_if_o[9]), .ZN(dp_n149) );
  OAI22_X1 dp_U354 ( .A1(dp_n109), .A2(dp_n551), .B1(dp_n3), .B2(dp_n149), 
        .ZN(dp_n684) );
  INV_X1 dp_U353 ( .A(IRAM_DATA[0]), .ZN(dp_n1055) );
  OAI22_X1 dp_U352 ( .A1(dp_n526), .A2(dp_n107), .B1(dp_n100), .B2(dp_n1055), 
        .ZN(dp_n649) );
  INV_X1 dp_U351 ( .A(IRAM_DATA[1]), .ZN(dp_n1054) );
  OAI22_X1 dp_U350 ( .A1(dp_n527), .A2(dp_n107), .B1(dp_n101), .B2(dp_n1054), 
        .ZN(dp_n650) );
  INV_X1 dp_U349 ( .A(IRAM_DATA[2]), .ZN(dp_n1053) );
  OAI22_X1 dp_U348 ( .A1(dp_n528), .A2(dp_n107), .B1(dp_n69), .B2(dp_n1053), 
        .ZN(dp_n651) );
  INV_X1 dp_U347 ( .A(IRAM_DATA[3]), .ZN(dp_n1052) );
  OAI22_X1 dp_U346 ( .A1(dp_n529), .A2(dp_n108), .B1(dp_n3), .B2(dp_n1052), 
        .ZN(dp_n652) );
  INV_X1 dp_U345 ( .A(IRAM_DATA[4]), .ZN(dp_n1051) );
  OAI22_X1 dp_U344 ( .A1(dp_n530), .A2(dp_n108), .B1(dp_n4), .B2(dp_n1051), 
        .ZN(dp_n653) );
  INV_X1 dp_U343 ( .A(IRAM_DATA[5]), .ZN(dp_n1050) );
  OAI22_X1 dp_U342 ( .A1(dp_n531), .A2(dp_n107), .B1(dp_n3), .B2(dp_n1050), 
        .ZN(dp_n654) );
  INV_X1 dp_U341 ( .A(IRAM_DATA[6]), .ZN(dp_n1049) );
  OAI22_X1 dp_U340 ( .A1(dp_n532), .A2(dp_n108), .B1(dp_n100), .B2(dp_n1049), 
        .ZN(dp_n655) );
  INV_X1 dp_U339 ( .A(IRAM_DATA[7]), .ZN(dp_n1048) );
  OAI22_X1 dp_U338 ( .A1(dp_n533), .A2(dp_n107), .B1(dp_n100), .B2(dp_n1048), 
        .ZN(dp_n656) );
  INV_X1 dp_U337 ( .A(IRAM_DATA[8]), .ZN(dp_n1047) );
  OAI22_X1 dp_U336 ( .A1(dp_n534), .A2(dp_n107), .B1(dp_n102), .B2(dp_n1047), 
        .ZN(dp_n657) );
  INV_X1 dp_U335 ( .A(IRAM_DATA[9]), .ZN(dp_n1046) );
  OAI22_X1 dp_U334 ( .A1(dp_n535), .A2(dp_n108), .B1(dp_n4), .B2(dp_n1046), 
        .ZN(dp_n658) );
  INV_X1 dp_U333 ( .A(IRAM_DATA[10]), .ZN(dp_n1045) );
  OAI22_X1 dp_U332 ( .A1(dp_n536), .A2(dp_n108), .B1(dp_n69), .B2(dp_n1045), 
        .ZN(dp_n659) );
  INV_X1 dp_U331 ( .A(IRAM_DATA[11]), .ZN(dp_n1044) );
  OAI22_X1 dp_U330 ( .A1(dp_n575), .A2(dp_n107), .B1(dp_n100), .B2(dp_n1044), 
        .ZN(dp_n660) );
  INV_X1 dp_U329 ( .A(IRAM_DATA[12]), .ZN(dp_n1043) );
  OAI22_X1 dp_U328 ( .A1(dp_n577), .A2(dp_n108), .B1(dp_n4), .B2(dp_n1043), 
        .ZN(dp_n661) );
  INV_X1 dp_U327 ( .A(IRAM_DATA[13]), .ZN(dp_n1042) );
  OAI22_X1 dp_U326 ( .A1(dp_n579), .A2(dp_n108), .B1(dp_n100), .B2(dp_n1042), 
        .ZN(dp_n662) );
  INV_X1 dp_U325 ( .A(IRAM_DATA[14]), .ZN(dp_n1041) );
  OAI22_X1 dp_U324 ( .A1(dp_n581), .A2(dp_n107), .B1(dp_n101), .B2(dp_n1041), 
        .ZN(dp_n663) );
  INV_X1 dp_U323 ( .A(IRAM_DATA[15]), .ZN(dp_n1040) );
  OAI22_X1 dp_U322 ( .A1(dp_n583), .A2(dp_n107), .B1(dp_n69), .B2(dp_n1040), 
        .ZN(dp_n664) );
  INV_X1 dp_U321 ( .A(IRAM_DATA[16]), .ZN(dp_n1039) );
  OAI22_X1 dp_U320 ( .A1(dp_n574), .A2(dp_n108), .B1(dp_n102), .B2(dp_n1039), 
        .ZN(dp_n665) );
  INV_X1 dp_U319 ( .A(IRAM_DATA[17]), .ZN(dp_n1038) );
  OAI22_X1 dp_U318 ( .A1(dp_n576), .A2(dp_n108), .B1(dp_n102), .B2(dp_n1038), 
        .ZN(dp_n666) );
  INV_X1 dp_U317 ( .A(IRAM_DATA[18]), .ZN(dp_n1037) );
  OAI22_X1 dp_U316 ( .A1(dp_n578), .A2(dp_n108), .B1(dp_n101), .B2(dp_n1037), 
        .ZN(dp_n667) );
  INV_X1 dp_U315 ( .A(IRAM_DATA[19]), .ZN(dp_n1036) );
  OAI22_X1 dp_U314 ( .A1(dp_n580), .A2(dp_n108), .B1(dp_n69), .B2(dp_n1036), 
        .ZN(dp_n668) );
  INV_X1 dp_U313 ( .A(IRAM_DATA[20]), .ZN(dp_n1035) );
  OAI22_X1 dp_U312 ( .A1(dp_n582), .A2(dp_n108), .B1(dp_n102), .B2(dp_n1035), 
        .ZN(dp_n669) );
  INV_X1 dp_U311 ( .A(IRAM_DATA[23]), .ZN(dp_n1032) );
  OAI22_X1 dp_U310 ( .A1(dp_n539), .A2(dp_n107), .B1(dp_n3), .B2(dp_n1032), 
        .ZN(dp_n672) );
  INV_X1 dp_U309 ( .A(IRAM_DATA[24]), .ZN(dp_n1031) );
  OAI22_X1 dp_U308 ( .A1(dp_n540), .A2(dp_n107), .B1(dp_n69), .B2(dp_n1031), 
        .ZN(dp_n673) );
  INV_X1 dp_U307 ( .A(IRAM_DATA[25]), .ZN(dp_n1030) );
  OAI22_X1 dp_U306 ( .A1(dp_n541), .A2(dp_n107), .B1(dp_n102), .B2(dp_n1030), 
        .ZN(dp_n674) );
  INV_X1 dp_U305 ( .A(IRAM_DATA[21]), .ZN(dp_n1034) );
  OAI22_X1 dp_U304 ( .A1(dp_n537), .A2(dp_n109), .B1(dp_n101), .B2(dp_n1034), 
        .ZN(dp_n670) );
  INV_X1 dp_U303 ( .A(IRAM_DATA[22]), .ZN(dp_n1033) );
  OAI22_X1 dp_U302 ( .A1(dp_n538), .A2(dp_n109), .B1(dp_n3), .B2(dp_n1033), 
        .ZN(dp_n671) );
  INV_X1 dp_U301 ( .A(dp_alu_out_ex_o[7]), .ZN(dp_n182) );
  OAI22_X1 dp_U300 ( .A1(dp_n870), .A2(dp_n73), .B1(dp_n67), .B2(dp_n182), 
        .ZN(dp_n934) );
  INV_X1 dp_U299 ( .A(dp_alu_out_ex_o[18]), .ZN(dp_n171) );
  OAI22_X1 dp_U298 ( .A1(dp_n859), .A2(dp_n72), .B1(dp_n67), .B2(dp_n171), 
        .ZN(dp_n923) );
  INV_X1 dp_U297 ( .A(dp_alu_out_ex_o[13]), .ZN(dp_n176) );
  OAI22_X1 dp_U296 ( .A1(dp_n864), .A2(dp_n72), .B1(dp_n67), .B2(dp_n176), 
        .ZN(dp_n928) );
  INV_X1 dp_U295 ( .A(dp_alu_out_ex_o[14]), .ZN(dp_n175) );
  OAI22_X1 dp_U294 ( .A1(dp_n863), .A2(dp_n72), .B1(dp_n67), .B2(dp_n175), 
        .ZN(dp_n927) );
  INV_X1 dp_U293 ( .A(dp_alu_out_ex_o[15]), .ZN(dp_n174) );
  OAI22_X1 dp_U292 ( .A1(dp_n862), .A2(dp_n72), .B1(dp_n67), .B2(dp_n174), 
        .ZN(dp_n926) );
  INV_X1 dp_U291 ( .A(dp_alu_out_ex_o[9]), .ZN(dp_n180) );
  OAI22_X1 dp_U290 ( .A1(dp_n868), .A2(dp_n72), .B1(dp_n67), .B2(dp_n180), 
        .ZN(dp_n932) );
  INV_X1 dp_U289 ( .A(dp_alu_out_ex_o[8]), .ZN(dp_n181) );
  OAI22_X1 dp_U288 ( .A1(dp_n869), .A2(dp_n73), .B1(dp_n67), .B2(dp_n181), 
        .ZN(dp_n933) );
  INV_X1 dp_U287 ( .A(dp_alu_out_ex_o[10]), .ZN(dp_n179) );
  OAI22_X1 dp_U286 ( .A1(dp_n867), .A2(dp_n72), .B1(dp_n67), .B2(dp_n179), 
        .ZN(dp_n931) );
  INV_X1 dp_U285 ( .A(dp_alu_out_ex_o[17]), .ZN(dp_n172) );
  OAI22_X1 dp_U284 ( .A1(dp_n860), .A2(dp_n72), .B1(dp_n172), .B2(dp_n67), 
        .ZN(dp_n924) );
  INV_X1 dp_U283 ( .A(dp_alu_out_ex_o[11]), .ZN(dp_n178) );
  OAI22_X1 dp_U282 ( .A1(dp_n866), .A2(dp_n72), .B1(dp_n67), .B2(dp_n178), 
        .ZN(dp_n930) );
  INV_X1 dp_U281 ( .A(dp_alu_out_ex_o[12]), .ZN(dp_n177) );
  OAI22_X1 dp_U280 ( .A1(dp_n865), .A2(dp_n72), .B1(dp_n67), .B2(dp_n177), 
        .ZN(dp_n929) );
  INV_X1 dp_U279 ( .A(dp_alu_out_ex_o[16]), .ZN(dp_n173) );
  OAI22_X1 dp_U278 ( .A1(dp_n861), .A2(dp_n72), .B1(dp_n173), .B2(dp_n67), 
        .ZN(dp_n925) );
  INV_X1 dp_U277 ( .A(dp_rd_fwd_ex_o[0]), .ZN(dp_n255) );
  OAI22_X1 dp_U276 ( .A1(dp_n71), .A2(dp_n293), .B1(dp_n67), .B2(dp_n255), 
        .ZN(dp_n1014) );
  OAI22_X1 dp_U275 ( .A1(dp_n872), .A2(dp_n73), .B1(dp_n67), .B2(dp_n184), 
        .ZN(dp_n936) );
  INV_X1 dp_U274 ( .A(dp_alu_out_ex_o[3]), .ZN(dp_n186) );
  OAI22_X1 dp_U273 ( .A1(dp_n874), .A2(dp_n73), .B1(dp_n67), .B2(dp_n186), 
        .ZN(dp_n938) );
  INV_X1 dp_U272 ( .A(dp_alu_out_ex_o[2]), .ZN(dp_n187) );
  OAI22_X1 dp_U271 ( .A1(dp_n875), .A2(dp_n73), .B1(dp_n67), .B2(dp_n187), 
        .ZN(dp_n939) );
  INV_X1 dp_U270 ( .A(dp_branch_t_ex_o), .ZN(dp_n292) );
  OAI22_X1 dp_U269 ( .A1(dp_n515), .A2(dp_n71), .B1(dp_n67), .B2(dp_n292), 
        .ZN(dp_n845) );
  INV_X1 dp_U268 ( .A(dp_rd_fwd_ex_o[1]), .ZN(dp_n256) );
  OAI22_X1 dp_U267 ( .A1(dp_n73), .A2(dp_n294), .B1(dp_n67), .B2(dp_n256), 
        .ZN(dp_n1013) );
  INV_X1 dp_U266 ( .A(dp_rd_fwd_ex_o[2]), .ZN(dp_n257) );
  OAI22_X1 dp_U265 ( .A1(dp_n73), .A2(dp_n295), .B1(dp_n67), .B2(dp_n257), 
        .ZN(dp_n1012) );
  INV_X1 dp_U264 ( .A(dp_rd_fwd_ex_o[3]), .ZN(dp_n258) );
  OAI22_X1 dp_U263 ( .A1(dp_n73), .A2(dp_n296), .B1(dp_n67), .B2(dp_n258), 
        .ZN(dp_n1011) );
  INV_X1 dp_U262 ( .A(dp_rd_fwd_ex_o[4]), .ZN(dp_n259) );
  OAI22_X1 dp_U261 ( .A1(dp_n73), .A2(dp_n297), .B1(dp_n67), .B2(dp_n259), 
        .ZN(dp_n1010) );
  OAI22_X1 dp_U260 ( .A1(dp_n873), .A2(dp_n73), .B1(dp_n67), .B2(dp_n185), 
        .ZN(dp_n937) );
  INV_X1 dp_U259 ( .A(dp_alu_out_ex_o[1]), .ZN(dp_n188) );
  OAI22_X1 dp_U258 ( .A1(dp_n876), .A2(dp_n73), .B1(dp_n67), .B2(dp_n188), 
        .ZN(dp_n940) );
  INV_X1 dp_U257 ( .A(dp_alu_out_ex_o[6]), .ZN(dp_n183) );
  OAI22_X1 dp_U256 ( .A1(dp_n871), .A2(dp_n73), .B1(dp_n67), .B2(dp_n183), 
        .ZN(dp_n935) );
  OAI221_X1 dp_U255 ( .B1(dp_n577), .B2(regrd_sel_i), .C1(dp_n576), .C2(
        dp_n1028), .A(dp_n1026), .ZN(dp_rd_fwd_id_o[1]) );
  INV_X1 dp_U254 ( .A(dp_rd_fwd_id_o[1]), .ZN(dp_n607) );
  OAI22_X1 dp_U253 ( .A1(dp_n99), .A2(dp_n415), .B1(dp_n77), .B2(dp_n607), 
        .ZN(dp_n713) );
  OAI221_X1 dp_U252 ( .B1(dp_n579), .B2(regrd_sel_i), .C1(dp_n578), .C2(
        dp_n1028), .A(dp_n1026), .ZN(dp_rd_fwd_id_o[2]) );
  INV_X1 dp_U251 ( .A(dp_rd_fwd_id_o[2]), .ZN(dp_n609) );
  OAI22_X1 dp_U250 ( .A1(dp_n99), .A2(dp_n416), .B1(dp_n80), .B2(dp_n609), 
        .ZN(dp_n714) );
  OAI221_X1 dp_U249 ( .B1(dp_n581), .B2(regrd_sel_i), .C1(dp_n580), .C2(
        dp_n1028), .A(dp_n1026), .ZN(dp_rd_fwd_id_o[3]) );
  INV_X1 dp_U248 ( .A(dp_rd_fwd_id_o[3]), .ZN(dp_n611) );
  OAI22_X1 dp_U247 ( .A1(dp_n99), .A2(dp_n417), .B1(dp_n76), .B2(dp_n611), 
        .ZN(dp_n715) );
  OAI221_X1 dp_U246 ( .B1(dp_n583), .B2(regrd_sel_i), .C1(dp_n582), .C2(
        dp_n1028), .A(dp_n1026), .ZN(dp_rd_fwd_id_o[4]) );
  INV_X1 dp_U245 ( .A(dp_rd_fwd_id_o[4]), .ZN(dp_n613) );
  OAI22_X1 dp_U244 ( .A1(dp_n99), .A2(dp_n418), .B1(dp_n78), .B2(dp_n613), 
        .ZN(dp_n716) );
  INV_X1 dp_U243 ( .A(dp_npc_id_o[0]), .ZN(dp_n626) );
  OAI22_X1 dp_U242 ( .A1(dp_n99), .A2(dp_n260), .B1(dp_n77), .B2(dp_n626), 
        .ZN(dp_n717) );
  INV_X1 dp_U241 ( .A(dp_npc_id_o[1]), .ZN(dp_n627) );
  OAI22_X1 dp_U240 ( .A1(dp_n99), .A2(dp_n261), .B1(dp_n78), .B2(dp_n627), 
        .ZN(dp_n718) );
  INV_X1 dp_U239 ( .A(dp_npc_id_o[2]), .ZN(dp_n628) );
  OAI22_X1 dp_U238 ( .A1(dp_n99), .A2(dp_n262), .B1(dp_n78), .B2(dp_n628), 
        .ZN(dp_n719) );
  AOI22_X1 dp_U237 ( .A1(dp_data_mem_ex_o[8]), .A2(dp_n51), .B1(dp_z_word[8]), 
        .B2(dp_n47), .ZN(dp_n392) );
  OAI221_X1 dp_U236 ( .B1(dp_n268), .B2(dp_n53), .C1(dp_n72), .C2(dp_n358), 
        .A(dp_n392), .ZN(dp_n996) );
  AOI22_X1 dp_U235 ( .A1(dp_data_mem_ex_o[9]), .A2(dp_n50), .B1(dp_z_word[9]), 
        .B2(dp_n47), .ZN(dp_n391) );
  OAI221_X1 dp_U234 ( .B1(dp_n269), .B2(dp_n53), .C1(dp_n73), .C2(dp_n357), 
        .A(dp_n391), .ZN(dp_n995) );
  AOI22_X1 dp_U233 ( .A1(dp_data_mem_ex_o[10]), .A2(dp_n50), .B1(dp_z_word[10]), .B2(dp_n47), .ZN(dp_n390) );
  OAI221_X1 dp_U232 ( .B1(dp_n270), .B2(dp_n53), .C1(dp_n71), .C2(dp_n356), 
        .A(dp_n390), .ZN(dp_n994) );
  AOI22_X1 dp_U231 ( .A1(dp_data_mem_ex_o[11]), .A2(dp_n49), .B1(dp_z_word[11]), .B2(dp_n47), .ZN(dp_n389) );
  OAI221_X1 dp_U230 ( .B1(dp_n271), .B2(dp_n53), .C1(dp_n72), .C2(dp_n355), 
        .A(dp_n389), .ZN(dp_n993) );
  AOI22_X1 dp_U229 ( .A1(dp_data_mem_ex_o[12]), .A2(dp_n51), .B1(dp_z_word[12]), .B2(dp_n47), .ZN(dp_n388) );
  OAI221_X1 dp_U228 ( .B1(dp_n272), .B2(dp_n53), .C1(dp_n73), .C2(dp_n354), 
        .A(dp_n388), .ZN(dp_n992) );
  AOI22_X1 dp_U227 ( .A1(dp_data_mem_ex_o[13]), .A2(dp_n49), .B1(dp_z_word[13]), .B2(dp_n47), .ZN(dp_n387) );
  OAI221_X1 dp_U226 ( .B1(dp_n273), .B2(dp_n53), .C1(dp_n73), .C2(dp_n353), 
        .A(dp_n387), .ZN(dp_n991) );
  AOI22_X1 dp_U225 ( .A1(dp_data_mem_ex_o[14]), .A2(dp_n51), .B1(dp_z_word[14]), .B2(dp_n47), .ZN(dp_n386) );
  OAI221_X1 dp_U224 ( .B1(dp_n274), .B2(dp_n53), .C1(dp_n73), .C2(dp_n352), 
        .A(dp_n386), .ZN(dp_n990) );
  AOI22_X1 dp_U223 ( .A1(dp_data_mem_ex_o[15]), .A2(dp_n49), .B1(dp_z_word[15]), .B2(dp_n47), .ZN(dp_n385) );
  OAI221_X1 dp_U222 ( .B1(dp_n275), .B2(dp_n53), .C1(dp_n71), .C2(dp_n351), 
        .A(dp_n385), .ZN(dp_n989) );
  AOI22_X1 dp_U221 ( .A1(dp_data_mem_ex_o[16]), .A2(dp_n51), .B1(dp_z_word[16]), .B2(dp_n47), .ZN(dp_n384) );
  OAI221_X1 dp_U220 ( .B1(dp_n276), .B2(dp_n53), .C1(dp_n72), .C2(dp_n350), 
        .A(dp_n384), .ZN(dp_n988) );
  AOI22_X1 dp_U219 ( .A1(dp_data_mem_ex_o[17]), .A2(dp_n49), .B1(dp_z_word[17]), .B2(dp_n47), .ZN(dp_n383) );
  OAI221_X1 dp_U218 ( .B1(dp_n277), .B2(dp_n53), .C1(dp_n71), .C2(dp_n349), 
        .A(dp_n383), .ZN(dp_n987) );
  AOI22_X1 dp_U217 ( .A1(dp_data_mem_ex_o[18]), .A2(dp_n51), .B1(dp_z_word[18]), .B2(dp_n47), .ZN(dp_n382) );
  OAI221_X1 dp_U216 ( .B1(dp_n278), .B2(dp_n53), .C1(dp_n73), .C2(dp_n348), 
        .A(dp_n382), .ZN(dp_n986) );
  AOI22_X1 dp_U215 ( .A1(dp_data_mem_ex_o[19]), .A2(dp_n49), .B1(dp_z_word[19]), .B2(dp_n47), .ZN(dp_n381) );
  AOI22_X1 dp_U214 ( .A1(dp_data_mem_ex_o[20]), .A2(dp_n49), .B1(dp_z_word[20]), .B2(dp_n46), .ZN(dp_n380) );
  OAI221_X1 dp_U213 ( .B1(dp_n280), .B2(dp_n52), .C1(dp_n71), .C2(dp_n346), 
        .A(dp_n380), .ZN(dp_n984) );
  AOI22_X1 dp_U212 ( .A1(dp_data_mem_ex_o[21]), .A2(dp_n51), .B1(dp_z_word[21]), .B2(dp_n46), .ZN(dp_n379) );
  OAI221_X1 dp_U211 ( .B1(dp_n281), .B2(dp_n52), .C1(dp_n73), .C2(dp_n345), 
        .A(dp_n379), .ZN(dp_n983) );
  AOI22_X1 dp_U210 ( .A1(dp_data_mem_ex_o[22]), .A2(dp_n49), .B1(dp_z_word[22]), .B2(dp_n46), .ZN(dp_n378) );
  OAI221_X1 dp_U209 ( .B1(dp_n282), .B2(dp_n52), .C1(dp_n71), .C2(dp_n344), 
        .A(dp_n378), .ZN(dp_n982) );
  AOI22_X1 dp_U208 ( .A1(dp_data_mem_ex_o[23]), .A2(dp_n51), .B1(dp_z_word[23]), .B2(dp_n46), .ZN(dp_n377) );
  OAI221_X1 dp_U207 ( .B1(dp_n283), .B2(dp_n52), .C1(dp_n72), .C2(dp_n343), 
        .A(dp_n377), .ZN(dp_n981) );
  AOI22_X1 dp_U206 ( .A1(dp_data_mem_ex_o[24]), .A2(dp_n49), .B1(dp_z_word[24]), .B2(dp_n46), .ZN(dp_n376) );
  OAI221_X1 dp_U205 ( .B1(dp_n284), .B2(dp_n52), .C1(dp_n73), .C2(dp_n342), 
        .A(dp_n376), .ZN(dp_n980) );
  AOI22_X1 dp_U204 ( .A1(dp_data_mem_ex_o[25]), .A2(dp_n49), .B1(dp_z_word[25]), .B2(dp_n46), .ZN(dp_n375) );
  OAI221_X1 dp_U203 ( .B1(dp_n285), .B2(dp_n52), .C1(dp_n71), .C2(dp_n341), 
        .A(dp_n375), .ZN(dp_n979) );
  AOI22_X1 dp_U202 ( .A1(dp_data_mem_ex_o[26]), .A2(dp_n51), .B1(dp_z_word[26]), .B2(dp_n46), .ZN(dp_n374) );
  OAI221_X1 dp_U201 ( .B1(dp_n286), .B2(dp_n52), .C1(dp_n71), .C2(dp_n340), 
        .A(dp_n374), .ZN(dp_n978) );
  AOI22_X1 dp_U200 ( .A1(dp_data_mem_ex_o[27]), .A2(dp_n49), .B1(dp_z_word[27]), .B2(dp_n46), .ZN(dp_n373) );
  OAI221_X1 dp_U199 ( .B1(dp_n287), .B2(dp_n52), .C1(dp_n72), .C2(dp_n339), 
        .A(dp_n373), .ZN(dp_n977) );
  AOI22_X1 dp_U198 ( .A1(dp_data_mem_ex_o[28]), .A2(dp_n51), .B1(dp_z_word[28]), .B2(dp_n46), .ZN(dp_n372) );
  OAI221_X1 dp_U197 ( .B1(dp_n288), .B2(dp_n52), .C1(dp_n73), .C2(dp_n338), 
        .A(dp_n372), .ZN(dp_n976) );
  AOI22_X1 dp_U196 ( .A1(dp_data_mem_ex_o[29]), .A2(dp_n49), .B1(dp_z_word[29]), .B2(dp_n46), .ZN(dp_n371) );
  OAI221_X1 dp_U195 ( .B1(dp_n289), .B2(dp_n52), .C1(dp_n71), .C2(dp_n337), 
        .A(dp_n371), .ZN(dp_n975) );
  AOI22_X1 dp_U194 ( .A1(dp_data_mem_ex_o[30]), .A2(dp_n51), .B1(dp_z_word[30]), .B2(dp_n46), .ZN(dp_n370) );
  OAI221_X1 dp_U193 ( .B1(dp_n290), .B2(dp_n52), .C1(dp_n72), .C2(dp_n336), 
        .A(dp_n370), .ZN(dp_n974) );
  AOI22_X1 dp_U192 ( .A1(dp_data_mem_ex_o[31]), .A2(dp_n50), .B1(dp_z_word[31]), .B2(dp_n46), .ZN(dp_n367) );
  OAI221_X1 dp_U191 ( .B1(dp_n291), .B2(dp_n52), .C1(dp_n72), .C2(dp_n335), 
        .A(dp_n367), .ZN(dp_n973) );
  AOI22_X1 dp_U190 ( .A1(dp_data_mem_ex_o[0]), .A2(dp_n50), .B1(dp_z_word[0]), 
        .B2(dp_n48), .ZN(dp_n401) );
  OAI221_X1 dp_U189 ( .B1(dp_n260), .B2(dp_n54), .C1(dp_n73), .C2(dp_n400), 
        .A(dp_n401), .ZN(dp_n1004) );
  AOI22_X1 dp_U188 ( .A1(dp_data_mem_ex_o[1]), .A2(dp_n50), .B1(dp_z_word[1]), 
        .B2(dp_n48), .ZN(dp_n399) );
  OAI221_X1 dp_U187 ( .B1(dp_n261), .B2(dp_n54), .C1(dp_n71), .C2(dp_n365), 
        .A(dp_n399), .ZN(dp_n1003) );
  AOI22_X1 dp_U186 ( .A1(dp_data_mem_ex_o[2]), .A2(dp_n50), .B1(dp_z_word[2]), 
        .B2(dp_n48), .ZN(dp_n398) );
  OAI221_X1 dp_U185 ( .B1(dp_n262), .B2(dp_n54), .C1(dp_n72), .C2(dp_n364), 
        .A(dp_n398), .ZN(dp_n1002) );
  AOI22_X1 dp_U184 ( .A1(dp_data_mem_ex_o[3]), .A2(dp_n50), .B1(dp_z_word[3]), 
        .B2(dp_n48), .ZN(dp_n397) );
  OAI221_X1 dp_U183 ( .B1(dp_n263), .B2(dp_n54), .C1(dp_n73), .C2(dp_n363), 
        .A(dp_n397), .ZN(dp_n1001) );
  AOI22_X1 dp_U182 ( .A1(dp_data_mem_ex_o[4]), .A2(dp_n50), .B1(dp_z_word[4]), 
        .B2(dp_n48), .ZN(dp_n396) );
  OAI221_X1 dp_U181 ( .B1(dp_n264), .B2(dp_n54), .C1(dp_n71), .C2(dp_n362), 
        .A(dp_n396), .ZN(dp_n1000) );
  AOI22_X1 dp_U180 ( .A1(dp_data_mem_ex_o[5]), .A2(dp_n50), .B1(dp_z_word[5]), 
        .B2(dp_n48), .ZN(dp_n395) );
  OAI221_X1 dp_U179 ( .B1(dp_n265), .B2(dp_n54), .C1(dp_n72), .C2(dp_n361), 
        .A(dp_n395), .ZN(dp_n999) );
  AOI22_X1 dp_U178 ( .A1(dp_data_mem_ex_o[6]), .A2(dp_n50), .B1(dp_z_word[6]), 
        .B2(dp_n48), .ZN(dp_n394) );
  OAI221_X1 dp_U177 ( .B1(dp_n266), .B2(dp_n54), .C1(dp_n73), .C2(dp_n360), 
        .A(dp_n394), .ZN(dp_n998) );
  AOI22_X1 dp_U176 ( .A1(dp_data_mem_ex_o[7]), .A2(dp_n50), .B1(dp_z_word[7]), 
        .B2(dp_n48), .ZN(dp_n393) );
  OAI221_X1 dp_U175 ( .B1(dp_n267), .B2(dp_n54), .C1(dp_n71), .C2(dp_n359), 
        .A(dp_n393), .ZN(dp_n997) );
  OAI22_X1 dp_U174 ( .A1(dp_n66), .A2(dp_n516), .B1(dp_n60), .B2(dp_n293), 
        .ZN(dp_n1009) );
  OAI22_X1 dp_U173 ( .A1(dp_n66), .A2(dp_n518), .B1(dp_n60), .B2(dp_n294), 
        .ZN(dp_n1008) );
  OAI22_X1 dp_U172 ( .A1(dp_n66), .A2(dp_n520), .B1(dp_n60), .B2(dp_n295), 
        .ZN(dp_n1007) );
  OAI22_X1 dp_U171 ( .A1(dp_n66), .A2(dp_n522), .B1(dp_n60), .B2(dp_n296), 
        .ZN(dp_n1006) );
  OAI22_X1 dp_U170 ( .A1(dp_n66), .A2(dp_n524), .B1(dp_n60), .B2(dp_n297), 
        .ZN(dp_n1005) );
  BUF_X1 dp_U169 ( .A(dp_n1029), .Z(dp_n24) );
  BUF_X1 dp_U168 ( .A(dp_n1029), .Z(dp_n23) );
  BUF_X1 dp_U167 ( .A(dp_n122), .Z(dp_n121) );
  BUF_X1 dp_U166 ( .A(dp_n122), .Z(dp_n119) );
  BUF_X1 dp_U165 ( .A(dp_n122), .Z(dp_n118) );
  BUF_X1 dp_U164 ( .A(dp_n122), .Z(dp_n117) );
  BUF_X1 dp_U163 ( .A(dp_n122), .Z(dp_n116) );
  BUF_X1 dp_U162 ( .A(dp_n122), .Z(dp_n115) );
  BUF_X1 dp_U161 ( .A(dp_n122), .Z(dp_n120) );
  AND2_X2 dp_U160 ( .A1(pipe_clear_n_i), .A2(dp_n112), .ZN(dp_n17) );
  NAND2_X1 dp_U159 ( .A1(pipe_clear_n_i), .A2(dp_n131), .ZN(dp_n132) );
  AND2_X2 dp_U158 ( .A1(pipe_ex_mem_en_i), .A2(pipe_clear_n_i), .ZN(dp_n16) );
  OAI22_X1 dp_U157 ( .A1(dp_n327), .A2(dp_n63), .B1(dp_n57), .B2(dp_n338), 
        .ZN(dp_n945) );
  OAI22_X1 dp_U156 ( .A1(dp_n328), .A2(dp_n63), .B1(dp_n57), .B2(dp_n337), 
        .ZN(dp_n944) );
  OAI22_X1 dp_U155 ( .A1(dp_n329), .A2(dp_n63), .B1(dp_n57), .B2(dp_n336), 
        .ZN(dp_n943) );
  OAI22_X1 dp_U154 ( .A1(dp_n330), .A2(dp_n63), .B1(dp_n57), .B2(dp_n335), 
        .ZN(dp_n942) );
  OAI22_X1 dp_U153 ( .A1(dp_n299), .A2(dp_n61), .B1(dp_n59), .B2(dp_n364), 
        .ZN(dp_n971) );
  OAI22_X1 dp_U152 ( .A1(dp_n300), .A2(dp_n61), .B1(dp_n59), .B2(dp_n363), 
        .ZN(dp_n970) );
  OAI22_X1 dp_U151 ( .A1(dp_n303), .A2(dp_n61), .B1(dp_n59), .B2(dp_n362), 
        .ZN(dp_n969) );
  OAI22_X1 dp_U150 ( .A1(dp_n304), .A2(dp_n61), .B1(dp_n59), .B2(dp_n361), 
        .ZN(dp_n968) );
  OAI22_X1 dp_U149 ( .A1(dp_n305), .A2(dp_n61), .B1(dp_n59), .B2(dp_n360), 
        .ZN(dp_n967) );
  OAI22_X1 dp_U148 ( .A1(dp_n306), .A2(dp_n61), .B1(dp_n59), .B2(dp_n359), 
        .ZN(dp_n966) );
  OAI22_X1 dp_U147 ( .A1(dp_n307), .A2(dp_n61), .B1(dp_n59), .B2(dp_n358), 
        .ZN(dp_n965) );
  OAI22_X1 dp_U146 ( .A1(dp_n308), .A2(dp_n61), .B1(dp_n59), .B2(dp_n357), 
        .ZN(dp_n964) );
  OAI22_X1 dp_U145 ( .A1(dp_n309), .A2(dp_n63), .B1(dp_n59), .B2(dp_n356), 
        .ZN(dp_n963) );
  OAI22_X1 dp_U144 ( .A1(dp_n310), .A2(dp_n62), .B1(dp_n59), .B2(dp_n355), 
        .ZN(dp_n962) );
  OAI22_X1 dp_U143 ( .A1(dp_n311), .A2(dp_n62), .B1(dp_n59), .B2(dp_n354), 
        .ZN(dp_n961) );
  OAI22_X1 dp_U142 ( .A1(dp_n312), .A2(dp_n62), .B1(dp_n59), .B2(dp_n353), 
        .ZN(dp_n960) );
  OAI22_X1 dp_U141 ( .A1(dp_n313), .A2(dp_n62), .B1(dp_n59), .B2(dp_n352), 
        .ZN(dp_n959) );
  OAI22_X1 dp_U140 ( .A1(dp_n314), .A2(dp_n62), .B1(dp_n58), .B2(dp_n351), 
        .ZN(dp_n958) );
  OAI22_X1 dp_U139 ( .A1(dp_n315), .A2(dp_n62), .B1(dp_n58), .B2(dp_n350), 
        .ZN(dp_n957) );
  OAI22_X1 dp_U138 ( .A1(dp_n316), .A2(dp_n62), .B1(dp_n58), .B2(dp_n349), 
        .ZN(dp_n956) );
  OAI22_X1 dp_U137 ( .A1(dp_n317), .A2(dp_n62), .B1(dp_n58), .B2(dp_n348), 
        .ZN(dp_n955) );
  OAI22_X1 dp_U136 ( .A1(dp_n318), .A2(dp_n62), .B1(dp_n58), .B2(dp_n347), 
        .ZN(dp_n954) );
  OAI22_X1 dp_U135 ( .A1(dp_n319), .A2(dp_n62), .B1(dp_n58), .B2(dp_n346), 
        .ZN(dp_n953) );
  OAI22_X1 dp_U134 ( .A1(dp_n320), .A2(dp_n62), .B1(dp_n58), .B2(dp_n345), 
        .ZN(dp_n952) );
  OAI22_X1 dp_U133 ( .A1(dp_n321), .A2(dp_n62), .B1(dp_n58), .B2(dp_n344), 
        .ZN(dp_n951) );
  OAI22_X1 dp_U132 ( .A1(dp_n322), .A2(dp_n63), .B1(dp_n58), .B2(dp_n343), 
        .ZN(dp_n950) );
  OAI22_X1 dp_U131 ( .A1(dp_n323), .A2(dp_n63), .B1(dp_n58), .B2(dp_n342), 
        .ZN(dp_n949) );
  OAI22_X1 dp_U130 ( .A1(dp_n324), .A2(dp_n63), .B1(dp_n58), .B2(dp_n341), 
        .ZN(dp_n948) );
  OAI22_X1 dp_U129 ( .A1(dp_n325), .A2(dp_n63), .B1(dp_n58), .B2(dp_n340), 
        .ZN(dp_n947) );
  OAI22_X1 dp_U128 ( .A1(dp_n326), .A2(dp_n63), .B1(dp_n58), .B2(dp_n339), 
        .ZN(dp_n946) );
  CLKBUF_X1 dp_U127 ( .A(dp_n366), .Z(dp_n54) );
  BUF_X1 dp_U126 ( .A(dp_n366), .Z(dp_n52) );
  NOR2_X1 dp_U125 ( .A1(dp_n1027), .A2(dp_n70), .ZN(dp_n369) );
  OAI22_X1 dp_U124 ( .A1(dp_n254), .A2(dp_n61), .B1(dp_n60), .B2(dp_n400), 
        .ZN(dp_n1015) );
  OAI22_X1 dp_U123 ( .A1(dp_n298), .A2(dp_n61), .B1(dp_n60), .B2(dp_n365), 
        .ZN(dp_n972) );
  NAND2_X1 dp_U122 ( .A1(pipe_clear_n_i), .A2(dp_n61), .ZN(dp_n302) );
  BUF_X1 dp_U121 ( .A(dp_n23), .Z(dp_n22) );
  BUF_X1 dp_U120 ( .A(dp_n24), .Z(dp_n18) );
  BUF_X1 dp_U119 ( .A(dp_n23), .Z(dp_n21) );
  BUF_X1 dp_U118 ( .A(dp_n23), .Z(dp_n20) );
  OR2_X1 dp_U117 ( .A1(pipe_if_id_en_i), .A2(dp_n142), .ZN(dp_n131) );
  INV_X1 dp_U116 ( .A(dp_n16), .ZN(dp_n70) );
  INV_X1 dp_U115 ( .A(dp_n69), .ZN(dp_n103) );
  BUF_X1 dp_U114 ( .A(dp_n369), .Z(dp_n48) );
  BUF_X1 dp_U113 ( .A(dp_n369), .Z(dp_n47) );
  BUF_X1 dp_U112 ( .A(dp_n369), .Z(dp_n46) );
  INV_X1 dp_U111 ( .A(dp_n17), .ZN(dp_n71) );
  INV_X1 dp_U110 ( .A(dp_n17), .ZN(dp_n72) );
  INV_X1 dp_U109 ( .A(dp_n17), .ZN(dp_n73) );
  BUF_X1 dp_U108 ( .A(dp_n68), .Z(dp_n106) );
  BUF_X1 dp_U107 ( .A(dp_n75), .Z(dp_n85) );
  BUF_X1 dp_U106 ( .A(dp_n74), .Z(dp_n77) );
  BUF_X1 dp_U105 ( .A(dp_n74), .Z(dp_n78) );
  BUF_X1 dp_U104 ( .A(dp_n74), .Z(dp_n79) );
  BUF_X1 dp_U103 ( .A(dp_n74), .Z(dp_n80) );
  BUF_X1 dp_U102 ( .A(dp_n74), .Z(dp_n76) );
  CLKBUF_X1 dp_U101 ( .A(dp_n301), .Z(dp_n66) );
  INV_X1 dp_U100 ( .A(dp_n103), .ZN(dp_n100) );
  CLKBUF_X1 dp_U99 ( .A(dp_n301), .Z(dp_n63) );
  CLKBUF_X1 dp_U98 ( .A(dp_n301), .Z(dp_n62) );
  CLKBUF_X1 dp_U97 ( .A(dp_n301), .Z(dp_n64) );
  CLKBUF_X1 dp_U96 ( .A(dp_n301), .Z(dp_n65) );
  BUF_X1 dp_U95 ( .A(dp_n105), .Z(dp_n107) );
  BUF_X1 dp_U94 ( .A(dp_n105), .Z(dp_n108) );
  BUF_X1 dp_U93 ( .A(dp_n88), .Z(dp_n91) );
  BUF_X1 dp_U92 ( .A(dp_n89), .Z(dp_n98) );
  BUF_X1 dp_U91 ( .A(dp_n89), .Z(dp_n97) );
  BUF_X1 dp_U90 ( .A(dp_n89), .Z(dp_n96) );
  BUF_X1 dp_U89 ( .A(dp_n89), .Z(dp_n95) );
  BUF_X1 dp_U88 ( .A(dp_n88), .Z(dp_n94) );
  BUF_X1 dp_U87 ( .A(dp_n88), .Z(dp_n93) );
  BUF_X1 dp_U86 ( .A(dp_n88), .Z(dp_n92) );
  BUF_X1 dp_U85 ( .A(dp_n105), .Z(dp_n109) );
  CLKBUF_X1 dp_U84 ( .A(dp_n68), .Z(dp_n105) );
  CLKBUF_X1 dp_U83 ( .A(dp_n131), .Z(dp_n89) );
  BUF_X2 dp_U82 ( .A(dp_n301), .Z(dp_n61) );
  CLKBUF_X1 dp_U81 ( .A(dp_n106), .Z(dp_n111) );
  OAI22_X4 dp_U80 ( .A1(dp_n115), .A2(dp_n331), .B1(dp_n114), .B2(dp_n254), 
        .ZN(dp_wr_data_id_i[0]) );
  OAI22_X4 dp_U79 ( .A1(dp_n117), .A2(dp_n332), .B1(dp_n113), .B2(dp_n298), 
        .ZN(dp_wr_data_id_i[1]) );
  OAI22_X4 dp_U78 ( .A1(dp_n119), .A2(dp_n333), .B1(dp_n113), .B2(dp_n299), 
        .ZN(dp_wr_data_id_i[2]) );
  OAI22_X4 dp_U77 ( .A1(dp_n120), .A2(dp_n334), .B1(dp_n113), .B2(dp_n300), 
        .ZN(dp_wr_data_id_i[3]) );
  OAI22_X4 dp_U76 ( .A1(dp_n115), .A2(dp_n408), .B1(dp_n114), .B2(dp_n309), 
        .ZN(dp_wr_data_id_i[10]) );
  OAI22_X4 dp_U75 ( .A1(dp_n116), .A2(dp_n519), .B1(wb_mux_sel_i), .B2(dp_n316), .ZN(dp_wr_data_id_i[17]) );
  OAI22_X4 dp_U74 ( .A1(dp_n120), .A2(dp_n402), .B1(dp_n113), .B2(dp_n303), 
        .ZN(dp_wr_data_id_i[4]) );
  OAI22_X4 dp_U73 ( .A1(dp_n115), .A2(dp_n409), .B1(dp_n114), .B2(dp_n310), 
        .ZN(dp_wr_data_id_i[11]) );
  OAI22_X4 dp_U72 ( .A1(dp_n116), .A2(dp_n521), .B1(wb_mux_sel_i), .B2(dp_n317), .ZN(dp_wr_data_id_i[18]) );
  OAI22_X4 dp_U71 ( .A1(dp_n120), .A2(dp_n403), .B1(dp_n113), .B2(dp_n304), 
        .ZN(dp_wr_data_id_i[5]) );
  OAI22_X4 dp_U70 ( .A1(dp_n115), .A2(dp_n410), .B1(dp_n114), .B2(dp_n311), 
        .ZN(dp_wr_data_id_i[12]) );
  OAI22_X4 dp_U69 ( .A1(dp_n117), .A2(dp_n523), .B1(dp_n113), .B2(dp_n318), 
        .ZN(dp_wr_data_id_i[19]) );
  OAI22_X4 dp_U68 ( .A1(dp_n120), .A2(dp_n404), .B1(dp_n113), .B2(dp_n305), 
        .ZN(dp_wr_data_id_i[6]) );
  OAI22_X4 dp_U67 ( .A1(dp_n115), .A2(dp_n411), .B1(dp_n114), .B2(dp_n312), 
        .ZN(dp_wr_data_id_i[13]) );
  OAI22_X4 dp_U66 ( .A1(dp_n117), .A2(dp_n525), .B1(dp_n113), .B2(dp_n319), 
        .ZN(dp_wr_data_id_i[20]) );
  INV_X2 dp_U65 ( .A(dp_n121), .ZN(dp_n113) );
  OAI22_X4 dp_U64 ( .A1(dp_n120), .A2(dp_n405), .B1(dp_n113), .B2(dp_n306), 
        .ZN(dp_wr_data_id_i[7]) );
  OAI22_X4 dp_U63 ( .A1(dp_n121), .A2(dp_n406), .B1(dp_n113), .B2(dp_n307), 
        .ZN(dp_wr_data_id_i[8]) );
  OAI22_X4 dp_U62 ( .A1(dp_n116), .A2(dp_n412), .B1(dp_n114), .B2(dp_n313), 
        .ZN(dp_wr_data_id_i[14]) );
  OAI22_X4 dp_U61 ( .A1(dp_n117), .A2(dp_n584), .B1(wb_mux_sel_i), .B2(dp_n320), .ZN(dp_wr_data_id_i[21]) );
  OAI22_X4 dp_U60 ( .A1(dp_n118), .A2(dp_n586), .B1(wb_mux_sel_i), .B2(dp_n322), .ZN(dp_wr_data_id_i[23]) );
  OAI22_X4 dp_U59 ( .A1(dp_n121), .A2(dp_n407), .B1(dp_n113), .B2(dp_n308), 
        .ZN(dp_wr_data_id_i[9]) );
  OAI22_X4 dp_U58 ( .A1(dp_n116), .A2(dp_n413), .B1(dp_n114), .B2(dp_n314), 
        .ZN(dp_wr_data_id_i[15]) );
  OAI22_X4 dp_U57 ( .A1(dp_n117), .A2(dp_n585), .B1(dp_n113), .B2(dp_n321), 
        .ZN(dp_wr_data_id_i[22]) );
  OAI22_X4 dp_U56 ( .A1(dp_n116), .A2(dp_n517), .B1(dp_n114), .B2(dp_n315), 
        .ZN(dp_wr_data_id_i[16]) );
  OAI22_X4 dp_U55 ( .A1(dp_n118), .A2(dp_n587), .B1(wb_mux_sel_i), .B2(dp_n323), .ZN(dp_wr_data_id_i[24]) );
  OAI22_X4 dp_U54 ( .A1(dp_n119), .A2(dp_n591), .B1(dp_n113), .B2(dp_n327), 
        .ZN(dp_wr_data_id_i[28]) );
  OAI22_X4 dp_U53 ( .A1(dp_n118), .A2(dp_n588), .B1(wb_mux_sel_i), .B2(dp_n324), .ZN(dp_wr_data_id_i[25]) );
  OAI22_X4 dp_U52 ( .A1(dp_n119), .A2(dp_n592), .B1(dp_n113), .B2(dp_n328), 
        .ZN(dp_wr_data_id_i[29]) );
  BUF_X2 dp_U51 ( .A(dp_n368), .Z(dp_n49) );
  BUF_X2 dp_U50 ( .A(dp_n368), .Z(dp_n50) );
  BUF_X2 dp_U49 ( .A(dp_n88), .Z(dp_n90) );
  BUF_X2 dp_U48 ( .A(dp_n132), .Z(dp_n75) );
  BUF_X2 dp_U47 ( .A(dp_n75), .Z(dp_n84) );
  BUF_X2 dp_U46 ( .A(dp_n368), .Z(dp_n51) );
  OR2_X1 dp_U45 ( .A1(pipe_if_id_en_i), .A2(dp_n142), .ZN(dp_n301) );
  INV_X4 dp_U44 ( .A(dp_n16), .ZN(dp_n67) );
  BUF_X2 dp_U43 ( .A(dp_n366), .Z(dp_n53) );
  INV_X1 dp_U42 ( .A(dp_n67), .ZN(dp_n15) );
  NAND3_X1 dp_U41 ( .A1(dp_n13), .A2(dp_n14), .A3(dp_n381), .ZN(dp_n985) );
  OR2_X1 dp_U40 ( .A1(dp_n72), .A2(dp_n347), .ZN(dp_n14) );
  OR2_X1 dp_U39 ( .A1(dp_n279), .A2(dp_n53), .ZN(dp_n13) );
  BUF_X2 dp_U38 ( .A(dp_n75), .Z(dp_n87) );
  BUF_X1 dp_U37 ( .A(dp_n131), .Z(dp_n88) );
  INV_X8 dp_U36 ( .A(RST), .ZN(dp_n1029) );
  OAI22_X1 dp_U35 ( .A1(dp_n119), .A2(dp_n1025), .B1(dp_n113), .B2(dp_n330), 
        .ZN(dp_wr_data_id_i[31]) );
  INV_X1 dp_U34 ( .A(dp_wr_data_id_i[31]), .ZN(dp_n11) );
  OAI22_X1 dp_U33 ( .A1(dp_n119), .A2(dp_n593), .B1(dp_n113), .B2(dp_n329), 
        .ZN(dp_wr_data_id_i[30]) );
  INV_X1 dp_U32 ( .A(dp_wr_data_id_i[30]), .ZN(dp_n9) );
  OAI22_X1 dp_U31 ( .A1(dp_n118), .A2(dp_n590), .B1(dp_n113), .B2(dp_n326), 
        .ZN(dp_wr_data_id_i[27]) );
  INV_X1 dp_U30 ( .A(dp_wr_data_id_i[27]), .ZN(dp_n7) );
  OAI22_X1 dp_U29 ( .A1(dp_n118), .A2(dp_n589), .B1(dp_n113), .B2(dp_n325), 
        .ZN(dp_wr_data_id_i[26]) );
  INV_X1 dp_U28 ( .A(dp_wr_data_id_i[26]), .ZN(dp_n5) );
  CLKBUF_X1 dp_U27 ( .A(dp_n24), .Z(dp_n19) );
  INV_X1 dp_U26 ( .A(dp_n103), .ZN(dp_n101) );
  INV_X1 dp_U25 ( .A(dp_n103), .ZN(dp_n4) );
  INV_X1 dp_U24 ( .A(dp_n103), .ZN(dp_n3) );
  NAND2_X2 dp_U23 ( .A1(dp_n106), .A2(pipe_clear_n_i), .ZN(dp_n69) );
  INV_X2 dp_U22 ( .A(dp_n69), .ZN(dp_n104) );
  BUF_X2 dp_U21 ( .A(dp_n302), .Z(dp_n60) );
  BUF_X2 dp_U20 ( .A(dp_n302), .Z(dp_n58) );
  BUF_X2 dp_U19 ( .A(dp_n302), .Z(dp_n59) );
  BUF_X2 dp_U18 ( .A(dp_n302), .Z(dp_n57) );
  BUF_X2 dp_U17 ( .A(dp_n302), .Z(dp_n56) );
  BUF_X2 dp_U16 ( .A(dp_n302), .Z(dp_n55) );
  BUF_X2 dp_U15 ( .A(dp_n74), .Z(dp_n81) );
  BUF_X2 dp_U14 ( .A(dp_n75), .Z(dp_n83) );
  BUF_X2 dp_U13 ( .A(dp_n75), .Z(dp_n82) );
  BUF_X2 dp_U12 ( .A(dp_n75), .Z(dp_n86) );
  BUF_X2 dp_U11 ( .A(dp_n106), .Z(dp_n110) );
  INV_X1 dp_U10 ( .A(dp_n11), .ZN(dp_n12) );
  INV_X1 dp_U9 ( .A(dp_n9), .ZN(dp_n10) );
  INV_X1 dp_U8 ( .A(dp_n7), .ZN(dp_n8) );
  INV_X1 dp_U7 ( .A(dp_n5), .ZN(dp_n6) );
  BUF_X1 dp_U6 ( .A(dp_n132), .Z(dp_n74) );
  DFFR_X2 dp_npc_id_i_reg_16_ ( .D(dp_n691), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[16]), .QN(dp_n558) );
  DFFR_X2 dp_npc_id_i_reg_17_ ( .D(dp_n692), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[17]), .QN(dp_n559) );
  DFFR_X2 dp_npc_id_i_reg_18_ ( .D(dp_n693), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[18]), .QN(dp_n560) );
  DFFR_X2 dp_npc_id_i_reg_19_ ( .D(dp_n694), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[19]), .QN(dp_n561) );
  DFFR_X2 dp_npc_id_i_reg_20_ ( .D(dp_n695), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[20]), .QN(dp_n562) );
  DFFR_X2 dp_npc_id_i_reg_21_ ( .D(dp_n696), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[21]), .QN(dp_n563) );
  DFFR_X2 dp_npc_id_i_reg_22_ ( .D(dp_n697), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[22]), .QN(dp_n564) );
  DFFR_X2 dp_npc_id_i_reg_23_ ( .D(dp_n698), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[23]), .QN(dp_n565) );
  DFFR_X2 dp_npc_id_i_reg_24_ ( .D(dp_n699), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[24]), .QN(dp_n566) );
  DFFR_X2 dp_npc_id_i_reg_26_ ( .D(dp_n701), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[26]), .QN(dp_n568) );
  DFFR_X2 dp_npc_id_i_reg_27_ ( .D(dp_n702), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[27]), .QN(dp_n569) );
  DFFR_X2 dp_npc_id_i_reg_25_ ( .D(dp_n700), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[25]), .QN(dp_n567) );
  DFFR_X2 dp_npc_id_i_reg_28_ ( .D(dp_n703), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[28]), .QN(dp_n570) );
  DFFR_X2 dp_npc_id_i_reg_29_ ( .D(dp_n704), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[29]), .QN(dp_n571) );
  DFFR_X2 dp_npc_id_i_reg_30_ ( .D(dp_n705), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[30]), .QN(dp_n572) );
  DFFR_X1 dp_data_mem_mem_i_reg_20_ ( .D(dp_n984), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[20]) );
  DFFR_X1 dp_data_mem_mem_i_reg_21_ ( .D(dp_n983), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[21]) );
  DFFR_X1 dp_data_mem_mem_i_reg_22_ ( .D(dp_n982), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[22]) );
  DFFR_X1 dp_data_mem_mem_i_reg_23_ ( .D(dp_n981), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[23]) );
  DFFR_X1 dp_data_mem_mem_i_reg_24_ ( .D(dp_n980), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[24]) );
  DFFR_X1 dp_data_mem_mem_i_reg_25_ ( .D(dp_n979), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[25]) );
  DFFR_X1 dp_data_mem_mem_i_reg_26_ ( .D(dp_n978), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[26]) );
  DFFR_X1 dp_data_mem_mem_i_reg_27_ ( .D(dp_n977), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[27]) );
  DFFR_X1 dp_data_mem_mem_i_reg_28_ ( .D(dp_n976), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[28]) );
  DFFR_X1 dp_data_mem_mem_i_reg_29_ ( .D(dp_n975), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[29]) );
  DFFR_X1 dp_data_mem_mem_i_reg_30_ ( .D(dp_n974), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[30]) );
  DFFR_X1 dp_data_mem_mem_i_reg_31_ ( .D(dp_n973), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[31]) );
  DFFR_X1 dp_data_mem_mem_i_reg_8_ ( .D(dp_n996), .CK(CLK), .RN(dp_n1029), .Q(
        DRAM_DATA[8]) );
  DFFR_X1 dp_data_mem_mem_i_reg_9_ ( .D(dp_n995), .CK(CLK), .RN(dp_n1029), .Q(
        DRAM_DATA[9]) );
  DFFR_X1 dp_data_mem_mem_i_reg_10_ ( .D(dp_n994), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[10]) );
  DFFR_X1 dp_data_mem_mem_i_reg_11_ ( .D(dp_n993), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[11]) );
  DFFR_X1 dp_data_mem_mem_i_reg_12_ ( .D(dp_n992), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[12]) );
  DFFR_X1 dp_data_mem_mem_i_reg_13_ ( .D(dp_n991), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[13]) );
  DFFR_X1 dp_data_mem_mem_i_reg_14_ ( .D(dp_n990), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[14]) );
  DFFR_X1 dp_data_mem_mem_i_reg_15_ ( .D(dp_n989), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[15]) );
  DFFR_X1 dp_data_mem_mem_i_reg_16_ ( .D(dp_n988), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[16]) );
  DFFR_X1 dp_data_mem_mem_i_reg_17_ ( .D(dp_n987), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[17]) );
  DFFR_X1 dp_data_mem_mem_i_reg_18_ ( .D(dp_n986), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[18]) );
  DFFR_X1 dp_data_mem_mem_i_reg_0_ ( .D(dp_n1004), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[0]) );
  DFFR_X1 dp_data_mem_mem_i_reg_1_ ( .D(dp_n1003), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[1]) );
  DFFR_X1 dp_data_mem_mem_i_reg_2_ ( .D(dp_n1002), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[2]) );
  DFFR_X1 dp_data_mem_mem_i_reg_3_ ( .D(dp_n1001), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[3]) );
  DFFR_X1 dp_data_mem_mem_i_reg_4_ ( .D(dp_n1000), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[4]) );
  DFFR_X1 dp_data_mem_mem_i_reg_5_ ( .D(dp_n999), .CK(CLK), .RN(dp_n1029), .Q(
        DRAM_DATA[5]) );
  DFFR_X1 dp_data_mem_mem_i_reg_6_ ( .D(dp_n998), .CK(CLK), .RN(dp_n1029), .Q(
        DRAM_DATA[6]) );
  DFFR_X1 dp_data_mem_mem_i_reg_7_ ( .D(dp_n997), .CK(CLK), .RN(dp_n1029), .Q(
        DRAM_DATA[7]) );
  DFFR_X1 dp_data_mem_wb_i_reg_10_ ( .D(dp_n963), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n309) );
  DFFR_X1 dp_data_mem_wb_i_reg_11_ ( .D(dp_n962), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n310) );
  DFFR_X1 dp_data_mem_wb_i_reg_12_ ( .D(dp_n961), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n311) );
  DFFR_X1 dp_data_mem_wb_i_reg_13_ ( .D(dp_n960), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n312) );
  DFFR_X1 dp_data_mem_wb_i_reg_14_ ( .D(dp_n959), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n313) );
  DFFR_X1 dp_data_mem_wb_i_reg_15_ ( .D(dp_n958), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n314) );
  DFFR_X1 dp_data_mem_wb_i_reg_16_ ( .D(dp_n957), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n315) );
  DFFR_X1 dp_data_mem_wb_i_reg_17_ ( .D(dp_n956), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n316) );
  DFFR_X1 dp_data_mem_wb_i_reg_18_ ( .D(dp_n955), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n317) );
  DFFR_X1 dp_data_mem_wb_i_reg_19_ ( .D(dp_n954), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n318) );
  DFFR_X1 dp_data_mem_wb_i_reg_20_ ( .D(dp_n953), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n319) );
  DFFR_X1 dp_data_mem_wb_i_reg_21_ ( .D(dp_n952), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n320) );
  DFFR_X1 dp_data_mem_wb_i_reg_22_ ( .D(dp_n951), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n321) );
  DFFR_X1 dp_data_mem_wb_i_reg_23_ ( .D(dp_n950), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n322) );
  DFFR_X1 dp_data_mem_wb_i_reg_24_ ( .D(dp_n949), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n323) );
  DFFR_X1 dp_data_mem_wb_i_reg_25_ ( .D(dp_n948), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n324) );
  DFFR_X1 dp_data_mem_wb_i_reg_26_ ( .D(dp_n947), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n325) );
  DFFR_X1 dp_data_mem_wb_i_reg_27_ ( .D(dp_n946), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n326) );
  DFFR_X1 dp_data_mem_mem_i_reg_19_ ( .D(dp_n985), .CK(CLK), .RN(dp_n1029), 
        .Q(DRAM_DATA[19]) );
  DFFR_X1 dp_data_mem_wb_i_reg_2_ ( .D(dp_n971), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n299) );
  DFFR_X1 dp_data_mem_wb_i_reg_3_ ( .D(dp_n970), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n300) );
  DFFR_X1 dp_data_mem_wb_i_reg_4_ ( .D(dp_n969), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n303) );
  DFFR_X1 dp_data_mem_wb_i_reg_5_ ( .D(dp_n968), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n304) );
  DFFR_X1 dp_data_mem_wb_i_reg_6_ ( .D(dp_n967), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n305) );
  DFFR_X1 dp_data_mem_wb_i_reg_7_ ( .D(dp_n966), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n306) );
  DFFR_X1 dp_data_mem_wb_i_reg_8_ ( .D(dp_n965), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n307) );
  DFFR_X1 dp_data_mem_wb_i_reg_9_ ( .D(dp_n964), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n308) );
  DFFR_X1 dp_alu_out_wb_i_reg_0_ ( .D(dp_n909), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n331) );
  DFFR_X1 dp_alu_out_wb_i_reg_1_ ( .D(dp_n908), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n332) );
  DFFR_X1 dp_alu_out_wb_i_reg_2_ ( .D(dp_n907), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n333) );
  DFFR_X1 dp_alu_out_wb_i_reg_3_ ( .D(dp_n906), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n334) );
  DFFR_X1 dp_alu_out_wb_i_reg_4_ ( .D(dp_n905), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n402) );
  DFFR_X1 dp_alu_out_wb_i_reg_5_ ( .D(dp_n904), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n403) );
  DFFR_X1 dp_alu_out_wb_i_reg_6_ ( .D(dp_n903), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n404) );
  DFFR_X1 dp_alu_out_wb_i_reg_7_ ( .D(dp_n902), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n405) );
  DFFR_X1 dp_alu_out_wb_i_reg_8_ ( .D(dp_n901), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n406) );
  DFFR_X1 dp_alu_out_wb_i_reg_9_ ( .D(dp_n900), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n407) );
  DFFR_X1 dp_alu_out_wb_i_reg_10_ ( .D(dp_n899), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n408) );
  DFFR_X1 dp_alu_out_wb_i_reg_11_ ( .D(dp_n898), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n409) );
  DFFR_X1 dp_alu_out_wb_i_reg_12_ ( .D(dp_n897), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n410) );
  DFFR_X1 dp_alu_out_wb_i_reg_13_ ( .D(dp_n896), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n411) );
  DFFR_X1 dp_alu_out_wb_i_reg_14_ ( .D(dp_n895), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n412) );
  DFFR_X1 dp_alu_out_wb_i_reg_15_ ( .D(dp_n894), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n413) );
  DFFR_X1 dp_alu_out_wb_i_reg_16_ ( .D(dp_n893), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n517) );
  DFFR_X1 dp_alu_out_wb_i_reg_17_ ( .D(dp_n892), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n519) );
  DFFR_X1 dp_alu_out_wb_i_reg_18_ ( .D(dp_n891), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n521) );
  DFFR_X1 dp_alu_out_wb_i_reg_19_ ( .D(dp_n890), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n523) );
  DFFR_X1 dp_alu_out_wb_i_reg_20_ ( .D(dp_n889), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n525) );
  DFFR_X1 dp_alu_out_wb_i_reg_21_ ( .D(dp_n888), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n584) );
  DFFR_X1 dp_alu_out_wb_i_reg_22_ ( .D(dp_n887), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n585) );
  DFFR_X1 dp_alu_out_wb_i_reg_23_ ( .D(dp_n886), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n586) );
  DFFR_X1 dp_alu_out_wb_i_reg_24_ ( .D(dp_n885), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n587) );
  DFFR_X1 dp_alu_out_wb_i_reg_25_ ( .D(dp_n884), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n588) );
  DFFR_X1 dp_alu_out_wb_i_reg_26_ ( .D(dp_n883), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n589) );
  DFFR_X1 dp_alu_out_wb_i_reg_27_ ( .D(dp_n882), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n590) );
  DFFR_X1 dp_alu_out_wb_i_reg_28_ ( .D(dp_n881), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n591) );
  DFFR_X1 dp_alu_out_wb_i_reg_29_ ( .D(dp_n880), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n592) );
  DFFR_X1 dp_alu_out_wb_i_reg_30_ ( .D(dp_n879), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n593) );
  DFFR_X1 dp_alu_out_wb_i_reg_31_ ( .D(dp_n878), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n1025) );
  DFFR_X1 dp_data_mem_wb_i_reg_28_ ( .D(dp_n945), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n327) );
  DFFR_X1 dp_data_mem_wb_i_reg_29_ ( .D(dp_n944), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n328) );
  DFFR_X1 dp_data_mem_wb_i_reg_30_ ( .D(dp_n943), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n329) );
  DFFR_X1 dp_data_mem_wb_i_reg_31_ ( .D(dp_n942), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n330) );
  DFFR_X1 dp_data_mem_wb_i_reg_0_ ( .D(dp_n1015), .CK(CLK), .RN(dp_n1029), 
        .QN(dp_n254) );
  DFFR_X1 dp_data_mem_wb_i_reg_1_ ( .D(dp_n972), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n298) );
  DFFR_X1 dp_npc_ex_i_reg_3_ ( .D(dp_n720), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[3]), .QN(dp_n263) );
  DFFR_X1 dp_npc_ex_i_reg_4_ ( .D(dp_n721), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[4]), .QN(dp_n264) );
  DFFR_X1 dp_npc_ex_i_reg_6_ ( .D(dp_n723), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[6]), .QN(dp_n266) );
  DFFR_X1 dp_npc_ex_i_reg_11_ ( .D(dp_n728), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[11]), .QN(dp_n271) );
  DFFR_X1 dp_npc_ex_i_reg_18_ ( .D(dp_n735), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[18]), .QN(dp_n278) );
  DFFR_X1 dp_npc_ex_i_reg_19_ ( .D(dp_n736), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[19]), .QN(dp_n279) );
  DFFR_X1 dp_npc_ex_i_reg_20_ ( .D(dp_n737), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[20]), .QN(dp_n280) );
  DFFR_X1 dp_npc_ex_i_reg_24_ ( .D(dp_n741), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[24]), .QN(dp_n284) );
  DFFR_X1 dp_npc_ex_i_reg_26_ ( .D(dp_n743), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[26]), .QN(dp_n286) );
  DFFR_X1 dp_npc_ex_i_reg_5_ ( .D(dp_n722), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[5]), .QN(dp_n265) );
  DFFR_X1 dp_npc_ex_i_reg_7_ ( .D(dp_n724), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[7]), .QN(dp_n267) );
  DFFR_X1 dp_npc_ex_i_reg_8_ ( .D(dp_n725), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[8]), .QN(dp_n268) );
  DFFR_X1 dp_npc_ex_i_reg_9_ ( .D(dp_n726), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[9]), .QN(dp_n269) );
  DFFR_X1 dp_npc_ex_i_reg_10_ ( .D(dp_n727), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[10]), .QN(dp_n270) );
  DFFR_X1 dp_npc_ex_i_reg_12_ ( .D(dp_n729), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[12]), .QN(dp_n272) );
  DFFR_X1 dp_npc_ex_i_reg_13_ ( .D(dp_n730), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[13]), .QN(dp_n273) );
  DFFR_X1 dp_npc_ex_i_reg_14_ ( .D(dp_n731), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[14]), .QN(dp_n274) );
  DFFR_X1 dp_npc_ex_i_reg_15_ ( .D(dp_n732), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[15]), .QN(dp_n275) );
  DFFR_X1 dp_npc_ex_i_reg_16_ ( .D(dp_n733), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[16]), .QN(dp_n276) );
  DFFR_X1 dp_npc_ex_i_reg_17_ ( .D(dp_n734), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[17]), .QN(dp_n277) );
  DFFR_X1 dp_npc_ex_i_reg_21_ ( .D(dp_n738), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[21]), .QN(dp_n281) );
  DFFR_X1 dp_npc_ex_i_reg_22_ ( .D(dp_n739), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[22]), .QN(dp_n282) );
  DFFR_X1 dp_npc_ex_i_reg_23_ ( .D(dp_n740), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[23]), .QN(dp_n283) );
  DFFR_X1 dp_npc_ex_i_reg_25_ ( .D(dp_n742), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[25]), .QN(dp_n285) );
  DFFR_X1 dp_npc_ex_i_reg_27_ ( .D(dp_n744), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[27]), .QN(dp_n287) );
  DFFR_X1 dp_npc_ex_i_reg_28_ ( .D(dp_n745), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[28]), .QN(dp_n288) );
  DFFR_X1 dp_npc_ex_i_reg_29_ ( .D(dp_n746), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[29]), .QN(dp_n289) );
  DFFR_X1 dp_npc_ex_i_reg_30_ ( .D(dp_n747), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[30]), .QN(dp_n290) );
  DFFR_X1 dp_npc_ex_i_reg_31_ ( .D(dp_n748), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[31]), .QN(dp_n291) );
  DFFR_X1 dp_npc_ex_i_reg_0_ ( .D(dp_n717), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[0]), .QN(dp_n260) );
  DFFR_X1 dp_npc_ex_i_reg_1_ ( .D(dp_n718), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[1]), .QN(dp_n261) );
  DFFR_X1 dp_npc_ex_i_reg_2_ ( .D(dp_n719), .CK(CLK), .RN(dp_n1029), .Q(
        dp_npc_ex_i[2]), .QN(dp_n262) );
  DFFR_X1 dp_rd_fwd_mem_i_reg_0_ ( .D(dp_n1014), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n293) );
  DFFR_X1 dp_rd_fwd_mem_i_reg_1_ ( .D(dp_n1013), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n294) );
  DFFR_X1 dp_rd_fwd_mem_i_reg_2_ ( .D(dp_n1012), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n295) );
  DFFR_X1 dp_rd_fwd_mem_i_reg_4_ ( .D(dp_n1010), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n297) );
  DFFR_X1 dp_rd_fwd_mem_i_reg_3_ ( .D(dp_n1011), .CK(CLK), .RN(dp_n1029), .QN(
        dp_n296) );
  TBUF_X1 dp_z_word_tri_31_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[31]) );
  TBUF_X1 dp_z_word_tri_30_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[30]) );
  TBUF_X1 dp_z_word_tri_29_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[29]) );
  TBUF_X1 dp_z_word_tri_28_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[28]) );
  TBUF_X1 dp_z_word_tri_27_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[27]) );
  TBUF_X1 dp_z_word_tri_26_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[26]) );
  TBUF_X1 dp_z_word_tri_25_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[25]) );
  TBUF_X1 dp_z_word_tri_24_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[24]) );
  TBUF_X1 dp_z_word_tri_23_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[23]) );
  TBUF_X1 dp_z_word_tri_22_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[22]) );
  TBUF_X1 dp_z_word_tri_21_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[21]) );
  TBUF_X1 dp_z_word_tri_20_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[20]) );
  TBUF_X1 dp_z_word_tri_19_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[19]) );
  TBUF_X1 dp_z_word_tri_18_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[18]) );
  TBUF_X1 dp_z_word_tri_17_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[17]) );
  TBUF_X1 dp_z_word_tri_16_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[16]) );
  TBUF_X1 dp_z_word_tri_15_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[15]) );
  TBUF_X1 dp_z_word_tri_14_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[14]) );
  TBUF_X1 dp_z_word_tri_13_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[13]) );
  TBUF_X1 dp_z_word_tri_12_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[12]) );
  TBUF_X1 dp_z_word_tri_11_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[11]) );
  TBUF_X1 dp_z_word_tri_10_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[10]) );
  TBUF_X1 dp_z_word_tri_9_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[9]) );
  TBUF_X1 dp_z_word_tri_8_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[8]) );
  TBUF_X1 dp_z_word_tri_7_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[7]) );
  TBUF_X1 dp_z_word_tri_6_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[6]) );
  TBUF_X1 dp_z_word_tri_5_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[5]) );
  TBUF_X1 dp_z_word_tri_4_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[4]) );
  TBUF_X1 dp_z_word_tri_3_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[3]) );
  TBUF_X1 dp_z_word_tri_2_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[2]) );
  TBUF_X1 dp_z_word_tri_1_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[1]) );
  TBUF_X1 dp_z_word_tri_0_ ( .A(1'b0), .EN(1'b1), .Z(dp_z_word[0]) );
  NOR3_X2 dp_U752 ( .A1(mem_in_en_i), .A2(npc_wb_en_i), .A3(dp_n70), .ZN(
        dp_n368) );
  NAND3_X1 dp_U753 ( .A1(dp_n16), .A2(dp_n1027), .A3(npc_wb_en_i), .ZN(dp_n366) );
  DFFR_X1 dp_npc_id_i_reg_31_ ( .D(dp_n706), .CK(CLK), .RN(dp_n25), .Q(
        dp_npc_id_o[31]), .QN(dp_n573) );
  DFFR_X1 dp_npc_id_i_reg_15_ ( .D(dp_n690), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[15]), .QN(dp_n557) );
  DFFR_X1 dp_npc_id_i_reg_14_ ( .D(dp_n689), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[14]), .QN(dp_n556) );
  DFFR_X1 dp_npc_id_i_reg_13_ ( .D(dp_n688), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[13]), .QN(dp_n555) );
  DFFR_X1 dp_npc_id_i_reg_12_ ( .D(dp_n687), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[12]), .QN(dp_n554) );
  DFFR_X1 dp_npc_id_i_reg_11_ ( .D(dp_n686), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[11]), .QN(dp_n553) );
  DFFR_X1 dp_npc_id_i_reg_10_ ( .D(dp_n685), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[10]), .QN(dp_n552) );
  DFFR_X1 dp_npc_id_i_reg_9_ ( .D(dp_n684), .CK(CLK), .RN(dp_n26), .Q(
        dp_npc_id_o[9]), .QN(dp_n551) );
  DFFR_X1 dp_npc_id_i_reg_8_ ( .D(dp_n683), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[8]), .QN(dp_n550) );
  DFFR_X1 dp_npc_id_i_reg_7_ ( .D(dp_n682), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[7]), .QN(dp_n549) );
  DFFR_X1 dp_npc_id_i_reg_6_ ( .D(dp_n681), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[6]), .QN(dp_n548) );
  DFFR_X1 dp_npc_id_i_reg_5_ ( .D(dp_n680), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[5]), .QN(dp_n547) );
  DFFR_X1 dp_npc_id_i_reg_4_ ( .D(dp_n679), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[4]), .QN(dp_n546) );
  DFFR_X1 dp_npc_id_i_reg_3_ ( .D(dp_n678), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[3]), .QN(dp_n545) );
  DFFR_X1 dp_npc_id_i_reg_2_ ( .D(dp_n677), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[2]), .QN(dp_n544) );
  DFFR_X1 dp_npc_id_i_reg_1_ ( .D(dp_n676), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[1]), .QN(dp_n543) );
  DFFR_X1 dp_npc_id_i_reg_0_ ( .D(dp_n675), .CK(CLK), .RN(dp_n27), .Q(
        dp_npc_id_o[0]), .QN(dp_n542) );
  DFFR_X1 dp_ir_reg_25_ ( .D(dp_n674), .CK(CLK), .RN(dp_n27), .Q(dp_ir_25_), 
        .QN(dp_n541) );
  DFFR_X1 dp_ir_reg_24_ ( .D(dp_n673), .CK(CLK), .RN(dp_n27), .Q(dp_ir_24_), 
        .QN(dp_n540) );
  DFFR_X1 dp_ir_reg_23_ ( .D(dp_n672), .CK(CLK), .RN(dp_n27), .Q(dp_ir_23_), 
        .QN(dp_n539) );
  DFFR_X1 dp_ir_reg_22_ ( .D(dp_n671), .CK(CLK), .RN(dp_n28), .Q(dp_ir_22_), 
        .QN(dp_n538) );
  DFFR_X1 dp_ir_reg_21_ ( .D(dp_n670), .CK(CLK), .RN(dp_n28), .Q(dp_ir_21_), 
        .QN(dp_n537) );
  DFFR_X1 dp_ir_reg_20_ ( .D(dp_n669), .CK(CLK), .RN(dp_n28), .Q(dp_ir_20_), 
        .QN(dp_n582) );
  DFFR_X1 dp_ir_reg_19_ ( .D(dp_n668), .CK(CLK), .RN(dp_n28), .Q(dp_ir_19_), 
        .QN(dp_n580) );
  DFFR_X1 dp_ir_reg_18_ ( .D(dp_n667), .CK(CLK), .RN(dp_n28), .Q(dp_ir_18_), 
        .QN(dp_n578) );
  DFFR_X1 dp_ir_reg_17_ ( .D(dp_n666), .CK(CLK), .RN(dp_n28), .Q(dp_ir_17_), 
        .QN(dp_n576) );
  DFFR_X1 dp_ir_reg_16_ ( .D(dp_n665), .CK(CLK), .RN(dp_n28), .Q(dp_ir_16_), 
        .QN(dp_n574) );
  DFFR_X1 dp_ir_reg_15_ ( .D(dp_n664), .CK(CLK), .RN(dp_n28), .Q(dp_ir_15_), 
        .QN(dp_n583) );
  DFFR_X1 dp_ir_reg_14_ ( .D(dp_n663), .CK(CLK), .RN(dp_n28), .Q(dp_ir_14_), 
        .QN(dp_n581) );
  DFFR_X1 dp_ir_reg_13_ ( .D(dp_n662), .CK(CLK), .RN(dp_n28), .Q(dp_ir_13_), 
        .QN(dp_n579) );
  DFFR_X1 dp_ir_reg_12_ ( .D(dp_n661), .CK(CLK), .RN(dp_n28), .Q(dp_ir_12_), 
        .QN(dp_n577) );
  DFFR_X1 dp_ir_reg_11_ ( .D(dp_n660), .CK(CLK), .RN(dp_n28), .Q(dp_ir_11_), 
        .QN(dp_n575) );
  DFFR_X1 dp_ir_reg_10_ ( .D(dp_n659), .CK(CLK), .RN(dp_n29), .Q(dp_ir_10_), 
        .QN(dp_n536) );
  DFFR_X1 dp_ir_reg_9_ ( .D(dp_n658), .CK(CLK), .RN(dp_n29), .Q(dp_ir_9_), 
        .QN(dp_n535) );
  DFFR_X1 dp_ir_reg_8_ ( .D(dp_n657), .CK(CLK), .RN(dp_n29), .Q(dp_ir_8_), 
        .QN(dp_n534) );
  DFFR_X1 dp_ir_reg_7_ ( .D(dp_n656), .CK(CLK), .RN(dp_n29), .Q(dp_ir_7_), 
        .QN(dp_n533) );
  DFFR_X1 dp_ir_reg_6_ ( .D(dp_n655), .CK(CLK), .RN(dp_n29), .Q(dp_ir_6_), 
        .QN(dp_n532) );
  DFFR_X1 dp_ir_reg_5_ ( .D(dp_n654), .CK(CLK), .RN(dp_n29), .Q(dp_ir_5_), 
        .QN(dp_n531) );
  DFFR_X1 dp_ir_reg_4_ ( .D(dp_n653), .CK(CLK), .RN(dp_n29), .Q(dp_ir_4_), 
        .QN(dp_n530) );
  DFFR_X1 dp_ir_reg_3_ ( .D(dp_n652), .CK(CLK), .RN(dp_n29), .Q(dp_ir_3_), 
        .QN(dp_n529) );
  DFFR_X1 dp_ir_reg_2_ ( .D(dp_n651), .CK(CLK), .RN(dp_n29), .Q(dp_ir_2_), 
        .QN(dp_n528) );
  DFFR_X1 dp_ir_reg_1_ ( .D(dp_n650), .CK(CLK), .RN(dp_n29), .Q(dp_ir_1_), 
        .QN(dp_n527) );
  DFFR_X1 dp_ir_reg_0_ ( .D(dp_n649), .CK(CLK), .RN(dp_n29), .Q(dp_ir_0_), 
        .QN(dp_n526) );
  DFFR_X1 dp_alu_out_mem_i_reg_31_ ( .D(dp_n910), .CK(CLK), .RN(dp_n29), .Q(
        DRAM_ADDRESS[31]), .QN(dp_n846) );
  DFFR_X1 dp_alu_out_mem_i_reg_30_ ( .D(dp_n911), .CK(CLK), .RN(dp_n30), .Q(
        DRAM_ADDRESS[30]), .QN(dp_n847) );
  DFFR_X1 dp_alu_out_mem_i_reg_29_ ( .D(dp_n912), .CK(CLK), .RN(dp_n30), .Q(
        DRAM_ADDRESS[29]), .QN(dp_n848) );
  DFFR_X1 dp_alu_out_mem_i_reg_28_ ( .D(dp_n913), .CK(CLK), .RN(dp_n30), .Q(
        DRAM_ADDRESS[28]), .QN(dp_n849) );
  DFFR_X1 dp_alu_out_mem_i_reg_27_ ( .D(dp_n914), .CK(CLK), .RN(dp_n30), .Q(
        DRAM_ADDRESS[27]), .QN(dp_n850) );
  DFFR_X1 dp_alu_out_mem_i_reg_26_ ( .D(dp_n915), .CK(CLK), .RN(dp_n30), .Q(
        DRAM_ADDRESS[26]), .QN(dp_n851) );
  DFFR_X1 dp_alu_out_mem_i_reg_25_ ( .D(dp_n916), .CK(CLK), .RN(dp_n30), .Q(
        DRAM_ADDRESS[25]), .QN(dp_n852) );
  DFFR_X1 dp_alu_out_mem_i_reg_24_ ( .D(dp_n917), .CK(CLK), .RN(dp_n31), .Q(
        DRAM_ADDRESS[24]), .QN(dp_n853) );
  DFFR_X1 dp_alu_out_mem_i_reg_23_ ( .D(dp_n918), .CK(CLK), .RN(dp_n31), .Q(
        DRAM_ADDRESS[23]), .QN(dp_n854) );
  DFFR_X1 dp_alu_out_mem_i_reg_22_ ( .D(dp_n919), .CK(CLK), .RN(dp_n31), .Q(
        DRAM_ADDRESS[22]), .QN(dp_n855) );
  DFFR_X1 dp_alu_out_mem_i_reg_21_ ( .D(dp_n920), .CK(CLK), .RN(dp_n31), .Q(
        DRAM_ADDRESS[21]), .QN(dp_n856) );
  DFFR_X1 dp_alu_out_mem_i_reg_20_ ( .D(dp_n921), .CK(CLK), .RN(dp_n31), .Q(
        DRAM_ADDRESS[20]), .QN(dp_n857) );
  DFFR_X1 dp_alu_out_mem_i_reg_19_ ( .D(dp_n922), .CK(CLK), .RN(dp_n31), .Q(
        DRAM_ADDRESS[19]), .QN(dp_n858) );
  DFFR_X1 dp_alu_out_mem_i_reg_18_ ( .D(dp_n923), .CK(CLK), .RN(dp_n32), .Q(
        DRAM_ADDRESS[18]), .QN(dp_n859) );
  DFFR_X1 dp_alu_out_mem_i_reg_17_ ( .D(dp_n924), .CK(CLK), .RN(dp_n32), .Q(
        DRAM_ADDRESS[17]), .QN(dp_n860) );
  DFFR_X1 dp_alu_out_mem_i_reg_16_ ( .D(dp_n925), .CK(CLK), .RN(dp_n32), .Q(
        DRAM_ADDRESS[16]), .QN(dp_n861) );
  DFFR_X1 dp_alu_out_mem_i_reg_15_ ( .D(dp_n926), .CK(CLK), .RN(dp_n32), .Q(
        DRAM_ADDRESS[15]), .QN(dp_n862) );
  DFFR_X1 dp_alu_out_mem_i_reg_14_ ( .D(dp_n927), .CK(CLK), .RN(dp_n32), .Q(
        DRAM_ADDRESS[14]), .QN(dp_n863) );
  DFFR_X1 dp_alu_out_mem_i_reg_13_ ( .D(dp_n928), .CK(CLK), .RN(dp_n32), .Q(
        DRAM_ADDRESS[13]), .QN(dp_n864) );
  DFFR_X1 dp_alu_out_mem_i_reg_12_ ( .D(dp_n929), .CK(CLK), .RN(dp_n33), .Q(
        DRAM_ADDRESS[12]), .QN(dp_n865) );
  DFFR_X1 dp_alu_out_mem_i_reg_11_ ( .D(dp_n930), .CK(CLK), .RN(dp_n33), .Q(
        DRAM_ADDRESS[11]), .QN(dp_n866) );
  DFFR_X1 dp_alu_out_mem_i_reg_10_ ( .D(dp_n931), .CK(CLK), .RN(dp_n33), .Q(
        DRAM_ADDRESS[10]), .QN(dp_n867) );
  DFFR_X1 dp_alu_out_mem_i_reg_9_ ( .D(dp_n932), .CK(CLK), .RN(dp_n33), .Q(
        DRAM_ADDRESS[9]), .QN(dp_n868) );
  DFFR_X1 dp_alu_out_mem_i_reg_8_ ( .D(dp_n933), .CK(CLK), .RN(dp_n33), .Q(
        DRAM_ADDRESS[8]), .QN(dp_n869) );
  DFFR_X1 dp_alu_out_mem_i_reg_7_ ( .D(dp_n934), .CK(CLK), .RN(dp_n33), .Q(
        DRAM_ADDRESS[7]), .QN(dp_n870) );
  DFFR_X1 dp_alu_out_mem_i_reg_6_ ( .D(dp_n935), .CK(CLK), .RN(dp_n34), .Q(
        DRAM_ADDRESS[6]), .QN(dp_n871) );
  DFFR_X1 dp_alu_out_mem_i_reg_5_ ( .D(dp_n936), .CK(CLK), .RN(dp_n34), .Q(
        DRAM_ADDRESS[5]), .QN(dp_n872) );
  DFFR_X1 dp_alu_out_mem_i_reg_4_ ( .D(dp_n937), .CK(CLK), .RN(dp_n34), .Q(
        DRAM_ADDRESS[4]), .QN(dp_n873) );
  DFFR_X1 dp_alu_out_mem_i_reg_3_ ( .D(dp_n938), .CK(CLK), .RN(dp_n34), .Q(
        DRAM_ADDRESS[3]), .QN(dp_n874) );
  DFFR_X1 dp_alu_out_mem_i_reg_2_ ( .D(dp_n939), .CK(CLK), .RN(dp_n34), .Q(
        DRAM_ADDRESS[2]), .QN(dp_n875) );
  DFFR_X1 dp_alu_out_mem_i_reg_1_ ( .D(dp_n940), .CK(CLK), .RN(dp_n34), .Q(
        DRAM_ADDRESS[1]), .QN(dp_n876) );
  DFFR_X1 dp_alu_out_mem_i_reg_0_ ( .D(dp_n941), .CK(CLK), .RN(dp_n24), .Q(
        DRAM_ADDRESS[0]), .QN(dp_n877) );
  DFFR_X1 dp_rd_fwd_wb_i_reg_4_ ( .D(dp_n1005), .CK(CLK), .RN(dp_n35), .Q(
        dp_rd_fwd_wb_i[4]), .QN(dp_n524) );
  DFFR_X1 dp_rd_fwd_wb_i_reg_3_ ( .D(dp_n1006), .CK(CLK), .RN(dp_n35), .Q(
        dp_rd_fwd_wb_i[3]), .QN(dp_n522) );
  DFFR_X1 dp_rd_fwd_wb_i_reg_2_ ( .D(dp_n1007), .CK(CLK), .RN(dp_n35), .Q(
        dp_rd_fwd_wb_i[2]), .QN(dp_n520) );
  DFFR_X1 dp_rd_fwd_wb_i_reg_1_ ( .D(dp_n1008), .CK(CLK), .RN(dp_n35), .Q(
        dp_rd_fwd_wb_i[1]), .QN(dp_n518) );
  DFFR_X1 dp_rd_fwd_wb_i_reg_0_ ( .D(dp_n1009), .CK(CLK), .RN(dp_n36), .Q(
        dp_rd_fwd_wb_i[0]), .QN(dp_n516) );
  DFFR_X1 dp_branch_t_mem_i_reg ( .D(dp_n845), .CK(CLK), .RN(dp_n36), .Q(
        is_zero_i), .QN(dp_n515) );
  DFFR_X1 dp_rf_out1_ex_i_reg_31_ ( .D(dp_n844), .CK(CLK), .RN(dp_n36), .Q(
        dp_rf_out1_ex_i[31]), .QN(dp_n514) );
  DFFR_X1 dp_rf_out1_ex_i_reg_30_ ( .D(dp_n843), .CK(CLK), .RN(dp_n36), .Q(
        dp_rf_out1_ex_i[30]), .QN(dp_n513) );
  DFFR_X1 dp_rf_out1_ex_i_reg_29_ ( .D(dp_n842), .CK(CLK), .RN(dp_n36), .Q(
        dp_rf_out1_ex_i[29]), .QN(dp_n512) );
  DFFR_X1 dp_rf_out1_ex_i_reg_28_ ( .D(dp_n841), .CK(CLK), .RN(dp_n36), .Q(
        dp_rf_out1_ex_i[28]), .QN(dp_n511) );
  DFFR_X1 dp_rf_out1_ex_i_reg_27_ ( .D(dp_n840), .CK(CLK), .RN(dp_n36), .Q(
        dp_rf_out1_ex_i[27]), .QN(dp_n510) );
  DFFR_X1 dp_rf_out1_ex_i_reg_26_ ( .D(dp_n839), .CK(CLK), .RN(dp_n36), .Q(
        dp_rf_out1_ex_i[26]), .QN(dp_n509) );
  DFFR_X1 dp_rf_out1_ex_i_reg_25_ ( .D(dp_n838), .CK(CLK), .RN(dp_n36), .Q(
        dp_rf_out1_ex_i[25]), .QN(dp_n508) );
  DFFR_X1 dp_rf_out1_ex_i_reg_24_ ( .D(dp_n837), .CK(CLK), .RN(dp_n36), .Q(
        dp_rf_out1_ex_i[24]), .QN(dp_n507) );
  DFFR_X1 dp_rf_out1_ex_i_reg_23_ ( .D(dp_n836), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[23]), .QN(dp_n506) );
  DFFR_X1 dp_rf_out1_ex_i_reg_22_ ( .D(dp_n835), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[22]), .QN(dp_n505) );
  DFFR_X1 dp_rf_out1_ex_i_reg_21_ ( .D(dp_n834), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[21]), .QN(dp_n504) );
  DFFR_X1 dp_rf_out1_ex_i_reg_20_ ( .D(dp_n833), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[20]), .QN(dp_n503) );
  DFFR_X1 dp_rf_out1_ex_i_reg_19_ ( .D(dp_n832), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[19]), .QN(dp_n502) );
  DFFR_X1 dp_rf_out1_ex_i_reg_18_ ( .D(dp_n831), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[18]), .QN(dp_n501) );
  DFFR_X1 dp_rf_out1_ex_i_reg_17_ ( .D(dp_n830), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[17]), .QN(dp_n500) );
  DFFR_X1 dp_rf_out1_ex_i_reg_16_ ( .D(dp_n829), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[16]), .QN(dp_n499) );
  DFFR_X1 dp_rf_out1_ex_i_reg_15_ ( .D(dp_n828), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[15]), .QN(dp_n498) );
  DFFR_X1 dp_rf_out1_ex_i_reg_14_ ( .D(dp_n827), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[14]), .QN(dp_n497) );
  DFFR_X1 dp_rf_out1_ex_i_reg_13_ ( .D(dp_n826), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[13]), .QN(dp_n496) );
  DFFR_X1 dp_rf_out1_ex_i_reg_12_ ( .D(dp_n825), .CK(CLK), .RN(dp_n37), .Q(
        dp_rf_out1_ex_i[12]), .QN(dp_n495) );
  DFFR_X1 dp_rf_out1_ex_i_reg_11_ ( .D(dp_n824), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[11]), .QN(dp_n494) );
  DFFR_X1 dp_rf_out1_ex_i_reg_10_ ( .D(dp_n823), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[10]), .QN(dp_n493) );
  DFFR_X1 dp_rf_out1_ex_i_reg_9_ ( .D(dp_n822), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[9]), .QN(dp_n492) );
  DFFR_X1 dp_rf_out1_ex_i_reg_8_ ( .D(dp_n821), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[8]), .QN(dp_n491) );
  DFFR_X1 dp_rf_out1_ex_i_reg_7_ ( .D(dp_n820), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[7]), .QN(dp_n490) );
  DFFR_X1 dp_rf_out1_ex_i_reg_6_ ( .D(dp_n819), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[6]), .QN(dp_n489) );
  DFFR_X1 dp_rf_out1_ex_i_reg_5_ ( .D(dp_n818), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[5]), .QN(dp_n488) );
  DFFR_X1 dp_rf_out1_ex_i_reg_4_ ( .D(dp_n817), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[4]), .QN(dp_n487) );
  DFFR_X1 dp_rf_out1_ex_i_reg_3_ ( .D(dp_n816), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[3]), .QN(dp_n486) );
  DFFR_X1 dp_rf_out1_ex_i_reg_2_ ( .D(dp_n815), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[2]), .QN(dp_n485) );
  DFFR_X1 dp_rf_out1_ex_i_reg_1_ ( .D(dp_n814), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[1]), .QN(dp_n484) );
  DFFR_X1 dp_rf_out1_ex_i_reg_0_ ( .D(dp_n813), .CK(CLK), .RN(dp_n38), .Q(
        dp_rf_out1_ex_i[0]), .QN(dp_n483) );
  DFFR_X1 dp_rf_out2_ex_i_reg_31_ ( .D(dp_n812), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[31]), .QN(dp_n482) );
  DFFR_X1 dp_rf_out2_ex_i_reg_30_ ( .D(dp_n811), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[30]), .QN(dp_n481) );
  DFFR_X1 dp_rf_out2_ex_i_reg_29_ ( .D(dp_n810), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[29]), .QN(dp_n480) );
  DFFR_X1 dp_rf_out2_ex_i_reg_28_ ( .D(dp_n809), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[28]), .QN(dp_n479) );
  DFFR_X1 dp_rf_out2_ex_i_reg_27_ ( .D(dp_n808), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[27]), .QN(dp_n478) );
  DFFR_X1 dp_rf_out2_ex_i_reg_26_ ( .D(dp_n807), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[26]), .QN(dp_n477) );
  DFFR_X1 dp_rf_out2_ex_i_reg_25_ ( .D(dp_n806), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[25]), .QN(dp_n476) );
  DFFR_X1 dp_rf_out2_ex_i_reg_24_ ( .D(dp_n805), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[24]), .QN(dp_n475) );
  DFFR_X1 dp_rf_out2_ex_i_reg_23_ ( .D(dp_n804), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[23]), .QN(dp_n474) );
  DFFR_X1 dp_rf_out2_ex_i_reg_22_ ( .D(dp_n803), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[22]), .QN(dp_n473) );
  DFFR_X1 dp_rf_out2_ex_i_reg_21_ ( .D(dp_n802), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[21]), .QN(dp_n472) );
  DFFR_X1 dp_rf_out2_ex_i_reg_20_ ( .D(dp_n801), .CK(CLK), .RN(dp_n39), .Q(
        dp_data_mem_ex_o[20]), .QN(dp_n471) );
  DFFR_X1 dp_rf_out2_ex_i_reg_19_ ( .D(dp_n800), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[19]), .QN(dp_n470) );
  DFFR_X1 dp_rf_out2_ex_i_reg_18_ ( .D(dp_n799), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[18]), .QN(dp_n469) );
  DFFR_X1 dp_rf_out2_ex_i_reg_17_ ( .D(dp_n798), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[17]), .QN(dp_n468) );
  DFFR_X1 dp_rf_out2_ex_i_reg_16_ ( .D(dp_n797), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[16]), .QN(dp_n467) );
  DFFR_X1 dp_rf_out2_ex_i_reg_15_ ( .D(dp_n796), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[15]), .QN(dp_n466) );
  DFFR_X1 dp_rf_out2_ex_i_reg_14_ ( .D(dp_n795), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[14]), .QN(dp_n465) );
  DFFR_X1 dp_rf_out2_ex_i_reg_13_ ( .D(dp_n794), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[13]), .QN(dp_n464) );
  DFFR_X1 dp_rf_out2_ex_i_reg_12_ ( .D(dp_n793), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[12]), .QN(dp_n463) );
  DFFR_X1 dp_rf_out2_ex_i_reg_11_ ( .D(dp_n792), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[11]), .QN(dp_n462) );
  DFFR_X1 dp_rf_out2_ex_i_reg_10_ ( .D(dp_n791), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[10]), .QN(dp_n461) );
  DFFR_X1 dp_rf_out2_ex_i_reg_9_ ( .D(dp_n790), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[9]), .QN(dp_n460) );
  DFFR_X1 dp_rf_out2_ex_i_reg_8_ ( .D(dp_n789), .CK(CLK), .RN(dp_n40), .Q(
        dp_data_mem_ex_o[8]), .QN(dp_n459) );
  DFFR_X1 dp_rf_out2_ex_i_reg_7_ ( .D(dp_n788), .CK(CLK), .RN(dp_n41), .Q(
        dp_data_mem_ex_o[7]), .QN(dp_n458) );
  DFFR_X1 dp_rf_out2_ex_i_reg_6_ ( .D(dp_n787), .CK(CLK), .RN(dp_n41), .Q(
        dp_data_mem_ex_o[6]), .QN(dp_n457) );
  DFFR_X1 dp_rf_out2_ex_i_reg_5_ ( .D(dp_n786), .CK(CLK), .RN(dp_n41), .Q(
        dp_data_mem_ex_o[5]), .QN(dp_n456) );
  DFFR_X1 dp_rf_out2_ex_i_reg_4_ ( .D(dp_n785), .CK(CLK), .RN(dp_n41), .Q(
        dp_data_mem_ex_o[4]), .QN(dp_n455) );
  DFFR_X1 dp_rf_out2_ex_i_reg_3_ ( .D(dp_n784), .CK(CLK), .RN(dp_n41), .Q(
        dp_data_mem_ex_o[3]), .QN(dp_n454) );
  DFFR_X1 dp_rf_out2_ex_i_reg_2_ ( .D(dp_n783), .CK(CLK), .RN(dp_n41), .Q(
        dp_data_mem_ex_o[2]), .QN(dp_n453) );
  DFFR_X1 dp_rf_out2_ex_i_reg_1_ ( .D(dp_n782), .CK(CLK), .RN(dp_n41), .Q(
        dp_data_mem_ex_o[1]), .QN(dp_n452) );
  DFFR_X1 dp_rf_out2_ex_i_reg_0_ ( .D(dp_n781), .CK(CLK), .RN(dp_n41), .Q(
        dp_data_mem_ex_o[0]), .QN(dp_n451) );
  DFFR_X1 dp_imm_ex_i_reg_31_ ( .D(dp_n780), .CK(CLK), .RN(dp_n41), .Q(
        dp_imm_ex_i[31]), .QN(dp_n450) );
  DFFR_X1 dp_imm_ex_i_reg_30_ ( .D(dp_n779), .CK(CLK), .RN(dp_n41), .Q(
        dp_imm_ex_i[30]), .QN(dp_n449) );
  DFFR_X1 dp_imm_ex_i_reg_29_ ( .D(dp_n778), .CK(CLK), .RN(dp_n41), .Q(
        dp_imm_ex_i[29]), .QN(dp_n448) );
  DFFR_X1 dp_imm_ex_i_reg_28_ ( .D(dp_n777), .CK(CLK), .RN(dp_n41), .Q(
        dp_imm_ex_i[28]), .QN(dp_n447) );
  DFFR_X1 dp_imm_ex_i_reg_27_ ( .D(dp_n776), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[27]), .QN(dp_n446) );
  DFFR_X1 dp_imm_ex_i_reg_26_ ( .D(dp_n775), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[26]), .QN(dp_n445) );
  DFFR_X1 dp_imm_ex_i_reg_25_ ( .D(dp_n774), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[25]), .QN(dp_n444) );
  DFFR_X1 dp_imm_ex_i_reg_24_ ( .D(dp_n773), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[24]), .QN(dp_n443) );
  DFFR_X1 dp_imm_ex_i_reg_23_ ( .D(dp_n772), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[23]), .QN(dp_n442) );
  DFFR_X1 dp_imm_ex_i_reg_22_ ( .D(dp_n771), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[22]), .QN(dp_n441) );
  DFFR_X1 dp_imm_ex_i_reg_21_ ( .D(dp_n770), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[21]), .QN(dp_n440) );
  DFFR_X1 dp_imm_ex_i_reg_20_ ( .D(dp_n769), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[20]), .QN(dp_n439) );
  DFFR_X1 dp_imm_ex_i_reg_19_ ( .D(dp_n768), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[19]), .QN(dp_n438) );
  DFFR_X1 dp_imm_ex_i_reg_18_ ( .D(dp_n767), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[18]), .QN(dp_n437) );
  DFFR_X1 dp_imm_ex_i_reg_17_ ( .D(dp_n766), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[17]), .QN(dp_n436) );
  DFFR_X1 dp_imm_ex_i_reg_16_ ( .D(dp_n765), .CK(CLK), .RN(dp_n42), .Q(
        dp_imm_ex_i[16]), .QN(dp_n435) );
  DFFR_X1 dp_imm_ex_i_reg_15_ ( .D(dp_n764), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[15]), .QN(dp_n434) );
  DFFR_X1 dp_imm_ex_i_reg_14_ ( .D(dp_n763), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[14]), .QN(dp_n433) );
  DFFR_X1 dp_imm_ex_i_reg_13_ ( .D(dp_n762), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[13]), .QN(dp_n432) );
  DFFR_X1 dp_imm_ex_i_reg_12_ ( .D(dp_n761), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[12]), .QN(dp_n431) );
  DFFR_X1 dp_imm_ex_i_reg_11_ ( .D(dp_n760), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[11]), .QN(dp_n430) );
  DFFR_X1 dp_imm_ex_i_reg_10_ ( .D(dp_n759), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[10]), .QN(dp_n429) );
  DFFR_X1 dp_imm_ex_i_reg_9_ ( .D(dp_n758), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[9]), .QN(dp_n428) );
  DFFR_X1 dp_imm_ex_i_reg_8_ ( .D(dp_n757), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[8]), .QN(dp_n427) );
  DFFR_X1 dp_imm_ex_i_reg_7_ ( .D(dp_n756), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[7]), .QN(dp_n426) );
  DFFR_X1 dp_imm_ex_i_reg_6_ ( .D(dp_n755), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[6]), .QN(dp_n425) );
  DFFR_X1 dp_imm_ex_i_reg_5_ ( .D(dp_n754), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[5]), .QN(dp_n424) );
  DFFR_X1 dp_imm_ex_i_reg_4_ ( .D(dp_n753), .CK(CLK), .RN(dp_n43), .Q(
        dp_imm_ex_i[4]), .QN(dp_n423) );
  DFFR_X1 dp_imm_ex_i_reg_3_ ( .D(dp_n752), .CK(CLK), .RN(dp_n44), .Q(
        dp_imm_ex_i[3]), .QN(dp_n422) );
  DFFR_X1 dp_imm_ex_i_reg_2_ ( .D(dp_n751), .CK(CLK), .RN(dp_n44), .Q(
        dp_imm_ex_i[2]), .QN(dp_n421) );
  DFFR_X1 dp_imm_ex_i_reg_1_ ( .D(dp_n750), .CK(CLK), .RN(dp_n44), .Q(
        dp_imm_ex_i[1]), .QN(dp_n420) );
  DFFR_X1 dp_imm_ex_i_reg_0_ ( .D(dp_n749), .CK(CLK), .RN(dp_n44), .Q(
        dp_imm_ex_i[0]), .QN(dp_n419) );
  DFFR_X1 dp_rd_fwd_ex_i_reg_4_ ( .D(dp_n716), .CK(CLK), .RN(dp_n45), .Q(
        dp_rd_fwd_ex_o[4]), .QN(dp_n418) );
  DFFR_X1 dp_rd_fwd_ex_i_reg_3_ ( .D(dp_n715), .CK(CLK), .RN(dp_n45), .Q(
        dp_rd_fwd_ex_o[3]), .QN(dp_n417) );
  DFFR_X1 dp_rd_fwd_ex_i_reg_2_ ( .D(dp_n714), .CK(CLK), .RN(dp_n45), .Q(
        dp_rd_fwd_ex_o[2]), .QN(dp_n416) );
  DFFR_X1 dp_rd_fwd_ex_i_reg_1_ ( .D(dp_n713), .CK(CLK), .RN(dp_n45), .Q(
        dp_rd_fwd_ex_o[1]), .QN(dp_n415) );
  DFFR_X1 dp_rd_fwd_ex_i_reg_0_ ( .D(dp_n712), .CK(CLK), .RN(dp_n45), .Q(
        dp_rd_fwd_ex_o[0]), .QN(dp_n414) );
  INV_X1 dp_if_stage_U59 ( .A(RST), .ZN(dp_if_stage_n41) );
  MUX2_X1 dp_if_stage_U58 ( .A(IRAM_ADDRESS[16]), .B(dp_npc_if_o[16]), .S(
        dp_if_stage_n39), .Z(dp_if_stage_n16) );
  MUX2_X1 dp_if_stage_U57 ( .A(IRAM_ADDRESS[17]), .B(dp_npc_if_o[17]), .S(
        dp_if_stage_n39), .Z(dp_if_stage_n15) );
  MUX2_X1 dp_if_stage_U56 ( .A(IRAM_ADDRESS[18]), .B(dp_npc_if_o[18]), .S(
        dp_if_stage_n39), .Z(dp_if_stage_n14) );
  MUX2_X1 dp_if_stage_U55 ( .A(IRAM_ADDRESS[19]), .B(dp_npc_if_o[19]), .S(
        dp_if_stage_n39), .Z(dp_if_stage_n13) );
  MUX2_X1 dp_if_stage_U54 ( .A(IRAM_ADDRESS[20]), .B(dp_npc_if_o[20]), .S(
        dp_if_stage_n39), .Z(dp_if_stage_n12) );
  MUX2_X1 dp_if_stage_U53 ( .A(IRAM_ADDRESS[21]), .B(dp_npc_if_o[21]), .S(
        dp_if_stage_n39), .Z(dp_if_stage_n11) );
  MUX2_X1 dp_if_stage_U52 ( .A(IRAM_ADDRESS[22]), .B(dp_npc_if_o[22]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n10) );
  MUX2_X1 dp_if_stage_U51 ( .A(IRAM_ADDRESS[23]), .B(dp_npc_if_o[23]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n9) );
  MUX2_X1 dp_if_stage_U50 ( .A(IRAM_ADDRESS[24]), .B(dp_npc_if_o[24]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n8) );
  MUX2_X1 dp_if_stage_U49 ( .A(IRAM_ADDRESS[25]), .B(dp_npc_if_o[25]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n7) );
  MUX2_X1 dp_if_stage_U48 ( .A(IRAM_ADDRESS[26]), .B(dp_npc_if_o[26]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n6) );
  MUX2_X1 dp_if_stage_U47 ( .A(IRAM_ADDRESS[27]), .B(dp_npc_if_o[27]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n5) );
  MUX2_X1 dp_if_stage_U46 ( .A(IRAM_ADDRESS[28]), .B(dp_npc_if_o[28]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n4) );
  MUX2_X1 dp_if_stage_U45 ( .A(IRAM_ADDRESS[29]), .B(dp_npc_if_o[29]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n3) );
  MUX2_X1 dp_if_stage_U44 ( .A(IRAM_ADDRESS[30]), .B(dp_npc_if_o[30]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n2) );
  MUX2_X1 dp_if_stage_U43 ( .A(IRAM_ADDRESS[31]), .B(dp_npc_if_o[31]), .S(
        dp_if_stage_n40), .Z(dp_if_stage_n1) );
  NAND2_X1 dp_if_stage_U42 ( .A1(dp_npc_if_o[0]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n32) );
  OAI21_X1 dp_if_stage_U41 ( .B1(dp_if_stage_n64), .B2(dp_if_stage_n39), .A(
        dp_if_stage_n32), .ZN(dp_if_stage_n97) );
  NAND2_X1 dp_if_stage_U40 ( .A1(dp_npc_if_o[1]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n31) );
  OAI21_X1 dp_if_stage_U39 ( .B1(dp_if_stage_n63), .B2(dp_if_stage_n39), .A(
        dp_if_stage_n31), .ZN(dp_if_stage_n95) );
  NAND2_X1 dp_if_stage_U38 ( .A1(dp_npc_if_o[2]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n30) );
  OAI21_X1 dp_if_stage_U37 ( .B1(dp_if_stage_n62), .B2(dp_if_stage_n39), .A(
        dp_if_stage_n30), .ZN(dp_if_stage_n94) );
  NAND2_X1 dp_if_stage_U36 ( .A1(dp_npc_if_o[3]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n29) );
  OAI21_X1 dp_if_stage_U35 ( .B1(dp_if_stage_n61), .B2(dp_if_stage_n39), .A(
        dp_if_stage_n29), .ZN(dp_if_stage_n93) );
  NAND2_X1 dp_if_stage_U34 ( .A1(dp_npc_if_o[4]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n28) );
  OAI21_X1 dp_if_stage_U33 ( .B1(dp_if_stage_n60), .B2(dp_if_stage_n39), .A(
        dp_if_stage_n28), .ZN(dp_if_stage_n92) );
  NAND2_X1 dp_if_stage_U32 ( .A1(dp_npc_if_o[5]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n27) );
  OAI21_X1 dp_if_stage_U31 ( .B1(dp_if_stage_n59), .B2(dp_if_stage_n39), .A(
        dp_if_stage_n27), .ZN(dp_if_stage_n91) );
  NAND2_X1 dp_if_stage_U30 ( .A1(dp_npc_if_o[6]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n26) );
  OAI21_X1 dp_if_stage_U29 ( .B1(dp_if_stage_n58), .B2(dp_if_stage_n39), .A(
        dp_if_stage_n26), .ZN(dp_if_stage_n90) );
  NAND2_X1 dp_if_stage_U28 ( .A1(dp_npc_if_o[7]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n25) );
  OAI21_X1 dp_if_stage_U27 ( .B1(dp_if_stage_n57), .B2(dp_if_stage_n39), .A(
        dp_if_stage_n25), .ZN(dp_if_stage_n89) );
  NAND2_X1 dp_if_stage_U26 ( .A1(dp_npc_if_o[8]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n24) );
  OAI21_X1 dp_if_stage_U25 ( .B1(dp_if_stage_n56), .B2(dp_if_stage_n38), .A(
        dp_if_stage_n24), .ZN(dp_if_stage_n88) );
  NAND2_X1 dp_if_stage_U24 ( .A1(dp_npc_if_o[9]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n23) );
  OAI21_X1 dp_if_stage_U23 ( .B1(dp_if_stage_n55), .B2(dp_if_stage_n38), .A(
        dp_if_stage_n23), .ZN(dp_if_stage_n87) );
  NAND2_X1 dp_if_stage_U22 ( .A1(dp_npc_if_o[10]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n22) );
  OAI21_X1 dp_if_stage_U21 ( .B1(dp_if_stage_n54), .B2(dp_if_stage_n38), .A(
        dp_if_stage_n22), .ZN(dp_if_stage_n86) );
  NAND2_X1 dp_if_stage_U20 ( .A1(dp_npc_if_o[11]), .A2(dp_if_stage_n37), .ZN(
        dp_if_stage_n21) );
  OAI21_X1 dp_if_stage_U19 ( .B1(dp_if_stage_n53), .B2(dp_if_stage_n38), .A(
        dp_if_stage_n21), .ZN(dp_if_stage_n85) );
  NAND2_X1 dp_if_stage_U18 ( .A1(dp_npc_if_o[12]), .A2(dp_if_stage_n38), .ZN(
        dp_if_stage_n20) );
  OAI21_X1 dp_if_stage_U17 ( .B1(dp_if_stage_n52), .B2(dp_if_stage_n38), .A(
        dp_if_stage_n20), .ZN(dp_if_stage_n84) );
  NAND2_X1 dp_if_stage_U16 ( .A1(dp_npc_if_o[13]), .A2(dp_if_stage_n38), .ZN(
        dp_if_stage_n19) );
  OAI21_X1 dp_if_stage_U15 ( .B1(dp_if_stage_n51), .B2(dp_if_stage_n38), .A(
        dp_if_stage_n19), .ZN(dp_if_stage_n83) );
  NAND2_X1 dp_if_stage_U14 ( .A1(dp_npc_if_o[14]), .A2(dp_if_stage_n38), .ZN(
        dp_if_stage_n18) );
  OAI21_X1 dp_if_stage_U13 ( .B1(dp_if_stage_n50), .B2(dp_if_stage_n38), .A(
        dp_if_stage_n18), .ZN(dp_if_stage_n82) );
  NAND2_X1 dp_if_stage_U12 ( .A1(dp_npc_if_o[15]), .A2(dp_if_stage_n38), .ZN(
        dp_if_stage_n17) );
  OAI21_X1 dp_if_stage_U11 ( .B1(dp_if_stage_n49), .B2(dp_if_stage_n38), .A(
        dp_if_stage_n17), .ZN(dp_if_stage_n81) );
  BUF_X1 dp_if_stage_U10 ( .A(dp_if_stage_n41), .Z(dp_if_stage_n33) );
  BUF_X1 dp_if_stage_U9 ( .A(dp_if_stage_n41), .Z(dp_if_stage_n34) );
  BUF_X1 dp_if_stage_U8 ( .A(dp_if_stage_n36), .Z(dp_if_stage_n40) );
  BUF_X1 dp_if_stage_U7 ( .A(dp_if_stage_n36), .Z(dp_if_stage_n39) );
  BUF_X1 dp_if_stage_U6 ( .A(dp_if_stage_n35), .Z(dp_if_stage_n38) );
  BUF_X1 dp_if_stage_U5 ( .A(dp_if_stage_n35), .Z(dp_if_stage_n37) );
  CLKBUF_X1 dp_if_stage_U4 ( .A(pipe_ex_mem_en_i), .Z(dp_if_stage_n35) );
  CLKBUF_X1 dp_if_stage_U3 ( .A(pipe_ex_mem_en_i), .Z(dp_if_stage_n36) );
  DFFR_X1 dp_if_stage_PC_i_reg_16_ ( .D(dp_if_stage_n16), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[16]) );
  DFFR_X1 dp_if_stage_PC_i_reg_17_ ( .D(dp_if_stage_n15), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[17]) );
  DFFR_X1 dp_if_stage_PC_i_reg_18_ ( .D(dp_if_stage_n14), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[18]) );
  DFFR_X1 dp_if_stage_PC_i_reg_19_ ( .D(dp_if_stage_n13), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[19]) );
  DFFR_X1 dp_if_stage_PC_i_reg_20_ ( .D(dp_if_stage_n12), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[20]) );
  DFFR_X1 dp_if_stage_PC_i_reg_21_ ( .D(dp_if_stage_n11), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[21]) );
  DFFR_X1 dp_if_stage_PC_i_reg_22_ ( .D(dp_if_stage_n10), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[22]) );
  DFFR_X1 dp_if_stage_PC_i_reg_23_ ( .D(dp_if_stage_n9), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[23]) );
  DFFR_X1 dp_if_stage_PC_i_reg_24_ ( .D(dp_if_stage_n8), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[24]) );
  DFFR_X1 dp_if_stage_PC_i_reg_25_ ( .D(dp_if_stage_n7), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[25]) );
  DFFR_X1 dp_if_stage_PC_i_reg_26_ ( .D(dp_if_stage_n6), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[26]) );
  DFFR_X1 dp_if_stage_PC_i_reg_27_ ( .D(dp_if_stage_n5), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[27]) );
  DFFR_X1 dp_if_stage_PC_i_reg_28_ ( .D(dp_if_stage_n4), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[28]) );
  DFFR_X1 dp_if_stage_PC_i_reg_29_ ( .D(dp_if_stage_n3), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[29]) );
  DFFR_X1 dp_if_stage_PC_i_reg_30_ ( .D(dp_if_stage_n2), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[30]) );
  DFFR_X1 dp_if_stage_PC_i_reg_31_ ( .D(dp_if_stage_n1), .CK(CLK), .RN(
        dp_if_stage_n41), .Q(IRAM_ADDRESS[31]) );
  DFFR_X1 dp_if_stage_PC_i_reg_15_ ( .D(dp_if_stage_n81), .CK(CLK), .RN(
        dp_if_stage_n34), .Q(IRAM_ADDRESS[15]), .QN(dp_if_stage_n49) );
  DFFR_X1 dp_if_stage_PC_i_reg_14_ ( .D(dp_if_stage_n82), .CK(CLK), .RN(
        dp_if_stage_n34), .Q(IRAM_ADDRESS[14]), .QN(dp_if_stage_n50) );
  DFFR_X1 dp_if_stage_PC_i_reg_13_ ( .D(dp_if_stage_n83), .CK(CLK), .RN(
        dp_if_stage_n34), .Q(IRAM_ADDRESS[13]), .QN(dp_if_stage_n51) );
  DFFR_X1 dp_if_stage_PC_i_reg_12_ ( .D(dp_if_stage_n84), .CK(CLK), .RN(
        dp_if_stage_n34), .Q(IRAM_ADDRESS[12]), .QN(dp_if_stage_n52) );
  DFFR_X1 dp_if_stage_PC_i_reg_11_ ( .D(dp_if_stage_n85), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[11]), .QN(dp_if_stage_n53) );
  DFFR_X1 dp_if_stage_PC_i_reg_10_ ( .D(dp_if_stage_n86), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[10]), .QN(dp_if_stage_n54) );
  DFFR_X1 dp_if_stage_PC_i_reg_9_ ( .D(dp_if_stage_n87), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[9]), .QN(dp_if_stage_n55) );
  DFFR_X1 dp_if_stage_PC_i_reg_8_ ( .D(dp_if_stage_n88), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[8]), .QN(dp_if_stage_n56) );
  DFFR_X1 dp_if_stage_PC_i_reg_7_ ( .D(dp_if_stage_n89), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[7]), .QN(dp_if_stage_n57) );
  DFFR_X1 dp_if_stage_PC_i_reg_6_ ( .D(dp_if_stage_n90), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[6]), .QN(dp_if_stage_n58) );
  DFFR_X1 dp_if_stage_PC_i_reg_5_ ( .D(dp_if_stage_n91), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[5]), .QN(dp_if_stage_n59) );
  DFFR_X1 dp_if_stage_PC_i_reg_4_ ( .D(dp_if_stage_n92), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[4]), .QN(dp_if_stage_n60) );
  DFFR_X1 dp_if_stage_PC_i_reg_3_ ( .D(dp_if_stage_n93), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[3]), .QN(dp_if_stage_n61) );
  DFFR_X1 dp_if_stage_PC_i_reg_2_ ( .D(dp_if_stage_n94), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[2]), .QN(dp_if_stage_n62) );
  DFFR_X1 dp_if_stage_PC_i_reg_1_ ( .D(dp_if_stage_n95), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[1]), .QN(dp_if_stage_n63) );
  DFFR_X1 dp_if_stage_PC_i_reg_0_ ( .D(dp_if_stage_n97), .CK(CLK), .RN(
        dp_if_stage_n33), .Q(IRAM_ADDRESS[0]), .QN(dp_if_stage_n64) );
  MUX2_X1 dp_if_stage_mux_U55 ( .A(dp_if_stage_NPC_4_i_31_), .B(
        DRAM_ADDRESS[31]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[31]) );
  MUX2_X1 dp_if_stage_mux_U54 ( .A(dp_if_stage_NPC_4_i_30_), .B(
        DRAM_ADDRESS[30]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[30]) );
  MUX2_X1 dp_if_stage_mux_U53 ( .A(dp_if_stage_NPC_4_i_29_), .B(
        DRAM_ADDRESS[29]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[29]) );
  MUX2_X1 dp_if_stage_mux_U52 ( .A(dp_if_stage_NPC_4_i_28_), .B(
        DRAM_ADDRESS[28]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[28]) );
  MUX2_X1 dp_if_stage_mux_U51 ( .A(dp_if_stage_NPC_4_i_27_), .B(
        DRAM_ADDRESS[27]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[27]) );
  MUX2_X1 dp_if_stage_mux_U50 ( .A(dp_if_stage_NPC_4_i_26_), .B(
        DRAM_ADDRESS[26]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[26]) );
  MUX2_X1 dp_if_stage_mux_U49 ( .A(dp_if_stage_NPC_4_i_25_), .B(
        DRAM_ADDRESS[25]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[25]) );
  MUX2_X1 dp_if_stage_mux_U48 ( .A(dp_if_stage_NPC_4_i_24_), .B(
        DRAM_ADDRESS[24]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[24]) );
  MUX2_X1 dp_if_stage_mux_U47 ( .A(dp_if_stage_NPC_4_i_23_), .B(
        DRAM_ADDRESS[23]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[23]) );
  MUX2_X1 dp_if_stage_mux_U46 ( .A(dp_if_stage_NPC_4_i_22_), .B(
        DRAM_ADDRESS[22]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[22]) );
  MUX2_X1 dp_if_stage_mux_U45 ( .A(dp_if_stage_NPC_4_i_21_), .B(
        DRAM_ADDRESS[21]), .S(jump_en_i), .Z(dp_npc_if_o[21]) );
  MUX2_X1 dp_if_stage_mux_U44 ( .A(dp_if_stage_NPC_4_i_20_), .B(
        DRAM_ADDRESS[20]), .S(jump_en_i), .Z(dp_npc_if_o[20]) );
  MUX2_X1 dp_if_stage_mux_U43 ( .A(dp_if_stage_NPC_4_i_19_), .B(
        DRAM_ADDRESS[19]), .S(jump_en_i), .Z(dp_npc_if_o[19]) );
  MUX2_X1 dp_if_stage_mux_U42 ( .A(dp_if_stage_NPC_4_i_18_), .B(
        DRAM_ADDRESS[18]), .S(jump_en_i), .Z(dp_npc_if_o[18]) );
  MUX2_X1 dp_if_stage_mux_U41 ( .A(dp_if_stage_NPC_4_i_17_), .B(
        DRAM_ADDRESS[17]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[17]) );
  MUX2_X1 dp_if_stage_mux_U40 ( .A(dp_if_stage_NPC_4_i_16_), .B(
        DRAM_ADDRESS[16]), .S(dp_if_stage_mux_n1), .Z(dp_npc_if_o[16]) );
  INV_X1 dp_if_stage_mux_U39 ( .A(jump_en_i), .ZN(dp_if_stage_mux_n7) );
  AOI22_X1 dp_if_stage_mux_U38 ( .A1(IRAM_ADDRESS[1]), .A2(dp_if_stage_mux_n3), 
        .B1(DRAM_ADDRESS[1]), .B2(jump_en_i), .ZN(dp_if_stage_mux_n54) );
  INV_X1 dp_if_stage_mux_U37 ( .A(dp_if_stage_mux_n54), .ZN(dp_npc_if_o[1]) );
  AOI22_X1 dp_if_stage_mux_U36 ( .A1(dp_if_stage_NPC_4_i_2_), .A2(
        dp_if_stage_mux_n4), .B1(DRAM_ADDRESS[2]), .B2(jump_en_i), .ZN(
        dp_if_stage_mux_n43) );
  INV_X1 dp_if_stage_mux_U35 ( .A(dp_if_stage_mux_n43), .ZN(dp_npc_if_o[2]) );
  AOI22_X1 dp_if_stage_mux_U34 ( .A1(dp_if_stage_NPC_4_i_3_), .A2(
        dp_if_stage_mux_n4), .B1(DRAM_ADDRESS[3]), .B2(dp_if_stage_mux_n1), 
        .ZN(dp_if_stage_mux_n40) );
  INV_X1 dp_if_stage_mux_U33 ( .A(dp_if_stage_mux_n40), .ZN(dp_npc_if_o[3]) );
  AOI22_X1 dp_if_stage_mux_U32 ( .A1(dp_if_stage_NPC_4_i_4_), .A2(
        dp_if_stage_mux_n4), .B1(DRAM_ADDRESS[4]), .B2(dp_if_stage_mux_n1), 
        .ZN(dp_if_stage_mux_n39) );
  INV_X1 dp_if_stage_mux_U31 ( .A(dp_if_stage_mux_n39), .ZN(dp_npc_if_o[4]) );
  AOI22_X1 dp_if_stage_mux_U30 ( .A1(dp_if_stage_NPC_4_i_5_), .A2(
        dp_if_stage_mux_n4), .B1(DRAM_ADDRESS[5]), .B2(dp_if_stage_mux_n1), 
        .ZN(dp_if_stage_mux_n38) );
  INV_X1 dp_if_stage_mux_U29 ( .A(dp_if_stage_mux_n38), .ZN(dp_npc_if_o[5]) );
  AOI22_X1 dp_if_stage_mux_U28 ( .A1(dp_if_stage_NPC_4_i_6_), .A2(
        dp_if_stage_mux_n5), .B1(DRAM_ADDRESS[6]), .B2(dp_if_stage_mux_n1), 
        .ZN(dp_if_stage_mux_n37) );
  INV_X1 dp_if_stage_mux_U27 ( .A(dp_if_stage_mux_n37), .ZN(dp_npc_if_o[6]) );
  AOI22_X1 dp_if_stage_mux_U26 ( .A1(dp_if_stage_NPC_4_i_8_), .A2(
        dp_if_stage_mux_n5), .B1(DRAM_ADDRESS[8]), .B2(jump_en_i), .ZN(
        dp_if_stage_mux_n35) );
  INV_X1 dp_if_stage_mux_U25 ( .A(dp_if_stage_mux_n35), .ZN(dp_npc_if_o[8]) );
  AOI22_X1 dp_if_stage_mux_U24 ( .A1(dp_if_stage_NPC_4_i_12_), .A2(
        dp_if_stage_mux_n2), .B1(DRAM_ADDRESS[12]), .B2(jump_en_i), .ZN(
        dp_if_stage_mux_n62) );
  INV_X1 dp_if_stage_mux_U23 ( .A(dp_if_stage_mux_n62), .ZN(dp_npc_if_o[12])
         );
  AOI22_X1 dp_if_stage_mux_U22 ( .A1(dp_if_stage_NPC_4_i_13_), .A2(
        dp_if_stage_mux_n3), .B1(DRAM_ADDRESS[13]), .B2(jump_en_i), .ZN(
        dp_if_stage_mux_n61) );
  INV_X1 dp_if_stage_mux_U21 ( .A(dp_if_stage_mux_n61), .ZN(dp_npc_if_o[13])
         );
  AOI22_X1 dp_if_stage_mux_U20 ( .A1(dp_if_stage_NPC_4_i_14_), .A2(
        dp_if_stage_mux_n3), .B1(DRAM_ADDRESS[14]), .B2(jump_en_i), .ZN(
        dp_if_stage_mux_n60) );
  INV_X1 dp_if_stage_mux_U19 ( .A(dp_if_stage_mux_n60), .ZN(dp_npc_if_o[14])
         );
  AOI22_X1 dp_if_stage_mux_U18 ( .A1(dp_if_stage_NPC_4_i_15_), .A2(
        dp_if_stage_mux_n3), .B1(DRAM_ADDRESS[15]), .B2(jump_en_i), .ZN(
        dp_if_stage_mux_n59) );
  INV_X1 dp_if_stage_mux_U17 ( .A(dp_if_stage_mux_n59), .ZN(dp_npc_if_o[15])
         );
  AOI22_X1 dp_if_stage_mux_U16 ( .A1(IRAM_ADDRESS[0]), .A2(dp_if_stage_mux_n2), 
        .B1(DRAM_ADDRESS[0]), .B2(dp_if_stage_mux_n1), .ZN(dp_if_stage_mux_n65) );
  INV_X1 dp_if_stage_mux_U15 ( .A(dp_if_stage_mux_n65), .ZN(dp_npc_if_o[0]) );
  AOI22_X1 dp_if_stage_mux_U14 ( .A1(dp_if_stage_NPC_4_i_10_), .A2(
        dp_if_stage_mux_n2), .B1(DRAM_ADDRESS[10]), .B2(dp_if_stage_mux_n1), 
        .ZN(dp_if_stage_mux_n64) );
  INV_X1 dp_if_stage_mux_U13 ( .A(dp_if_stage_mux_n64), .ZN(dp_npc_if_o[10])
         );
  AOI22_X1 dp_if_stage_mux_U12 ( .A1(dp_if_stage_NPC_4_i_11_), .A2(
        dp_if_stage_mux_n2), .B1(DRAM_ADDRESS[11]), .B2(dp_if_stage_mux_n1), 
        .ZN(dp_if_stage_mux_n63) );
  INV_X1 dp_if_stage_mux_U11 ( .A(dp_if_stage_mux_n63), .ZN(dp_npc_if_o[11])
         );
  AOI22_X1 dp_if_stage_mux_U10 ( .A1(dp_if_stage_NPC_4_i_9_), .A2(
        dp_if_stage_mux_n5), .B1(dp_if_stage_mux_n1), .B2(DRAM_ADDRESS[9]), 
        .ZN(dp_if_stage_mux_n34) );
  INV_X1 dp_if_stage_mux_U9 ( .A(dp_if_stage_mux_n34), .ZN(dp_npc_if_o[9]) );
  AOI22_X1 dp_if_stage_mux_U8 ( .A1(dp_if_stage_NPC_4_i_7_), .A2(
        dp_if_stage_mux_n5), .B1(DRAM_ADDRESS[7]), .B2(dp_if_stage_mux_n1), 
        .ZN(dp_if_stage_mux_n36) );
  INV_X1 dp_if_stage_mux_U7 ( .A(dp_if_stage_mux_n36), .ZN(dp_npc_if_o[7]) );
  BUF_X1 dp_if_stage_mux_U6 ( .A(dp_if_stage_mux_n7), .Z(dp_if_stage_mux_n6)
         );
  BUF_X1 dp_if_stage_mux_U5 ( .A(dp_if_stage_mux_n7), .Z(dp_if_stage_mux_n2)
         );
  BUF_X1 dp_if_stage_mux_U4 ( .A(dp_if_stage_mux_n7), .Z(dp_if_stage_mux_n3)
         );
  BUF_X1 dp_if_stage_mux_U3 ( .A(dp_if_stage_mux_n7), .Z(dp_if_stage_mux_n4)
         );
  BUF_X1 dp_if_stage_mux_U2 ( .A(dp_if_stage_mux_n7), .Z(dp_if_stage_mux_n5)
         );
  INV_X1 dp_if_stage_mux_U1 ( .A(dp_if_stage_mux_n6), .ZN(dp_if_stage_mux_n1)
         );
  XNOR2_X1 dp_if_stage_add_77_U91 ( .A(dp_if_stage_add_77_n58), .B(
        dp_if_stage_add_77_n56), .ZN(dp_if_stage_NPC_4_i_10_) );
  XNOR2_X1 dp_if_stage_add_77_U90 ( .A(dp_if_stage_add_77_n57), .B(
        dp_if_stage_add_77_n55), .ZN(dp_if_stage_NPC_4_i_11_) );
  INV_X1 dp_if_stage_add_77_U89 ( .A(dp_if_stage_add_77_n11), .ZN(
        dp_if_stage_add_77_n54) );
  XNOR2_X1 dp_if_stage_add_77_U88 ( .A(dp_if_stage_add_77_n52), .B(
        dp_if_stage_add_77_n51), .ZN(dp_if_stage_NPC_4_i_13_) );
  XNOR2_X1 dp_if_stage_add_77_U87 ( .A(dp_if_stage_add_77_n50), .B(
        dp_if_stage_add_77_n48), .ZN(dp_if_stage_NPC_4_i_15_) );
  INV_X1 dp_if_stage_add_77_U86 ( .A(dp_if_stage_add_77_n47), .ZN(
        dp_if_stage_add_77_n44) );
  NAND3_X1 dp_if_stage_add_77_U85 ( .A1(IRAM_ADDRESS[18]), .A2(
        IRAM_ADDRESS[19]), .A3(IRAM_ADDRESS[17]), .ZN(dp_if_stage_add_77_n38)
         );
  NAND3_X1 dp_if_stage_add_77_U84 ( .A1(IRAM_ADDRESS[22]), .A2(
        IRAM_ADDRESS[23]), .A3(IRAM_ADDRESS[21]), .ZN(dp_if_stage_add_77_n32)
         );
  NAND3_X1 dp_if_stage_add_77_U83 ( .A1(IRAM_ADDRESS[26]), .A2(
        IRAM_ADDRESS[27]), .A3(IRAM_ADDRESS[25]), .ZN(dp_if_stage_add_77_n26)
         );
  XNOR2_X1 dp_if_stage_add_77_U82 ( .A(dp_if_stage_add_77_n14), .B(
        dp_if_stage_add_77_n13), .ZN(dp_if_stage_NPC_4_i_5_) );
  XNOR2_X1 dp_if_stage_add_77_U81 ( .A(dp_if_stage_add_77_n59), .B(
        dp_if_stage_add_77_n11), .ZN(dp_if_stage_NPC_4_i_8_) );
  XNOR2_X1 dp_if_stage_add_77_U80 ( .A(dp_if_stage_add_77_n10), .B(
        IRAM_ADDRESS[9]), .ZN(dp_if_stage_NPC_4_i_9_) );
  INV_X1 dp_if_stage_add_77_U79 ( .A(IRAM_ADDRESS[31]), .ZN(
        dp_if_stage_add_77_n18) );
  INV_X1 dp_if_stage_add_77_U78 ( .A(IRAM_ADDRESS[9]), .ZN(
        dp_if_stage_add_77_n61) );
  INV_X1 dp_if_stage_add_77_U77 ( .A(IRAM_ADDRESS[19]), .ZN(
        dp_if_stage_add_77_n39) );
  INV_X1 dp_if_stage_add_77_U76 ( .A(IRAM_ADDRESS[23]), .ZN(
        dp_if_stage_add_77_n33) );
  INV_X1 dp_if_stage_add_77_U75 ( .A(IRAM_ADDRESS[27]), .ZN(
        dp_if_stage_add_77_n27) );
  INV_X1 dp_if_stage_add_77_U74 ( .A(IRAM_ADDRESS[29]), .ZN(
        dp_if_stage_add_77_n23) );
  INV_X1 dp_if_stage_add_77_U73 ( .A(IRAM_ADDRESS[11]), .ZN(
        dp_if_stage_add_77_n57) );
  INV_X1 dp_if_stage_add_77_U72 ( .A(IRAM_ADDRESS[30]), .ZN(
        dp_if_stage_add_77_n20) );
  INV_X1 dp_if_stage_add_77_U71 ( .A(IRAM_ADDRESS[28]), .ZN(
        dp_if_stage_add_77_n24) );
  INV_X1 dp_if_stage_add_77_U70 ( .A(IRAM_ADDRESS[20]), .ZN(
        dp_if_stage_add_77_n36) );
  INV_X1 dp_if_stage_add_77_U69 ( .A(IRAM_ADDRESS[24]), .ZN(
        dp_if_stage_add_77_n30) );
  INV_X1 dp_if_stage_add_77_U68 ( .A(IRAM_ADDRESS[5]), .ZN(
        dp_if_stage_add_77_n14) );
  INV_X1 dp_if_stage_add_77_U67 ( .A(IRAM_ADDRESS[13]), .ZN(
        dp_if_stage_add_77_n52) );
  INV_X1 dp_if_stage_add_77_U66 ( .A(IRAM_ADDRESS[15]), .ZN(
        dp_if_stage_add_77_n50) );
  INV_X1 dp_if_stage_add_77_U65 ( .A(IRAM_ADDRESS[10]), .ZN(
        dp_if_stage_add_77_n58) );
  INV_X1 dp_if_stage_add_77_U64 ( .A(IRAM_ADDRESS[4]), .ZN(
        dp_if_stage_add_77_n60) );
  XNOR2_X1 dp_if_stage_add_77_U63 ( .A(dp_if_stage_add_77_n35), .B(
        dp_if_stage_add_77_n36), .ZN(dp_if_stage_NPC_4_i_20_) );
  XNOR2_X1 dp_if_stage_add_77_U62 ( .A(dp_if_stage_add_77_n29), .B(
        dp_if_stage_add_77_n30), .ZN(dp_if_stage_NPC_4_i_24_) );
  XNOR2_X1 dp_if_stage_add_77_U61 ( .A(dp_if_stage_add_77_n22), .B(
        dp_if_stage_add_77_n24), .ZN(dp_if_stage_NPC_4_i_28_) );
  XNOR2_X1 dp_if_stage_add_77_U60 ( .A(dp_if_stage_add_77_n19), .B(
        dp_if_stage_add_77_n20), .ZN(dp_if_stage_NPC_4_i_30_) );
  XOR2_X1 dp_if_stage_add_77_U59 ( .A(dp_if_stage_add_77_n7), .B(
        IRAM_ADDRESS[18]), .Z(dp_if_stage_NPC_4_i_18_) );
  AND2_X1 dp_if_stage_add_77_U58 ( .A1(IRAM_ADDRESS[18]), .A2(
        dp_if_stage_add_77_n7), .ZN(dp_if_stage_add_77_n9) );
  XNOR2_X1 dp_if_stage_add_77_U57 ( .A(dp_if_stage_add_77_n9), .B(
        dp_if_stage_add_77_n39), .ZN(dp_if_stage_NPC_4_i_19_) );
  XOR2_X1 dp_if_stage_add_77_U56 ( .A(IRAM_ADDRESS[21]), .B(
        dp_if_stage_add_77_n34), .Z(dp_if_stage_NPC_4_i_21_) );
  XOR2_X1 dp_if_stage_add_77_U55 ( .A(IRAM_ADDRESS[16]), .B(
        dp_if_stage_add_77_n41), .Z(dp_if_stage_NPC_4_i_16_) );
  XOR2_X1 dp_if_stage_add_77_U54 ( .A(IRAM_ADDRESS[17]), .B(
        dp_if_stage_add_77_n40), .Z(dp_if_stage_NPC_4_i_17_) );
  XOR2_X1 dp_if_stage_add_77_U53 ( .A(dp_if_stage_add_77_n6), .B(
        IRAM_ADDRESS[22]), .Z(dp_if_stage_NPC_4_i_22_) );
  XOR2_X1 dp_if_stage_add_77_U52 ( .A(IRAM_ADDRESS[25]), .B(
        dp_if_stage_add_77_n28), .Z(dp_if_stage_NPC_4_i_25_) );
  XOR2_X1 dp_if_stage_add_77_U51 ( .A(dp_if_stage_add_77_n5), .B(
        IRAM_ADDRESS[26]), .Z(dp_if_stage_NPC_4_i_26_) );
  XNOR2_X1 dp_if_stage_add_77_U50 ( .A(IRAM_ADDRESS[29]), .B(
        dp_if_stage_add_77_n21), .ZN(dp_if_stage_NPC_4_i_29_) );
  INV_X1 dp_if_stage_add_77_U49 ( .A(IRAM_ADDRESS[2]), .ZN(
        dp_if_stage_NPC_4_i_2_) );
  INV_X1 dp_if_stage_add_77_U48 ( .A(IRAM_ADDRESS[8]), .ZN(
        dp_if_stage_add_77_n59) );
  INV_X1 dp_if_stage_add_77_U47 ( .A(IRAM_ADDRESS[3]), .ZN(
        dp_if_stage_add_77_n16) );
  AND2_X1 dp_if_stage_add_77_U46 ( .A1(IRAM_ADDRESS[6]), .A2(
        dp_if_stage_add_77_n12), .ZN(dp_if_stage_add_77_n8) );
  AND2_X1 dp_if_stage_add_77_U45 ( .A1(IRAM_ADDRESS[17]), .A2(
        dp_if_stage_add_77_n40), .ZN(dp_if_stage_add_77_n7) );
  AND2_X1 dp_if_stage_add_77_U44 ( .A1(IRAM_ADDRESS[21]), .A2(
        dp_if_stage_add_77_n34), .ZN(dp_if_stage_add_77_n6) );
  AND2_X1 dp_if_stage_add_77_U43 ( .A1(IRAM_ADDRESS[25]), .A2(
        dp_if_stage_add_77_n28), .ZN(dp_if_stage_add_77_n5) );
  NAND2_X1 dp_if_stage_add_77_U42 ( .A1(dp_if_stage_add_77_n11), .A2(
        IRAM_ADDRESS[8]), .ZN(dp_if_stage_add_77_n10) );
  NAND2_X1 dp_if_stage_add_77_U41 ( .A1(dp_if_stage_add_77_n29), .A2(
        IRAM_ADDRESS[24]), .ZN(dp_if_stage_add_77_n25) );
  NAND2_X1 dp_if_stage_add_77_U40 ( .A1(dp_if_stage_add_77_n35), .A2(
        IRAM_ADDRESS[20]), .ZN(dp_if_stage_add_77_n31) );
  NAND2_X1 dp_if_stage_add_77_U39 ( .A1(dp_if_stage_add_77_n41), .A2(
        IRAM_ADDRESS[16]), .ZN(dp_if_stage_add_77_n37) );
  NAND2_X1 dp_if_stage_add_77_U38 ( .A1(dp_if_stage_add_77_n22), .A2(
        IRAM_ADDRESS[28]), .ZN(dp_if_stage_add_77_n21) );
  AND2_X1 dp_if_stage_add_77_U37 ( .A1(dp_if_stage_add_77_n56), .A2(
        IRAM_ADDRESS[10]), .ZN(dp_if_stage_add_77_n55) );
  AND2_X1 dp_if_stage_add_77_U36 ( .A1(dp_if_stage_add_77_n49), .A2(
        IRAM_ADDRESS[14]), .ZN(dp_if_stage_add_77_n48) );
  OR2_X1 dp_if_stage_add_77_U35 ( .A1(dp_if_stage_NPC_4_i_2_), .A2(
        dp_if_stage_add_77_n16), .ZN(dp_if_stage_add_77_n4) );
  NOR2_X1 dp_if_stage_add_77_U34 ( .A1(dp_if_stage_add_77_n60), .A2(
        dp_if_stage_add_77_n4), .ZN(dp_if_stage_add_77_n13) );
  AND2_X1 dp_if_stage_add_77_U33 ( .A1(IRAM_ADDRESS[12]), .A2(
        dp_if_stage_add_77_n53), .ZN(dp_if_stage_add_77_n51) );
  NOR2_X1 dp_if_stage_add_77_U32 ( .A1(dp_if_stage_add_77_n23), .A2(
        dp_if_stage_add_77_n21), .ZN(dp_if_stage_add_77_n19) );
  NOR2_X1 dp_if_stage_add_77_U31 ( .A1(dp_if_stage_add_77_n25), .A2(
        dp_if_stage_add_77_n26), .ZN(dp_if_stage_add_77_n22) );
  NOR2_X1 dp_if_stage_add_77_U30 ( .A1(dp_if_stage_add_77_n31), .A2(
        dp_if_stage_add_77_n32), .ZN(dp_if_stage_add_77_n29) );
  NOR2_X1 dp_if_stage_add_77_U29 ( .A1(dp_if_stage_add_77_n37), .A2(
        dp_if_stage_add_77_n38), .ZN(dp_if_stage_add_77_n35) );
  NAND4_X1 dp_if_stage_add_77_U28 ( .A1(IRAM_ADDRESS[11]), .A2(
        IRAM_ADDRESS[10]), .A3(IRAM_ADDRESS[9]), .A4(IRAM_ADDRESS[8]), .ZN(
        dp_if_stage_add_77_n47) );
  NAND2_X1 dp_if_stage_add_77_U27 ( .A1(dp_if_stage_add_77_n44), .A2(
        dp_if_stage_add_77_n45), .ZN(dp_if_stage_add_77_n42) );
  NAND4_X1 dp_if_stage_add_77_U26 ( .A1(IRAM_ADDRESS[12]), .A2(
        IRAM_ADDRESS[13]), .A3(IRAM_ADDRESS[14]), .A4(IRAM_ADDRESS[15]), .ZN(
        dp_if_stage_add_77_n43) );
  NOR2_X1 dp_if_stage_add_77_U25 ( .A1(dp_if_stage_add_77_n42), .A2(
        dp_if_stage_add_77_n43), .ZN(dp_if_stage_add_77_n41) );
  NAND4_X1 dp_if_stage_add_77_U24 ( .A1(IRAM_ADDRESS[4]), .A2(IRAM_ADDRESS[5]), 
        .A3(IRAM_ADDRESS[6]), .A4(IRAM_ADDRESS[7]), .ZN(dp_if_stage_add_77_n46) );
  AND2_X1 dp_if_stage_add_77_U23 ( .A1(dp_if_stage_add_77_n51), .A2(
        IRAM_ADDRESS[13]), .ZN(dp_if_stage_add_77_n49) );
  AND2_X1 dp_if_stage_add_77_U22 ( .A1(dp_if_stage_add_77_n13), .A2(
        IRAM_ADDRESS[5]), .ZN(dp_if_stage_add_77_n12) );
  INV_X1 dp_if_stage_add_77_U21 ( .A(dp_if_stage_add_77_n4), .ZN(
        dp_if_stage_add_77_n15) );
  INV_X1 dp_if_stage_add_77_U20 ( .A(dp_if_stage_add_77_n31), .ZN(
        dp_if_stage_add_77_n34) );
  INV_X1 dp_if_stage_add_77_U19 ( .A(dp_if_stage_add_77_n25), .ZN(
        dp_if_stage_add_77_n28) );
  INV_X1 dp_if_stage_add_77_U18 ( .A(dp_if_stage_add_77_n37), .ZN(
        dp_if_stage_add_77_n40) );
  NOR2_X1 dp_if_stage_add_77_U17 ( .A1(dp_if_stage_add_77_n4), .A2(
        dp_if_stage_add_77_n46), .ZN(dp_if_stage_add_77_n45) );
  NOR2_X1 dp_if_stage_add_77_U16 ( .A1(dp_if_stage_add_77_n61), .A2(
        dp_if_stage_add_77_n10), .ZN(dp_if_stage_add_77_n56) );
  NOR2_X1 dp_if_stage_add_77_U15 ( .A1(dp_if_stage_add_77_n54), .A2(
        dp_if_stage_add_77_n47), .ZN(dp_if_stage_add_77_n53) );
  NOR2_X1 dp_if_stage_add_77_U14 ( .A1(dp_if_stage_add_77_n4), .A2(
        dp_if_stage_add_77_n46), .ZN(dp_if_stage_add_77_n11) );
  XOR2_X1 dp_if_stage_add_77_U13 ( .A(dp_if_stage_add_77_n16), .B(
        dp_if_stage_NPC_4_i_2_), .Z(dp_if_stage_NPC_4_i_3_) );
  XOR2_X1 dp_if_stage_add_77_U12 ( .A(IRAM_ADDRESS[4]), .B(
        dp_if_stage_add_77_n15), .Z(dp_if_stage_NPC_4_i_4_) );
  XOR2_X1 dp_if_stage_add_77_U11 ( .A(IRAM_ADDRESS[6]), .B(
        dp_if_stage_add_77_n12), .Z(dp_if_stage_NPC_4_i_6_) );
  XOR2_X1 dp_if_stage_add_77_U10 ( .A(IRAM_ADDRESS[7]), .B(
        dp_if_stage_add_77_n8), .Z(dp_if_stage_NPC_4_i_7_) );
  XOR2_X1 dp_if_stage_add_77_U9 ( .A(IRAM_ADDRESS[12]), .B(
        dp_if_stage_add_77_n53), .Z(dp_if_stage_NPC_4_i_12_) );
  XOR2_X1 dp_if_stage_add_77_U8 ( .A(IRAM_ADDRESS[14]), .B(
        dp_if_stage_add_77_n49), .Z(dp_if_stage_NPC_4_i_14_) );
  NAND2_X1 dp_if_stage_add_77_U7 ( .A1(IRAM_ADDRESS[22]), .A2(
        dp_if_stage_add_77_n6), .ZN(dp_if_stage_add_77_n3) );
  XOR2_X1 dp_if_stage_add_77_U6 ( .A(dp_if_stage_add_77_n3), .B(
        dp_if_stage_add_77_n33), .Z(dp_if_stage_NPC_4_i_23_) );
  NAND2_X1 dp_if_stage_add_77_U5 ( .A1(IRAM_ADDRESS[26]), .A2(
        dp_if_stage_add_77_n5), .ZN(dp_if_stage_add_77_n2) );
  XOR2_X1 dp_if_stage_add_77_U4 ( .A(dp_if_stage_add_77_n2), .B(
        dp_if_stage_add_77_n27), .Z(dp_if_stage_NPC_4_i_27_) );
  NAND2_X1 dp_if_stage_add_77_U3 ( .A1(dp_if_stage_add_77_n19), .A2(
        IRAM_ADDRESS[30]), .ZN(dp_if_stage_add_77_n1) );
  XOR2_X1 dp_if_stage_add_77_U2 ( .A(dp_if_stage_add_77_n1), .B(
        dp_if_stage_add_77_n18), .Z(dp_if_stage_NPC_4_i_31_) );
  XOR2_X1 dp_id_stage_U147 ( .A(dp_rd_fwd_wb_i[4]), .B(dp_id_stage_n27), .Z(
        dp_id_stage_p_addr_wRD[4]) );
  NOR2_X1 dp_id_stage_U146 ( .A1(dp_rd_fwd_wb_i[3]), .A2(dp_id_stage_n26), 
        .ZN(dp_id_stage_n27) );
  XNOR2_X1 dp_id_stage_U145 ( .A(dp_rd_fwd_wb_i[3]), .B(dp_id_stage_n26), .ZN(
        dp_id_stage_p_addr_wRD[3]) );
  OAI21_X1 dp_id_stage_U144 ( .B1(dp_id_stage_n25), .B2(dp_id_stage_n28), .A(
        dp_id_stage_n26), .ZN(dp_id_stage_p_addr_wRD[2]) );
  NAND2_X1 dp_id_stage_U143 ( .A1(dp_id_stage_n25), .A2(dp_id_stage_n28), .ZN(
        dp_id_stage_n26) );
  AOI21_X1 dp_id_stage_U142 ( .B1(dp_rd_fwd_wb_i[0]), .B2(dp_rd_fwd_wb_i[1]), 
        .A(dp_id_stage_n25), .ZN(dp_id_stage_n24) );
  NOR2_X1 dp_id_stage_U141 ( .A1(dp_rd_fwd_wb_i[1]), .A2(dp_rd_fwd_wb_i[0]), 
        .ZN(dp_id_stage_n25) );
  XOR2_X1 dp_id_stage_U140 ( .A(dp_ir_20_), .B(dp_id_stage_n15), .Z(
        dp_id_stage_p_addr_wRS2[4]) );
  NOR2_X1 dp_id_stage_U139 ( .A1(dp_ir_19_), .A2(dp_id_stage_n14), .ZN(
        dp_id_stage_n15) );
  XNOR2_X1 dp_id_stage_U138 ( .A(dp_ir_19_), .B(dp_id_stage_n14), .ZN(
        dp_id_stage_p_addr_wRS2[3]) );
  OAI21_X1 dp_id_stage_U137 ( .B1(dp_id_stage_n13), .B2(dp_id_stage_n16), .A(
        dp_id_stage_n14), .ZN(dp_id_stage_p_addr_wRS2[2]) );
  NAND2_X1 dp_id_stage_U136 ( .A1(dp_id_stage_n13), .A2(dp_id_stage_n16), .ZN(
        dp_id_stage_n14) );
  AOI21_X1 dp_id_stage_U135 ( .B1(dp_ir_16_), .B2(dp_ir_17_), .A(
        dp_id_stage_n13), .ZN(dp_id_stage_n12) );
  NOR2_X1 dp_id_stage_U134 ( .A1(dp_ir_17_), .A2(dp_ir_16_), .ZN(
        dp_id_stage_n13) );
  XOR2_X1 dp_id_stage_U133 ( .A(dp_ir_25_), .B(dp_id_stage_n10), .Z(
        dp_id_stage_p_addr_wRS1[4]) );
  NOR2_X1 dp_id_stage_U132 ( .A1(dp_ir_24_), .A2(dp_id_stage_n9), .ZN(
        dp_id_stage_n10) );
  XNOR2_X1 dp_id_stage_U131 ( .A(dp_ir_24_), .B(dp_id_stage_n9), .ZN(
        dp_id_stage_p_addr_wRS1[3]) );
  OAI21_X1 dp_id_stage_U130 ( .B1(dp_id_stage_n8), .B2(dp_id_stage_n11), .A(
        dp_id_stage_n9), .ZN(dp_id_stage_p_addr_wRS1[2]) );
  NAND2_X1 dp_id_stage_U129 ( .A1(dp_id_stage_n8), .A2(dp_id_stage_n11), .ZN(
        dp_id_stage_n9) );
  AOI21_X1 dp_id_stage_U128 ( .B1(dp_ir_21_), .B2(dp_ir_22_), .A(
        dp_id_stage_n8), .ZN(dp_id_stage_n7) );
  NOR2_X1 dp_id_stage_U127 ( .A1(dp_ir_22_), .A2(dp_ir_21_), .ZN(
        dp_id_stage_n8) );
  INV_X1 dp_id_stage_U126 ( .A(dp_ir_23_), .ZN(dp_id_stage_n11) );
  INV_X1 dp_id_stage_U125 ( .A(dp_ir_18_), .ZN(dp_id_stage_n16) );
  INV_X1 dp_id_stage_U124 ( .A(dp_id_stage_n7), .ZN(dp_id_stage_p_addr_wRS1[1]) );
  INV_X1 dp_id_stage_U123 ( .A(dp_ir_21_), .ZN(dp_id_stage_p_addr_wRS1[0]) );
  INV_X1 dp_id_stage_U122 ( .A(dp_id_stage_n12), .ZN(
        dp_id_stage_p_addr_wRS2[1]) );
  INV_X1 dp_id_stage_U121 ( .A(dp_ir_16_), .ZN(dp_id_stage_p_addr_wRS2[0]) );
  INV_X1 dp_id_stage_U120 ( .A(dp_rd_fwd_wb_i[2]), .ZN(dp_id_stage_n28) );
  INV_X1 dp_id_stage_U119 ( .A(dp_rd_fwd_wb_i[0]), .ZN(
        dp_id_stage_p_addr_wRD[0]) );
  OR3_X1 dp_id_stage_U118 ( .A1(dp_ir_20_), .A2(dp_ir_19_), .A3(dp_ir_18_), 
        .ZN(dp_id_stage_n18) );
  OR3_X1 dp_id_stage_U117 ( .A1(dp_ir_17_), .A2(dp_ir_16_), .A3(
        dp_id_stage_n18), .ZN(dp_id_stage_n17) );
  OR3_X1 dp_id_stage_U116 ( .A1(dp_ir_25_), .A2(dp_ir_24_), .A3(dp_ir_23_), 
        .ZN(dp_id_stage_n20) );
  OR3_X1 dp_id_stage_U115 ( .A1(dp_ir_22_), .A2(dp_ir_21_), .A3(
        dp_id_stage_n20), .ZN(dp_id_stage_n19) );
  INV_X1 dp_id_stage_U114 ( .A(dp_id_stage_n24), .ZN(dp_id_stage_p_addr_wRD[1]) );
  INV_X1 dp_id_stage_U113 ( .A(imm_uns_i), .ZN(dp_id_stage_n39) );
  INV_X1 dp_id_stage_U112 ( .A(dp_ir_22_), .ZN(dp_id_stage_n35) );
  OAI21_X1 dp_id_stage_U111 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n35), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[22]) );
  AND2_X1 dp_id_stage_U110 ( .A1(dp_id_stage_out2_i[3]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[3]) );
  AND2_X1 dp_id_stage_U109 ( .A1(dp_id_stage_out2_i[4]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[4]) );
  AND2_X1 dp_id_stage_U108 ( .A1(dp_id_stage_out2_i[5]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[5]) );
  AND2_X1 dp_id_stage_U107 ( .A1(dp_id_stage_out2_i[6]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[6]) );
  AND2_X1 dp_id_stage_U106 ( .A1(dp_id_stage_out2_i[7]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[7]) );
  AND2_X1 dp_id_stage_U105 ( .A1(dp_id_stage_out2_i[8]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[8]) );
  AND2_X1 dp_id_stage_U104 ( .A1(dp_id_stage_out2_i[9]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[9]) );
  AND2_X1 dp_id_stage_U103 ( .A1(dp_id_stage_out2_i[10]), .A2(dp_id_stage_n6), 
        .ZN(dp_rf_out2_id_o[10]) );
  AND2_X1 dp_id_stage_U102 ( .A1(dp_id_stage_out2_i[11]), .A2(dp_id_stage_n6), 
        .ZN(dp_rf_out2_id_o[11]) );
  AND2_X1 dp_id_stage_U101 ( .A1(dp_id_stage_out2_i[12]), .A2(dp_id_stage_n6), 
        .ZN(dp_rf_out2_id_o[12]) );
  AND2_X1 dp_id_stage_U100 ( .A1(dp_id_stage_out2_i[13]), .A2(dp_id_stage_n6), 
        .ZN(dp_rf_out2_id_o[13]) );
  AND2_X1 dp_id_stage_U99 ( .A1(dp_id_stage_out2_i[14]), .A2(dp_id_stage_n6), 
        .ZN(dp_rf_out2_id_o[14]) );
  AND2_X1 dp_id_stage_U98 ( .A1(dp_id_stage_out2_i[15]), .A2(dp_id_stage_n6), 
        .ZN(dp_rf_out2_id_o[15]) );
  AND2_X1 dp_id_stage_U97 ( .A1(dp_id_stage_out2_i[16]), .A2(dp_id_stage_n6), 
        .ZN(dp_rf_out2_id_o[16]) );
  AND2_X1 dp_id_stage_U96 ( .A1(dp_id_stage_out2_i[17]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[17]) );
  AND2_X1 dp_id_stage_U95 ( .A1(dp_id_stage_out2_i[18]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[18]) );
  AND2_X1 dp_id_stage_U94 ( .A1(dp_id_stage_out2_i[19]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[19]) );
  AND2_X1 dp_id_stage_U93 ( .A1(dp_id_stage_out2_i[20]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[20]) );
  AND2_X1 dp_id_stage_U92 ( .A1(dp_id_stage_out2_i[21]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[21]) );
  AND2_X1 dp_id_stage_U91 ( .A1(dp_id_stage_out1_i[0]), .A2(dp_id_stage_n3), 
        .ZN(dp_rf_out1_id_o[0]) );
  AND2_X1 dp_id_stage_U90 ( .A1(dp_id_stage_out2_i[22]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[22]) );
  AND2_X1 dp_id_stage_U89 ( .A1(dp_id_stage_out2_i[23]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[23]) );
  AND2_X1 dp_id_stage_U88 ( .A1(dp_id_stage_out2_i[24]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[24]) );
  AND2_X1 dp_id_stage_U87 ( .A1(dp_id_stage_out2_i[25]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[25]) );
  AND2_X1 dp_id_stage_U86 ( .A1(dp_id_stage_out2_i[26]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[26]) );
  AND2_X1 dp_id_stage_U85 ( .A1(dp_id_stage_out2_i[27]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[27]) );
  AND2_X1 dp_id_stage_U84 ( .A1(dp_id_stage_out2_i[28]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[28]) );
  AND2_X1 dp_id_stage_U83 ( .A1(dp_id_stage_out2_i[29]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[29]) );
  AND2_X1 dp_id_stage_U82 ( .A1(dp_id_stage_out2_i[30]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[30]) );
  AND2_X1 dp_id_stage_U81 ( .A1(dp_id_stage_out2_i[31]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[31]) );
  AND2_X1 dp_id_stage_U80 ( .A1(dp_id_stage_out1_i[1]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[1]) );
  AND2_X1 dp_id_stage_U79 ( .A1(dp_id_stage_out1_i[2]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[2]) );
  AND2_X1 dp_id_stage_U78 ( .A1(dp_id_stage_out1_i[3]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[3]) );
  AND2_X1 dp_id_stage_U77 ( .A1(dp_id_stage_out1_i[4]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[4]) );
  AND2_X1 dp_id_stage_U76 ( .A1(dp_id_stage_out1_i[5]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[5]) );
  AND2_X1 dp_id_stage_U75 ( .A1(dp_id_stage_out1_i[6]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[6]) );
  AND2_X1 dp_id_stage_U74 ( .A1(dp_id_stage_out1_i[7]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[7]) );
  AND2_X1 dp_id_stage_U73 ( .A1(dp_id_stage_out1_i[8]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[8]) );
  AND2_X1 dp_id_stage_U72 ( .A1(dp_id_stage_out1_i[9]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[9]) );
  AND2_X1 dp_id_stage_U71 ( .A1(dp_id_stage_out1_i[10]), .A2(dp_id_stage_n3), 
        .ZN(dp_rf_out1_id_o[10]) );
  AND2_X1 dp_id_stage_U70 ( .A1(dp_id_stage_out1_i[11]), .A2(dp_id_stage_n3), 
        .ZN(dp_rf_out1_id_o[11]) );
  AND2_X1 dp_id_stage_U69 ( .A1(dp_id_stage_out1_i[12]), .A2(dp_id_stage_n3), 
        .ZN(dp_rf_out1_id_o[12]) );
  AND2_X1 dp_id_stage_U68 ( .A1(dp_id_stage_out1_i[13]), .A2(dp_id_stage_n3), 
        .ZN(dp_rf_out1_id_o[13]) );
  AND2_X1 dp_id_stage_U67 ( .A1(dp_id_stage_out1_i[14]), .A2(dp_id_stage_n3), 
        .ZN(dp_rf_out1_id_o[14]) );
  AND2_X1 dp_id_stage_U66 ( .A1(dp_id_stage_out1_i[15]), .A2(dp_id_stage_n3), 
        .ZN(dp_rf_out1_id_o[15]) );
  AND2_X1 dp_id_stage_U65 ( .A1(dp_id_stage_out1_i[16]), .A2(dp_id_stage_n3), 
        .ZN(dp_rf_out1_id_o[16]) );
  AND2_X1 dp_id_stage_U64 ( .A1(dp_id_stage_out1_i[17]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[17]) );
  AND2_X1 dp_id_stage_U63 ( .A1(dp_id_stage_out1_i[18]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[18]) );
  AND2_X1 dp_id_stage_U62 ( .A1(dp_id_stage_out1_i[19]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[19]) );
  AND2_X1 dp_id_stage_U61 ( .A1(dp_id_stage_out1_i[20]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[20]) );
  AND2_X1 dp_id_stage_U60 ( .A1(dp_id_stage_out1_i[21]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[21]) );
  AND2_X1 dp_id_stage_U59 ( .A1(dp_id_stage_out1_i[22]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[22]) );
  AND2_X1 dp_id_stage_U58 ( .A1(dp_id_stage_out1_i[23]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[23]) );
  AND2_X1 dp_id_stage_U57 ( .A1(dp_id_stage_out1_i[24]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[24]) );
  INV_X1 dp_id_stage_U56 ( .A(dp_ir_16_), .ZN(dp_id_stage_n29) );
  OAI21_X1 dp_id_stage_U55 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n29), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[16]) );
  INV_X1 dp_id_stage_U54 ( .A(dp_ir_19_), .ZN(dp_id_stage_n32) );
  OAI21_X1 dp_id_stage_U53 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n32), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[19]) );
  INV_X1 dp_id_stage_U52 ( .A(dp_ir_20_), .ZN(dp_id_stage_n33) );
  OAI21_X1 dp_id_stage_U51 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n33), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[20]) );
  INV_X1 dp_id_stage_U50 ( .A(dp_ir_23_), .ZN(dp_id_stage_n36) );
  OAI21_X1 dp_id_stage_U49 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n36), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[23]) );
  INV_X1 dp_id_stage_U48 ( .A(dp_ir_18_), .ZN(dp_id_stage_n31) );
  OAI21_X1 dp_id_stage_U47 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n31), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[18]) );
  INV_X1 dp_id_stage_U46 ( .A(dp_ir_21_), .ZN(dp_id_stage_n34) );
  OAI21_X1 dp_id_stage_U45 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n34), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[21]) );
  INV_X1 dp_id_stage_U44 ( .A(dp_ir_24_), .ZN(dp_id_stage_n37) );
  OAI21_X1 dp_id_stage_U43 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n37), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[24]) );
  INV_X1 dp_id_stage_U42 ( .A(dp_ir_17_), .ZN(dp_id_stage_n30) );
  OAI21_X1 dp_id_stage_U41 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n30), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[17]) );
  AND2_X1 dp_id_stage_U40 ( .A1(dp_id_stage_out1_i[31]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[31]) );
  AND2_X1 dp_id_stage_U39 ( .A1(dp_id_stage_out1_i[26]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[26]) );
  AND2_X1 dp_id_stage_U38 ( .A1(dp_id_stage_out1_i[29]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[29]) );
  AND2_X1 dp_id_stage_U37 ( .A1(dp_id_stage_out1_i[25]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[25]) );
  AND2_X1 dp_id_stage_U36 ( .A1(dp_id_stage_out1_i[27]), .A2(dp_id_stage_n2), 
        .ZN(dp_rf_out1_id_o[27]) );
  AND2_X1 dp_id_stage_U35 ( .A1(dp_id_stage_out1_i[28]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[28]) );
  AND2_X1 dp_id_stage_U34 ( .A1(dp_id_stage_out1_i[30]), .A2(dp_id_stage_n1), 
        .ZN(dp_rf_out1_id_o[30]) );
  AND2_X1 dp_id_stage_U33 ( .A1(dp_id_stage_out2_i[0]), .A2(dp_id_stage_n6), 
        .ZN(dp_rf_out2_id_o[0]) );
  AND2_X1 dp_id_stage_U32 ( .A1(dp_id_stage_out2_i[1]), .A2(dp_id_stage_n5), 
        .ZN(dp_rf_out2_id_o[1]) );
  AND2_X1 dp_id_stage_U31 ( .A1(dp_id_stage_out2_i[2]), .A2(dp_id_stage_n4), 
        .ZN(dp_rf_out2_id_o[2]) );
  AND2_X1 dp_id_stage_U30 ( .A1(dp_ir_14_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[14]) );
  AND2_X1 dp_id_stage_U29 ( .A1(dp_ir_1_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[1]) );
  AND2_X1 dp_id_stage_U28 ( .A1(dp_ir_2_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[2]) );
  AND2_X1 dp_id_stage_U27 ( .A1(dp_ir_4_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[4]) );
  AND2_X1 dp_id_stage_U26 ( .A1(dp_ir_5_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[5]) );
  AND2_X1 dp_id_stage_U25 ( .A1(dp_ir_7_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[7]) );
  AND2_X1 dp_id_stage_U24 ( .A1(dp_ir_11_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[11]) );
  AND2_X1 dp_id_stage_U23 ( .A1(dp_ir_0_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[0]) );
  AND2_X1 dp_id_stage_U22 ( .A1(dp_ir_3_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[3]) );
  AND2_X1 dp_id_stage_U21 ( .A1(dp_ir_6_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[6]) );
  AND2_X1 dp_id_stage_U20 ( .A1(dp_ir_8_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[8]) );
  AND2_X1 dp_id_stage_U19 ( .A1(dp_ir_9_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[9]) );
  AND2_X1 dp_id_stage_U18 ( .A1(dp_ir_10_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[10]) );
  AND2_X1 dp_id_stage_U17 ( .A1(dp_ir_12_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[12]) );
  AND2_X1 dp_id_stage_U16 ( .A1(dp_ir_13_), .A2(dp_id_stage_n21), .ZN(
        dp_imm_id_o[13]) );
  AND2_X1 dp_id_stage_U15 ( .A1(dp_id_stage_n21), .A2(dp_ir_15_), .ZN(
        dp_imm_id_o[15]) );
  NAND2_X1 dp_id_stage_U14 ( .A1(imm_isoff_i), .A2(dp_id_stage_n22), .ZN(
        dp_id_stage_n21) );
  NAND2_X1 dp_id_stage_U13 ( .A1(imm_isoff_i), .A2(dp_id_stage_n39), .ZN(
        dp_id_stage_n22) );
  INV_X1 dp_id_stage_U12 ( .A(imm_isoff_i), .ZN(dp_id_stage_n40) );
  NAND3_X1 dp_id_stage_U11 ( .A1(dp_id_stage_n40), .A2(dp_id_stage_n39), .A3(
        dp_ir_15_), .ZN(dp_id_stage_n23) );
  INV_X1 dp_id_stage_U10 ( .A(dp_ir_25_), .ZN(dp_id_stage_n38) );
  OAI21_X1 dp_id_stage_U9 ( .B1(dp_id_stage_n22), .B2(dp_id_stage_n38), .A(
        dp_id_stage_n23), .ZN(dp_imm_id_o[31]) );
  BUF_X1 dp_id_stage_U8 ( .A(dp_id_stage_n17), .Z(dp_id_stage_n6) );
  BUF_X1 dp_id_stage_U7 ( .A(dp_id_stage_n19), .Z(dp_id_stage_n3) );
  BUF_X1 dp_id_stage_U6 ( .A(dp_id_stage_n17), .Z(dp_id_stage_n5) );
  BUF_X1 dp_id_stage_U5 ( .A(dp_id_stage_n17), .Z(dp_id_stage_n4) );
  BUF_X1 dp_id_stage_U4 ( .A(dp_id_stage_n19), .Z(dp_id_stage_n2) );
  BUF_X1 dp_id_stage_U3 ( .A(dp_id_stage_n19), .Z(dp_id_stage_n1) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U46 ( .A(1'b0), .ZN(
        dp_id_stage_regfile_ControlUnit_n41) );
  AND2_X1 dp_id_stage_regfile_ControlUnit_U45 ( .A1(
        dp_id_stage_regfile_canrestore), .A2(1'b0), .ZN(
        dp_id_stage_regfile_ControlUnit_n24) );
  OAI22_X1 dp_id_stage_regfile_ControlUnit_U44 ( .A1(
        dp_id_stage_regfile_cansave), .A2(dp_id_stage_regfile_ControlUnit_n41), 
        .B1(1'b0), .B2(dp_id_stage_regfile_ControlUnit_n24), .ZN(
        dp_id_stage_regfile_ControlUnit_n23) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U43 ( .A(dp_id_stage_regfile_end_sf), 
        .ZN(dp_id_stage_regfile_ControlUnit_n16) );
  AND3_X1 dp_id_stage_regfile_ControlUnit_U42 ( .A1(
        dp_id_stage_regfile_ControlUnit_n13), .A2(
        dp_id_stage_regfile_ControlUnit_n12), .A3(
        dp_id_stage_regfile_ControlUnit_current_state_3_), .ZN(
        dp_id_stage_regfile_cnt_swp) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U41 ( .A1(1'b0), .A2(
        dp_id_stage_regfile_ControlUnit_n6), .ZN(
        dp_id_stage_regfile_ControlUnit_n19) );
  AOI21_X1 dp_id_stage_regfile_ControlUnit_U40 ( .B1(
        dp_id_stage_regfile_ControlUnit_n17), .B2(
        dp_id_stage_regfile_ControlUnit_n19), .A(RST), .ZN(
        dp_id_stage_regfile_ControlUnit_next_state[1]) );
  AOI21_X1 dp_id_stage_regfile_ControlUnit_U39 ( .B1(
        dp_id_stage_regfile_ControlUnit_n17), .B2(
        dp_id_stage_regfile_ControlUnit_n18), .A(RST), .ZN(
        dp_id_stage_regfile_ControlUnit_next_state[2]) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U38 ( .A(
        dp_id_stage_regfile_ControlUnit_n26), .ZN(
        dp_id_stage_regfile_ControlUnit_n15) );
  AOI21_X1 dp_id_stage_regfile_ControlUnit_U37 ( .B1(
        dp_id_stage_regfile_ControlUnit_n6), .B2(
        dp_id_stage_regfile_ControlUnit_n23), .A(dp_id_stage_regfile_rd_cu), 
        .ZN(dp_id_stage_regfile_ControlUnit_n22) );
  AOI22_X1 dp_id_stage_regfile_ControlUnit_U36 ( .A1(
        dp_id_stage_regfile_ControlUnit_n15), .A2(
        dp_id_stage_regfile_ControlUnit_n12), .B1(
        dp_id_stage_regfile_ControlUnit_n25), .B2(
        dp_id_stage_regfile_ControlUnit_n14), .ZN(
        dp_id_stage_regfile_ControlUnit_n21) );
  AOI21_X1 dp_id_stage_regfile_ControlUnit_U35 ( .B1(
        dp_id_stage_regfile_ControlUnit_n21), .B2(
        dp_id_stage_regfile_ControlUnit_n22), .A(RST), .ZN(
        dp_id_stage_regfile_ControlUnit_next_state[0]) );
  NOR3_X1 dp_id_stage_regfile_ControlUnit_U34 ( .A1(
        dp_id_stage_regfile_ControlUnit_n16), .A2(RST), .A3(
        dp_id_stage_regfile_ControlUnit_n9), .ZN(
        dp_id_stage_regfile_ControlUnit_next_state[3]) );
  AOI21_X1 dp_id_stage_regfile_ControlUnit_U33 ( .B1(
        dp_id_stage_regfile_ControlUnit_n13), .B2(
        dp_id_stage_regfile_ControlUnit_current_state_3_), .A(
        dp_id_stage_regfile_ControlUnit_n27), .ZN(
        dp_id_stage_regfile_ControlUnit_n26) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U32 ( .A(
        dp_id_stage_regfile_ControlUnit_n29), .ZN(dp_id_stage_regfile_wr_cu)
         );
  NOR2_X1 dp_id_stage_regfile_ControlUnit_U31 ( .A1(
        dp_id_stage_regfile_ControlUnit_n14), .A2(
        dp_id_stage_regfile_ControlUnit_current_state_2_), .ZN(
        dp_id_stage_regfile_ControlUnit_n40) );
  AND2_X2 dp_id_stage_regfile_ControlUnit_U30 ( .A1(
        dp_id_stage_regfile_ControlUnit_n1), .A2(
        dp_id_stage_regfile_ControlUnit_n13), .ZN(
        dp_id_stage_regfile_ControlUnit_n25) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U29 ( .A(
        dp_id_stage_regfile_up_dwn_cwp), .ZN(
        dp_id_stage_regfile_ControlUnit_n5) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U28 ( .A1(
        dp_id_stage_regfile_ControlUnit_n35), .A2(
        dp_id_stage_regfile_ControlUnit_n5), .ZN(
        dp_id_stage_regfile_up_dwn_rest) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U27 ( .A1(
        dp_id_stage_regfile_ControlUnit_n35), .A2(
        dp_id_stage_regfile_ControlUnit_n29), .ZN(rf_fill_i) );
  AND3_X1 dp_id_stage_regfile_ControlUnit_U26 ( .A1(
        dp_id_stage_regfile_ControlUnit_n38), .A2(
        dp_id_stage_regfile_ControlUnit_n32), .A3(
        dp_id_stage_regfile_ControlUnit_n39), .ZN(
        dp_id_stage_regfile_ControlUnit_n34) );
  NAND4_X1 dp_id_stage_regfile_ControlUnit_U25 ( .A1(
        dp_id_stage_regfile_ControlUnit_n30), .A2(
        dp_id_stage_regfile_ControlUnit_n31), .A3(
        dp_id_stage_regfile_ControlUnit_n32), .A4(
        dp_id_stage_regfile_ControlUnit_n9), .ZN(
        dp_id_stage_regfile_up_dwn_swp) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U24 ( .A1(
        dp_id_stage_regfile_ControlUnit_n37), .A2(
        dp_id_stage_regfile_ControlUnit_n28), .ZN(rf_spill_i) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U23 ( .A(rf_spill_i), .ZN(
        dp_id_stage_regfile_ControlUnit_n4) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U22 ( .A1(
        dp_id_stage_regfile_ControlUnit_n30), .A2(
        dp_id_stage_regfile_ControlUnit_n4), .ZN(dp_id_stage_regfile_sel_wp)
         );
  INV_X1 dp_id_stage_regfile_ControlUnit_U21 ( .A(
        dp_id_stage_regfile_ControlUnit_n28), .ZN(dp_id_stage_regfile_rd_cu)
         );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U20 ( .A1(
        dp_id_stage_regfile_ControlUnit_n40), .A2(
        dp_id_stage_regfile_ControlUnit_n25), .ZN(
        dp_id_stage_regfile_ControlUnit_n38) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U19 ( .A1(
        dp_id_stage_regfile_ControlUnit_n36), .A2(
        dp_id_stage_regfile_ControlUnit_n33), .ZN(dp_id_stage_regfile_cnt_save) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U18 ( .A1(
        dp_id_stage_regfile_ControlUnit_n37), .A2(
        dp_id_stage_regfile_ControlUnit_n35), .ZN(
        dp_id_stage_regfile_ControlUnit_n20) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U17 ( .A(
        dp_id_stage_regfile_ControlUnit_n32), .ZN(dp_id_stage_regfile_rst_rf)
         );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U16 ( .A1(
        dp_id_stage_regfile_ControlUnit_n40), .A2(
        dp_id_stage_regfile_ControlUnit_n27), .ZN(
        dp_id_stage_regfile_ControlUnit_n37) );
  NOR2_X1 dp_id_stage_regfile_ControlUnit_U15 ( .A1(
        dp_id_stage_regfile_cnt_swp), .A2(dp_id_stage_regfile_rf_enable), .ZN(
        dp_id_stage_regfile_ControlUnit_n39) );
  AOI21_X1 dp_id_stage_regfile_ControlUnit_U14 ( .B1(
        dp_id_stage_regfile_ControlUnit_n16), .B2(
        dp_id_stage_regfile_rf_enable), .A(dp_id_stage_regfile_ControlUnit_n20), .ZN(dp_id_stage_regfile_ControlUnit_n17) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U13 ( .A1(
        dp_id_stage_regfile_ControlUnit_n29), .A2(
        dp_id_stage_regfile_ControlUnit_n28), .ZN(
        dp_id_stage_regfile_rf_enable) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U12 ( .A(
        dp_id_stage_regfile_ControlUnit_n20), .ZN(
        dp_id_stage_regfile_ControlUnit_n3) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U11 ( .A(dp_id_stage_regfile_cnt_save), .ZN(dp_id_stage_regfile_ControlUnit_n10) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U10 ( .A(
        dp_id_stage_regfile_rf_enable), .ZN(dp_id_stage_regfile_ControlUnit_n9) );
  INV_X1 dp_id_stage_regfile_ControlUnit_U9 ( .A(
        dp_id_stage_regfile_ControlUnit_n38), .ZN(
        dp_id_stage_regfile_ControlUnit_n6) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U8 ( .A1(
        dp_id_stage_regfile_ControlUnit_n39), .A2(
        dp_id_stage_regfile_ControlUnit_n31), .ZN(dp_id_stage_regfile_rst_swp)
         );
  NAND4_X1 dp_id_stage_regfile_ControlUnit_U7 ( .A1(
        dp_id_stage_regfile_ControlUnit_n39), .A2(
        dp_id_stage_regfile_ControlUnit_n37), .A3(
        dp_id_stage_regfile_ControlUnit_n38), .A4(
        dp_id_stage_regfile_ControlUnit_n10), .ZN(
        dp_id_stage_regfile_rst_spill_fill) );
  NAND2_X1 dp_id_stage_regfile_ControlUnit_U6 ( .A1(
        dp_id_stage_regfile_ControlUnit_n3), .A2(
        dp_id_stage_regfile_ControlUnit_n10), .ZN(dp_id_stage_regfile_cnt_cwp)
         );
  NOR2_X1 dp_id_stage_regfile_ControlUnit_U5 ( .A1(
        dp_id_stage_regfile_ControlUnit_n6), .A2(dp_id_stage_regfile_cnt_cwp), 
        .ZN(dp_id_stage_regfile_ControlUnit_n31) );
  INV_X2 dp_id_stage_regfile_ControlUnit_U4 ( .A(
        dp_id_stage_regfile_ControlUnit_n31), .ZN(dp_id_stage_regfile_cpu_work) );
  NOR2_X1 dp_id_stage_regfile_ControlUnit_U3 ( .A1(
        dp_id_stage_regfile_ControlUnit_n13), .A2(
        dp_id_stage_regfile_ControlUnit_current_state_3_), .ZN(
        dp_id_stage_regfile_ControlUnit_n27) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U56 ( .A1(
        dp_id_stage_regfile_ControlUnit_current_state_2_), .A2(
        dp_id_stage_regfile_ControlUnit_current_state_0_), .A3(
        dp_id_stage_regfile_ControlUnit_n25), .ZN(
        dp_id_stage_regfile_ControlUnit_n35) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U55 ( .A1(
        dp_id_stage_regfile_ControlUnit_n14), .A2(
        dp_id_stage_regfile_ControlUnit_n12), .A3(
        dp_id_stage_regfile_ControlUnit_n27), .ZN(
        dp_id_stage_regfile_ControlUnit_n36) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U54 ( .A1(
        dp_id_stage_regfile_ControlUnit_current_state_2_), .A2(
        dp_id_stage_regfile_ControlUnit_n14), .A3(
        dp_id_stage_regfile_ControlUnit_n25), .ZN(
        dp_id_stage_regfile_ControlUnit_n33) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U53 ( .A1(
        dp_id_stage_regfile_ControlUnit_n27), .A2(
        dp_id_stage_regfile_ControlUnit_n14), .A3(
        dp_id_stage_regfile_ControlUnit_current_state_2_), .ZN(
        dp_id_stage_regfile_ControlUnit_n29) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U52 ( .A1(
        dp_id_stage_regfile_ControlUnit_n14), .A2(
        dp_id_stage_regfile_ControlUnit_n12), .A3(
        dp_id_stage_regfile_ControlUnit_n25), .ZN(
        dp_id_stage_regfile_ControlUnit_n32) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U51 ( .A1(
        dp_id_stage_regfile_ControlUnit_current_state_0_), .A2(
        dp_id_stage_regfile_ControlUnit_n27), .A3(
        dp_id_stage_regfile_ControlUnit_current_state_2_), .ZN(
        dp_id_stage_regfile_ControlUnit_n28) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U50 ( .A1(
        dp_id_stage_regfile_ControlUnit_n40), .A2(
        dp_id_stage_regfile_ControlUnit_n13), .A3(
        dp_id_stage_regfile_ControlUnit_current_state_3_), .ZN(
        dp_id_stage_regfile_ControlUnit_n30) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U49 ( .A1(
        dp_id_stage_regfile_ControlUnit_n36), .A2(
        dp_id_stage_regfile_ControlUnit_n37), .A3(
        dp_id_stage_regfile_ControlUnit_n34), .ZN(
        dp_id_stage_regfile_up_dwn_cwp) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U48 ( .A1(
        dp_id_stage_regfile_ControlUnit_n3), .A2(
        dp_id_stage_regfile_ControlUnit_n33), .A3(
        dp_id_stage_regfile_ControlUnit_n34), .ZN(
        dp_id_stage_regfile_up_dwn_save) );
  NAND3_X1 dp_id_stage_regfile_ControlUnit_U47 ( .A1(
        dp_id_stage_regfile_ControlUnit_n6), .A2(
        dp_id_stage_regfile_ControlUnit_n41), .A3(1'b0), .ZN(
        dp_id_stage_regfile_ControlUnit_n18) );
  DFF_X1 dp_id_stage_regfile_ControlUnit_current_state_reg_3_ ( .D(
        dp_id_stage_regfile_ControlUnit_next_state[3]), .CK(CLK), .Q(
        dp_id_stage_regfile_ControlUnit_current_state_3_), .QN(
        dp_id_stage_regfile_ControlUnit_n1) );
  DFF_X1 dp_id_stage_regfile_ControlUnit_current_state_reg_2_ ( .D(
        dp_id_stage_regfile_ControlUnit_next_state[2]), .CK(CLK), .Q(
        dp_id_stage_regfile_ControlUnit_current_state_2_), .QN(
        dp_id_stage_regfile_ControlUnit_n12) );
  DFF_X1 dp_id_stage_regfile_ControlUnit_current_state_reg_1_ ( .D(
        dp_id_stage_regfile_ControlUnit_next_state[1]), .CK(CLK), .QN(
        dp_id_stage_regfile_ControlUnit_n13) );
  DFF_X1 dp_id_stage_regfile_ControlUnit_current_state_reg_0_ ( .D(
        dp_id_stage_regfile_ControlUnit_next_state[0]), .CK(CLK), .Q(
        dp_id_stage_regfile_ControlUnit_current_state_0_), .QN(
        dp_id_stage_regfile_ControlUnit_n14) );
  AND3_X1 dp_id_stage_regfile_DataPath_U4 ( .A1(
        dp_id_stage_regfile_DataPath_addr_sf_in_1_), .A2(
        dp_id_stage_regfile_DataPath_addr_sf_in_0_), .A3(
        dp_id_stage_regfile_DataPath_addr_sf_in_2_), .ZN(
        dp_id_stage_regfile_end_sf) );
  INV_X1 dp_id_stage_regfile_DataPath_U3 ( .A(
        dp_id_stage_regfile_DataPath_CWP_0_), .ZN(
        dp_id_stage_regfile_DataPath_cwp_1_0_) );
  AOI21_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U20 ( .B1(
        dp_id_stage_p_addr_wRS1[3]), .B2(dp_id_stage_p_addr_wRS1[2]), .A(
        dp_id_stage_p_addr_wRS1[4]), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_N1) );
  XNOR2_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U19 ( .A(
        dp_id_stage_p_addr_wRS1[3]), .B(dp_id_stage_regfile_DataPath_CWP_0_), 
        .ZN(dp_id_stage_regfile_DataPath_Conv_RD1_n18) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U18 ( .A(
        dp_id_stage_p_addr_wRS1[3]), .B(dp_id_stage_p_addr_wRS1[2]), .Z(
        dp_id_stage_regfile_DataPath_Conv_RD1_n4) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U17 ( .A1(
        dp_id_stage_p_addr_wRS1[3]), .A2(dp_id_stage_p_addr_wRS1[2]), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_n3) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U16 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_RD1_N5), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD1_n8), .B1(
        dp_id_stage_p_addr_wRS1[2]), .B2(
        dp_id_stage_regfile_DataPath_Conv_RD1_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_n20) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U15 ( .A(
        dp_id_stage_regfile_DataPath_Conv_RD1_n20), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd1_p[2]) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U14 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_RD1_n1), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD1_n8), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd1_p[4]) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U13 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_RD1_n2), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD1_n8), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd1_p[5]) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U12 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_RD1_n4), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD1_n8), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_n19) );
  OAI21_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U11 ( .B1(
        dp_id_stage_regfile_DataPath_Conv_RD1_n18), .B2(
        dp_id_stage_regfile_DataPath_Conv_RD1_n8), .A(
        dp_id_stage_regfile_DataPath_Conv_RD1_n19), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd1_p[3]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U10 ( .A1(
        dp_id_stage_p_addr_wRS1[1]), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD1_n8), .B1(
        dp_id_stage_p_addr_wRS1[1]), .B2(
        dp_id_stage_regfile_DataPath_Conv_RD1_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_n21) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U9 ( .A(
        dp_id_stage_regfile_DataPath_Conv_RD1_n21), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd1_p[1]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U8 ( .A1(
        dp_id_stage_p_addr_wRS1[0]), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD1_n8), .B1(
        dp_id_stage_p_addr_wRS1[0]), .B2(
        dp_id_stage_regfile_DataPath_Conv_RD1_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_n22) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U7 ( .A(
        dp_id_stage_regfile_DataPath_Conv_RD1_n22), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd1_p[0]) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U6 ( .A(
        dp_id_stage_p_addr_wRS1[2]), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_N5) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U5 ( .A(
        dp_id_stage_regfile_DataPath_Conv_RD1_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_n8) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U4 ( .A1(
        dp_id_stage_p_addr_wRS1[4]), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD1_n3), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD1_n2) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Conv_RD1_U3 ( .A(
        dp_id_stage_p_addr_wRS1[4]), .B(
        dp_id_stage_regfile_DataPath_Conv_RD1_n3), .Z(
        dp_id_stage_regfile_DataPath_Conv_RD1_n1) );
  AOI21_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U20 ( .B1(
        dp_id_stage_p_addr_wRS2[3]), .B2(dp_id_stage_p_addr_wRS2[2]), .A(
        dp_id_stage_p_addr_wRS2[4]), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_N1) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U19 ( .A1(
        dp_id_stage_p_addr_wRS2[1]), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD2_n8), .B1(
        dp_id_stage_p_addr_wRS2[1]), .B2(
        dp_id_stage_regfile_DataPath_Conv_RD2_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_n10) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U18 ( .A(
        dp_id_stage_regfile_DataPath_Conv_RD2_n10), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd2_p[1]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U17 ( .A1(
        dp_id_stage_p_addr_wRS2[0]), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD2_n8), .B1(
        dp_id_stage_p_addr_wRS2[0]), .B2(
        dp_id_stage_regfile_DataPath_Conv_RD2_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_n9) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U16 ( .A(
        dp_id_stage_regfile_DataPath_Conv_RD2_n9), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd2_p[0]) );
  XNOR2_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U15 ( .A(
        dp_id_stage_p_addr_wRS2[3]), .B(dp_id_stage_regfile_DataPath_CWP_0_), 
        .ZN(dp_id_stage_regfile_DataPath_Conv_RD2_n13) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U14 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_RD2_n1), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD2_n8), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_n12) );
  OAI21_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U13 ( .B1(
        dp_id_stage_regfile_DataPath_Conv_RD2_n13), .B2(
        dp_id_stage_regfile_DataPath_Conv_RD2_n8), .A(
        dp_id_stage_regfile_DataPath_Conv_RD2_n12), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd2_p[3]) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U12 ( .A1(
        dp_id_stage_p_addr_wRS2[3]), .A2(dp_id_stage_p_addr_wRS2[2]), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_n4) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U11 ( .A1(
        dp_id_stage_p_addr_wRS2[4]), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD2_n4), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_n3) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U10 ( .A(
        dp_id_stage_p_addr_wRS2[4]), .B(
        dp_id_stage_regfile_DataPath_Conv_RD2_n4), .Z(
        dp_id_stage_regfile_DataPath_Conv_RD2_n2) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U9 ( .A(
        dp_id_stage_p_addr_wRS2[2]), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_N5) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U8 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_RD2_N5), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD2_n8), .B1(
        dp_id_stage_p_addr_wRS2[2]), .B2(
        dp_id_stage_regfile_DataPath_Conv_RD2_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_n11) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U7 ( .A(
        dp_id_stage_regfile_DataPath_Conv_RD2_n11), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd2_p[2]) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U6 ( .A(
        dp_id_stage_regfile_DataPath_Conv_RD2_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_RD2_n8) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U5 ( .A(
        dp_id_stage_p_addr_wRS2[3]), .B(dp_id_stage_p_addr_wRS2[2]), .Z(
        dp_id_stage_regfile_DataPath_Conv_RD2_n1) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U4 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_RD2_n3), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD2_n8), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd2_p[5]) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_RD2_U3 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_RD2_n2), .A2(
        dp_id_stage_regfile_DataPath_Conv_RD2_n8), .ZN(
        dp_id_stage_regfile_DataPath_addr_rd2_p[4]) );
  AOI21_X1 dp_id_stage_regfile_DataPath_Conv_W_U20 ( .B1(
        dp_id_stage_p_addr_wRD[3]), .B2(dp_id_stage_p_addr_wRD[2]), .A(
        dp_id_stage_p_addr_wRD[4]), .ZN(dp_id_stage_regfile_DataPath_Conv_W_N1) );
  XNOR2_X1 dp_id_stage_regfile_DataPath_Conv_W_U19 ( .A(
        dp_id_stage_p_addr_wRD[3]), .B(dp_id_stage_regfile_DataPath_CWP_0_), 
        .ZN(dp_id_stage_regfile_DataPath_Conv_W_n13) );
  OAI21_X1 dp_id_stage_regfile_DataPath_Conv_W_U18 ( .B1(
        dp_id_stage_regfile_DataPath_Conv_W_n13), .B2(
        dp_id_stage_regfile_DataPath_Conv_W_n8), .A(
        dp_id_stage_regfile_DataPath_Conv_W_n12), .ZN(
        dp_id_stage_regfile_DataPath_addr_w_p[3]) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Conv_W_U17 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_W_n3), .A2(
        dp_id_stage_regfile_DataPath_Conv_W_n8), .ZN(
        dp_id_stage_regfile_DataPath_Conv_W_n12) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_W_U16 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_W_n2), .A2(
        dp_id_stage_regfile_DataPath_Conv_W_n8), .ZN(
        dp_id_stage_regfile_DataPath_addr_w_p[5]) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_W_U15 ( .A1(
        dp_id_stage_p_addr_wRD[3]), .A2(dp_id_stage_p_addr_wRD[2]), .ZN(
        dp_id_stage_regfile_DataPath_Conv_W_n4) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_W_U14 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_W_n1), .A2(
        dp_id_stage_regfile_DataPath_Conv_W_n8), .ZN(
        dp_id_stage_regfile_DataPath_addr_w_p[4]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_W_U13 ( .A1(
        dp_id_stage_p_addr_wRD[1]), .A2(dp_id_stage_regfile_DataPath_Conv_W_n8), .B1(dp_id_stage_p_addr_wRD[1]), .B2(dp_id_stage_regfile_DataPath_Conv_W_N1), 
        .ZN(dp_id_stage_regfile_DataPath_Conv_W_n10) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_W_U12 ( .A(
        dp_id_stage_regfile_DataPath_Conv_W_n10), .ZN(
        dp_id_stage_regfile_DataPath_addr_w_p[1]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_W_U11 ( .A1(
        dp_id_stage_p_addr_wRD[0]), .A2(dp_id_stage_regfile_DataPath_Conv_W_n8), .B1(dp_id_stage_p_addr_wRD[0]), .B2(dp_id_stage_regfile_DataPath_Conv_W_N1), 
        .ZN(dp_id_stage_regfile_DataPath_Conv_W_n9) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_W_U10 ( .A(
        dp_id_stage_regfile_DataPath_Conv_W_n9), .ZN(
        dp_id_stage_regfile_DataPath_addr_w_p[0]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Conv_W_U9 ( .A1(
        dp_id_stage_regfile_DataPath_Conv_W_N5), .A2(
        dp_id_stage_regfile_DataPath_Conv_W_n8), .B1(dp_id_stage_p_addr_wRD[2]), .B2(dp_id_stage_regfile_DataPath_Conv_W_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_W_n11) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_W_U8 ( .A(
        dp_id_stage_regfile_DataPath_Conv_W_n11), .ZN(
        dp_id_stage_regfile_DataPath_addr_w_p[2]) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_W_U7 ( .A(dp_id_stage_p_addr_wRD[2]), .ZN(dp_id_stage_regfile_DataPath_Conv_W_N5) );
  INV_X1 dp_id_stage_regfile_DataPath_Conv_W_U6 ( .A(
        dp_id_stage_regfile_DataPath_Conv_W_N1), .ZN(
        dp_id_stage_regfile_DataPath_Conv_W_n8) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Conv_W_U5 ( .A(
        dp_id_stage_p_addr_wRD[3]), .B(dp_id_stage_p_addr_wRD[2]), .Z(
        dp_id_stage_regfile_DataPath_Conv_W_n3) );
  AND2_X1 dp_id_stage_regfile_DataPath_Conv_W_U4 ( .A1(
        dp_id_stage_p_addr_wRD[4]), .A2(dp_id_stage_regfile_DataPath_Conv_W_n4), .ZN(dp_id_stage_regfile_DataPath_Conv_W_n2) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Conv_W_U3 ( .A(
        dp_id_stage_p_addr_wRD[4]), .B(dp_id_stage_regfile_DataPath_Conv_W_n4), 
        .Z(dp_id_stage_regfile_DataPath_Conv_W_n1) );
  AOI21_X1 dp_id_stage_regfile_DataPath_SF_converter_U20 ( .B1(1'b0), .B2(
        dp_id_stage_regfile_DataPath_addr_sf_in_2_), .A(1'b0), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_N1) );
  AND2_X1 dp_id_stage_regfile_DataPath_SF_converter_U19 ( .A1(1'b0), .A2(
        dp_id_stage_regfile_DataPath_SF_converter_n2), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_n4) );
  XOR2_X1 dp_id_stage_regfile_DataPath_SF_converter_U18 ( .A(1'b0), .B(
        dp_id_stage_regfile_DataPath_SF_converter_n2), .Z(
        dp_id_stage_regfile_DataPath_SF_converter_n3) );
  AND2_X1 dp_id_stage_regfile_DataPath_SF_converter_U17 ( .A1(1'b0), .A2(
        dp_id_stage_regfile_DataPath_addr_sf_in_2_), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_n2) );
  INV_X1 dp_id_stage_regfile_DataPath_SF_converter_U16 ( .A(
        dp_id_stage_regfile_DataPath_addr_sf_in_2_), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_N5) );
  AOI22_X1 dp_id_stage_regfile_DataPath_SF_converter_U15 ( .A1(
        dp_id_stage_regfile_DataPath_SF_converter_N5), .A2(
        dp_id_stage_regfile_DataPath_SF_converter_n10), .B1(
        dp_id_stage_regfile_DataPath_addr_sf_in_2_), .B2(
        dp_id_stage_regfile_DataPath_SF_converter_N1), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_n7) );
  INV_X1 dp_id_stage_regfile_DataPath_SF_converter_U14 ( .A(
        dp_id_stage_regfile_DataPath_SF_converter_n7), .ZN(
        dp_id_stage_regfile_DataPath_spill_fill_addr_2_) );
  AOI22_X1 dp_id_stage_regfile_DataPath_SF_converter_U13 ( .A1(
        dp_id_stage_regfile_DataPath_addr_sf_in_1_), .A2(
        dp_id_stage_regfile_DataPath_SF_converter_n10), .B1(
        dp_id_stage_regfile_DataPath_addr_sf_in_1_), .B2(
        dp_id_stage_regfile_DataPath_SF_converter_N1), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_n6) );
  INV_X1 dp_id_stage_regfile_DataPath_SF_converter_U12 ( .A(
        dp_id_stage_regfile_DataPath_SF_converter_n6), .ZN(
        dp_id_stage_regfile_DataPath_spill_fill_addr_1_) );
  AOI22_X1 dp_id_stage_regfile_DataPath_SF_converter_U11 ( .A1(
        dp_id_stage_regfile_DataPath_addr_sf_in_0_), .A2(
        dp_id_stage_regfile_DataPath_SF_converter_n10), .B1(
        dp_id_stage_regfile_DataPath_addr_sf_in_0_), .B2(
        dp_id_stage_regfile_DataPath_SF_converter_N1), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_n5) );
  INV_X1 dp_id_stage_regfile_DataPath_SF_converter_U10 ( .A(
        dp_id_stage_regfile_DataPath_SF_converter_n5), .ZN(
        dp_id_stage_regfile_DataPath_spill_fill_addr_0_) );
  XNOR2_X1 dp_id_stage_regfile_DataPath_SF_converter_U9 ( .A(1'b0), .B(
        dp_id_stage_regfile_DataPath_sf_wp_0_), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_n9) );
  NAND2_X1 dp_id_stage_regfile_DataPath_SF_converter_U8 ( .A1(
        dp_id_stage_regfile_DataPath_SF_converter_n1), .A2(
        dp_id_stage_regfile_DataPath_SF_converter_n10), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_n8) );
  OAI21_X1 dp_id_stage_regfile_DataPath_SF_converter_U7 ( .B1(
        dp_id_stage_regfile_DataPath_SF_converter_n9), .B2(
        dp_id_stage_regfile_DataPath_SF_converter_n10), .A(
        dp_id_stage_regfile_DataPath_SF_converter_n8), .ZN(
        dp_id_stage_regfile_DataPath_spill_fill_addr_3_) );
  INV_X1 dp_id_stage_regfile_DataPath_SF_converter_U6 ( .A(
        dp_id_stage_regfile_DataPath_SF_converter_N1), .ZN(
        dp_id_stage_regfile_DataPath_SF_converter_n10) );
  XOR2_X1 dp_id_stage_regfile_DataPath_SF_converter_U5 ( .A(1'b0), .B(
        dp_id_stage_regfile_DataPath_addr_sf_in_2_), .Z(
        dp_id_stage_regfile_DataPath_SF_converter_n1) );
  AND2_X1 dp_id_stage_regfile_DataPath_SF_converter_U4 ( .A1(
        dp_id_stage_regfile_DataPath_SF_converter_n3), .A2(
        dp_id_stage_regfile_DataPath_SF_converter_n10), .ZN(
        dp_id_stage_regfile_DataPath_spill_fill_addr_4_) );
  AND2_X1 dp_id_stage_regfile_DataPath_SF_converter_U3 ( .A1(
        dp_id_stage_regfile_DataPath_SF_converter_n4), .A2(
        dp_id_stage_regfile_DataPath_SF_converter_n10), .ZN(
        dp_id_stage_regfile_DataPath_spill_fill_addr_5_) );
  INV_X1 dp_id_stage_regfile_DataPath_Cwp_counter_U6 ( .A(1'b0), .ZN(
        dp_id_stage_regfile_DataPath_Cwp_counter_n2) );
  INV_X1 dp_id_stage_regfile_DataPath_Cwp_counter_U5 ( .A(
        dp_id_stage_regfile_rst_swp), .ZN(
        dp_id_stage_regfile_DataPath_Cwp_counter_n4) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Cwp_counter_U4 ( .A1(
        dp_id_stage_regfile_DataPath_Cwp_counter_n3), .A2(
        dp_id_stage_regfile_DataPath_Cwp_counter_n2), .B1(1'b0), .B2(1'b0), 
        .ZN(dp_id_stage_regfile_DataPath_Cwp_counter_n1) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Cwp_counter_U3 ( .A1(
        dp_id_stage_regfile_DataPath_Cwp_counter_n1), .A2(
        dp_id_stage_regfile_DataPath_Cwp_counter_n4), .ZN(
        dp_id_stage_regfile_DataPath_Cwp_counter_n5) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Cwp_counter_U7 ( .A(
        dp_id_stage_regfile_cnt_cwp), .B(dp_id_stage_regfile_DataPath_CWP_0_), 
        .Z(dp_id_stage_regfile_DataPath_Cwp_counter_n3) );
  DFF_X1 dp_id_stage_regfile_DataPath_Cwp_counter_Q_reg_0_ ( .D(
        dp_id_stage_regfile_DataPath_Cwp_counter_n5), .CK(CLK), .Q(
        dp_id_stage_regfile_DataPath_CWP_0_) );
  INV_X1 dp_id_stage_regfile_DataPath_Swp_counter_U6 ( .A(1'b0), .ZN(
        dp_id_stage_regfile_DataPath_Swp_counter_n2) );
  INV_X1 dp_id_stage_regfile_DataPath_Swp_counter_U5 ( .A(
        dp_id_stage_regfile_rst_swp), .ZN(
        dp_id_stage_regfile_DataPath_Swp_counter_n4) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Swp_counter_U4 ( .A1(
        dp_id_stage_regfile_DataPath_Swp_counter_n7), .A2(
        dp_id_stage_regfile_DataPath_Swp_counter_n2), .B1(1'b0), .B2(1'b0), 
        .ZN(dp_id_stage_regfile_DataPath_Swp_counter_n8) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Swp_counter_U3 ( .A1(
        dp_id_stage_regfile_DataPath_Swp_counter_n8), .A2(
        dp_id_stage_regfile_DataPath_Swp_counter_n4), .ZN(
        dp_id_stage_regfile_DataPath_Swp_counter_n6) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Swp_counter_U7 ( .A(
        dp_id_stage_regfile_cnt_swp), .B(
        dp_id_stage_regfile_DataPath_Swp_counter_Q_0_), .Z(
        dp_id_stage_regfile_DataPath_Swp_counter_n7) );
  DFF_X1 dp_id_stage_regfile_DataPath_Swp_counter_Q_reg_0_ ( .D(
        dp_id_stage_regfile_DataPath_Swp_counter_n6), .CK(CLK), .Q(
        dp_id_stage_regfile_DataPath_Swp_counter_Q_0_) );
  INV_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U18 ( .A(1'b0), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n4) );
  XNOR2_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U17 ( .A(1'b1), .B(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n11), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n10) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U16 ( .A1(
        dp_id_stage_regfile_DataPath_addr_sf_in_1_), .A2(
        dp_id_stage_regfile_DataPath_addr_sf_in_0_), .B1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n11), .B2(1'b1), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n9) );
  XNOR2_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U15 ( .A(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n9), .B(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n10), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n7) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U14 ( .A1(1'b0), 
        .A2(1'b0), .B1(dp_id_stage_regfile_DataPath_Spill_fill_counter_n1), 
        .B2(dp_id_stage_regfile_DataPath_Spill_fill_counter_n4), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n18) );
  OR2_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U13 ( .A1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n14), .A2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n18), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n17) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U12 ( .A1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n1), .A2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n12), .B1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n16), .B2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n17), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n21) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U11 ( .A1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n10), .A2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n4), .B1(1'b0), .B2(
        1'b0), .ZN(dp_id_stage_regfile_DataPath_Spill_fill_counter_n15) );
  OR2_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U10 ( .A1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n14), .A2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n15), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n13) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U9 ( .A1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n3), .A2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n12), .B1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n16), .B2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n13), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n20) );
  OAI21_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U8 ( .B1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n7), .B2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n2), .A(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n8), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n6) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U7 ( .A1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n6), .A2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n4), .B1(1'b0), .B2(
        1'b0), .ZN(dp_id_stage_regfile_DataPath_Spill_fill_counter_n5) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U6 ( .A1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n2), .A2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n12), .B1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n5), .B2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n16), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n19) );
  NOR3_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U5 ( .A1(
        dp_id_stage_regfile_rf_enable), .A2(1'b0), .A3(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n16), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n14) );
  INV_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U4 ( .A(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n14), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n12) );
  INV_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U3 ( .A(
        dp_id_stage_regfile_rst_spill_fill), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n16) );
  XOR2_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U23 ( .A(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n3), .B(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n1), .Z(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n11) );
  NAND3_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_U22 ( .A1(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n7), .A2(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n2), .A3(
        dp_id_stage_regfile_rf_enable), .ZN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n8) );
  DFF_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_Q_reg_2_ ( .D(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n19), .CK(CLK), .Q(
        dp_id_stage_regfile_DataPath_addr_sf_in_2_), .QN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n2) );
  DFF_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_Q_reg_1_ ( .D(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n20), .CK(CLK), .Q(
        dp_id_stage_regfile_DataPath_addr_sf_in_1_), .QN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n3) );
  DFF_X1 dp_id_stage_regfile_DataPath_Spill_fill_counter_Q_reg_0_ ( .D(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n21), .CK(CLK), .Q(
        dp_id_stage_regfile_DataPath_addr_sf_in_0_), .QN(
        dp_id_stage_regfile_DataPath_Spill_fill_counter_n1) );
  INV_X1 dp_id_stage_regfile_DataPath_CANSAVE_counter_U6 ( .A(
        dp_id_stage_regfile_rst_rf), .ZN(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n4) );
  AOI22_X1 dp_id_stage_regfile_DataPath_CANSAVE_counter_U5 ( .A1(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n7), .A2(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n4), .B1(
        dp_id_stage_regfile_rst_rf), .B2(1'b0), .ZN(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n8) );
  INV_X1 dp_id_stage_regfile_DataPath_CANSAVE_counter_U4 ( .A(1'b1), .ZN(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n2) );
  NOR2_X1 dp_id_stage_regfile_DataPath_CANSAVE_counter_U3 ( .A1(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n8), .A2(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n2), .ZN(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n6) );
  XOR2_X1 dp_id_stage_regfile_DataPath_CANSAVE_counter_U7 ( .A(
        dp_id_stage_regfile_cnt_save), .B(dp_id_stage_regfile_cansave), .Z(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n7) );
  DFF_X1 dp_id_stage_regfile_DataPath_CANSAVE_counter_Q_reg_0_ ( .D(
        dp_id_stage_regfile_DataPath_CANSAVE_counter_n6), .CK(CLK), .Q(
        dp_id_stage_regfile_cansave) );
  INV_X1 dp_id_stage_regfile_DataPath_CANRESTORE_counter_U6 ( .A(1'b0), .ZN(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n2) );
  INV_X1 dp_id_stage_regfile_DataPath_CANRESTORE_counter_U5 ( .A(
        dp_id_stage_regfile_rst_swp), .ZN(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n4) );
  AOI22_X1 dp_id_stage_regfile_DataPath_CANRESTORE_counter_U4 ( .A1(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n7), .A2(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n2), .B1(1'b0), .B2(
        1'b0), .ZN(dp_id_stage_regfile_DataPath_CANRESTORE_counter_n8) );
  NOR2_X1 dp_id_stage_regfile_DataPath_CANRESTORE_counter_U3 ( .A1(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n8), .A2(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n4), .ZN(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n6) );
  XOR2_X1 dp_id_stage_regfile_DataPath_CANRESTORE_counter_U7 ( .A(
        dp_id_stage_regfile_cnt_save), .B(dp_id_stage_regfile_canrestore), .Z(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n7) );
  DFF_X1 dp_id_stage_regfile_DataPath_CANRESTORE_counter_Q_reg_0_ ( .D(
        dp_id_stage_regfile_DataPath_CANRESTORE_counter_n6), .CK(CLK), .Q(
        dp_id_stage_regfile_canrestore) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_rd_U13 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_2_), .A2(
        dp_id_stage_regfile_DataPath_Mux_rd_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_rd1_p[2]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd_n11) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd_U12 ( .A(
        dp_id_stage_regfile_DataPath_Mux_rd_n11), .ZN(
        dp_id_stage_regfile_DataPath_mux_rd_out[2]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_rd_U11 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_4_), .A2(
        dp_id_stage_regfile_DataPath_Mux_rd_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_rd1_p[4]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd_n9) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd_U10 ( .A(
        dp_id_stage_regfile_DataPath_Mux_rd_n9), .ZN(
        dp_id_stage_regfile_DataPath_mux_rd_out[4]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_rd_U9 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_5_), .A2(
        dp_id_stage_regfile_DataPath_Mux_rd_n1), .B1(
        dp_id_stage_regfile_cpu_work), .B2(
        dp_id_stage_regfile_DataPath_addr_rd1_p[5]), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd_n8) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd_U8 ( .A(
        dp_id_stage_regfile_DataPath_Mux_rd_n8), .ZN(
        dp_id_stage_regfile_DataPath_mux_rd_out[5]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_rd_U7 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_3_), .A2(
        dp_id_stage_regfile_DataPath_Mux_rd_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_rd1_p[3]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd_n10) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd_U6 ( .A(
        dp_id_stage_regfile_DataPath_Mux_rd_n10), .ZN(
        dp_id_stage_regfile_DataPath_mux_rd_out[3]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_rd_U5 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_1_), .A2(
        dp_id_stage_regfile_DataPath_Mux_rd_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_rd1_p[1]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd_n12) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd_U4 ( .A(
        dp_id_stage_regfile_DataPath_Mux_rd_n12), .ZN(
        dp_id_stage_regfile_DataPath_mux_rd_out[1]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_rd_U3 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_0_), .A2(
        dp_id_stage_regfile_DataPath_Mux_rd_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_rd1_p[0]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd_n13) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd_U2 ( .A(
        dp_id_stage_regfile_DataPath_Mux_rd_n13), .ZN(
        dp_id_stage_regfile_DataPath_mux_rd_out[0]) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd_U1 ( .A(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd_n1) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_wr_U13 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_3_), .A2(
        dp_id_stage_regfile_DataPath_Mux_wr_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_w_p[3]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_n5) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_U12 ( .A(
        dp_id_stage_regfile_DataPath_Mux_wr_n5), .ZN(
        dp_id_stage_regfile_DataPath_mux_wr_out[3]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_wr_U11 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_5_), .A2(
        dp_id_stage_regfile_DataPath_Mux_wr_n1), .B1(
        dp_id_stage_regfile_cpu_work), .B2(
        dp_id_stage_regfile_DataPath_addr_w_p[5]), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_n7) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_U10 ( .A(
        dp_id_stage_regfile_DataPath_Mux_wr_n7), .ZN(
        dp_id_stage_regfile_DataPath_mux_wr_out[5]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_wr_U9 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_4_), .A2(
        dp_id_stage_regfile_DataPath_Mux_wr_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_w_p[4]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_n6) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_U8 ( .A(
        dp_id_stage_regfile_DataPath_Mux_wr_n6), .ZN(
        dp_id_stage_regfile_DataPath_mux_wr_out[4]) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_wr_U7 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_1_), .A2(
        dp_id_stage_regfile_DataPath_Mux_wr_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_w_p[1]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_n3) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_wr_U6 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_0_), .A2(
        dp_id_stage_regfile_DataPath_Mux_wr_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_w_p[0]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_n2) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_wr_U5 ( .A1(
        dp_id_stage_regfile_DataPath_spill_fill_addr_2_), .A2(
        dp_id_stage_regfile_DataPath_Mux_wr_n1), .B1(
        dp_id_stage_regfile_DataPath_addr_w_p[2]), .B2(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_n4) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_U4 ( .A(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_n1) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_U3 ( .A(
        dp_id_stage_regfile_DataPath_Mux_wr_n4), .ZN(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_U2 ( .A(
        dp_id_stage_regfile_DataPath_Mux_wr_n3), .ZN(
        dp_id_stage_regfile_DataPath_mux_wr_out[1]) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_U1 ( .A(
        dp_id_stage_regfile_DataPath_Mux_wr_n2), .ZN(
        dp_id_stage_regfile_DataPath_mux_wr_out[0]) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_sf_U3 ( .A(
        dp_id_stage_regfile_sel_wp), .ZN(
        dp_id_stage_regfile_DataPath_Mux_sf_n1) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_sf_U2 ( .A1(
        dp_id_stage_regfile_DataPath_CWP_0_), .A2(
        dp_id_stage_regfile_DataPath_Mux_sf_n1), .B1(
        dp_id_stage_regfile_sel_wp), .B2(dp_id_stage_regfile_DataPath_cwp_1_0_), .ZN(dp_id_stage_regfile_DataPath_Mux_sf_n3) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_sf_U1 ( .A(
        dp_id_stage_regfile_DataPath_Mux_sf_n3), .ZN(
        dp_id_stage_regfile_DataPath_sf_wp_0_) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd1_control_U3 ( .A(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd1_control_n2) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_rd1_control_U2 ( .A1(
        dp_id_stage_regfile_rd_cu), .A2(
        dp_id_stage_regfile_DataPath_Mux_rd1_control_n2), .B1(
        dp_id_stage_regfile_cpu_work), .B2(rf_rs1_en_i), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd1_control_n3) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd1_control_U1 ( .A(
        dp_id_stage_regfile_DataPath_Mux_rd1_control_n3), .ZN(
        dp_id_stage_regfile_DataPath_mux_rd1_control_out) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd2_control_U3 ( .A(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd2_control_n2) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_rd2_control_U2 ( .A1(1'b0), .A2(
        dp_id_stage_regfile_DataPath_Mux_rd2_control_n2), .B1(
        dp_id_stage_regfile_cpu_work), .B2(rf_rs2_en_i), .ZN(
        dp_id_stage_regfile_DataPath_Mux_rd2_control_n4) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_rd2_control_U1 ( .A(
        dp_id_stage_regfile_DataPath_Mux_rd2_control_n4), .ZN(
        dp_id_stage_regfile_DataPath_mux_rd2_control_out) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_wr_control_U3 ( .A1(
        dp_id_stage_regfile_wr_cu), .A2(
        dp_id_stage_regfile_DataPath_Mux_wr_control_n2), .B1(
        dp_id_stage_regfile_cpu_work), .B2(rf_we_i), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_control_n4) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_control_U2 ( .A(
        dp_id_stage_regfile_DataPath_Mux_wr_control_n4), .ZN(
        dp_id_stage_regfile_DataPath_mux_wr_control_out) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_wr_control_U1 ( .A(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_wr_control_n2) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_en_control_U3 ( .A(
        dp_id_stage_regfile_cpu_work), .ZN(
        dp_id_stage_regfile_DataPath_Mux_en_control_n2) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Mux_en_control_U2 ( .A1(
        dp_id_stage_regfile_rf_enable), .A2(
        dp_id_stage_regfile_DataPath_Mux_en_control_n2), .B1(
        dp_id_stage_regfile_cpu_work), .B2(1'b1), .ZN(
        dp_id_stage_regfile_DataPath_Mux_en_control_n4) );
  INV_X1 dp_id_stage_regfile_DataPath_Mux_en_control_U1 ( .A(
        dp_id_stage_regfile_DataPath_Mux_en_control_n4), .ZN(
        dp_id_stage_regfile_DataPath_mux_en_control_out) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3825 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4227), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3824 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4217), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3823 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4207), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3822 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4144), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3821 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4134), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3820 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4124), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3819 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4114), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3818 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4042), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3817 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4032), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3816 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3982), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3815 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3950), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3814 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3900), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3813 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3890), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3812 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1189), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1188) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3811 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1189), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3810 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1189), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3809 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1189), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1185) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3808 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1200), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3807 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1200), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3806 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1200), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3805 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1200), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3804 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1200), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3803 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1200), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1179) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3802 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1202), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3801 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1202), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3800 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1202), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1176) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3799 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1202), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3798 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1202), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3797 ( .A1(
        dp_id_stage_regfile_DataPath_mux_rd2_control_out), .A2(
        dp_id_stage_regfile_DataPath_mux_en_control_out), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N429) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3796 ( .A1(
        dp_id_stage_regfile_DataPath_mux_rd1_control_out), .A2(
        dp_id_stage_regfile_DataPath_mux_en_control_out), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N428) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3795 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n450), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n418), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2553), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2541) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3794 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2523), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2524), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2525), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2526), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2522) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3793 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2541), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2542), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2543), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2544), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2521) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3792 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2521), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2522), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N396) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3791 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n450), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n418), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3180), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3168) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3790 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3150), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3151), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3152), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3153), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3149) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3789 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3168), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3169), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3170), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3171), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3148) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3788 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3148), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3149), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N328) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3787 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n451), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n419), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2520), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2513) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3786 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2505), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2506), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2507), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2508), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2504) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3785 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2513), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2514), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2515), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2516), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2503) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3784 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2503), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2504), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N397) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3783 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n451), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n419), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3147), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3140) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3782 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3132), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3133), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3134), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3135), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3131) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3781 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3140), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3141), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3142), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3143), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3130) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3780 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3130), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3131), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N329) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3779 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n452), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n420), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2502), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2495) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3778 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2487), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2488), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2489), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2490), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2486) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3777 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2495), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2496), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2497), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2498), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2485) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3776 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2485), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2486), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N398) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3775 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n452), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n420), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3129), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3122) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3774 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3114), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3115), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3116), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3117), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3113) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3773 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3122), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3123), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3124), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3125), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3112) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3772 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3112), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3113), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N330) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3771 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n453), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n421), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2484), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2477) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3770 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2469), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2470), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2471), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2472), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2468) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3769 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2477), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2478), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2479), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2480), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2467) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3768 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2467), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2468), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N399) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3767 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n453), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n421), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3111), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3104) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3766 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3096), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3097), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3098), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3099), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3095) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3765 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3104), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3105), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3106), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3107), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3094) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3764 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3094), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3095), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N331) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3763 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n454), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n422), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2466), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2459) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3762 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2451), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2452), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2453), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2454), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2450) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3761 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2459), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2460), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2461), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2462), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2449) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3760 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2449), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2450), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N400) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3759 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n454), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n422), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3093), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3086) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3758 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3078), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3079), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3080), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3081), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3077) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3757 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3086), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3087), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3088), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3089), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3076) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3756 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3076), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3077), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N332) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3755 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n455), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n423), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2448), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2441) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3754 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2433), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2434), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2435), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2436), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2432) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3753 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2441), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2442), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2443), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2444), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2431) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3752 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2431), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2432), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N401) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3751 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n455), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n423), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3075), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3068) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3750 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3060), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3061), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3062), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3063), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3059) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3749 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3068), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3069), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3070), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3071), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3058) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3748 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3058), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3059), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N333) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3747 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n456), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n424), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2430), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2423) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3746 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2415), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2416), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2417), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2418), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2414) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3745 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2423), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2424), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2425), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2426), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2413) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3744 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2413), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2414), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N402) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3743 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n456), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n424), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3057), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3050) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3742 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3042), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3043), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3044), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3045), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3041) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3741 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3050), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3051), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3052), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3053), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3040) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3740 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3040), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3041), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N334) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3739 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n457), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n425), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2412), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2405) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3738 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2397), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2398), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2399), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2400), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2396) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3737 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2405), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2406), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2407), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2408), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2395) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3736 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2395), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2396), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N403) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3735 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n457), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n425), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3039), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3032) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3734 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3024), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3025), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3026), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3027), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3023) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3733 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3032), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3033), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3034), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3035), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3022) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3732 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3022), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3023), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N335) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3731 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n458), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n426), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2394), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2387) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3730 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2379), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2380), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2381), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2382), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2378) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3729 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2387), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2388), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2389), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2390), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2377) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3728 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2377), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2378), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N404) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3727 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n458), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n426), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3021), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3014) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3726 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3006), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3007), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3008), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3009), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3005) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3725 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3014), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3015), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n3016), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n3017), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3004) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3724 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3004), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3005), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N336) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3723 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n459), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n427), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2376), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2369) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3722 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2361), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2362), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2363), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2364), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2360) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3721 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2369), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2370), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2371), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2372), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2359) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3720 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2359), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2360), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N405) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3719 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n459), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n427), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3003), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2996) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3718 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2988), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2989), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2990), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2991), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2987) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3717 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2996), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2997), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2998), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2999), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2986) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3716 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2986), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2987), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N337) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3715 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n460), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n428), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2358), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2351) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3714 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2344), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2345), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2346), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2342) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3713 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2351), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2352), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2353), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2354), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2341) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3712 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2341), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2342), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N406) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3711 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n460), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n428), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2985), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2978) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3710 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2970), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2971), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2972), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2973), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2969) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3709 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2978), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2979), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2980), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2981), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2968) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3708 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2968), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2969), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N338) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3707 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n461), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n429), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2340), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2333) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3706 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2325), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2326), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2327), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2328), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2324) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3705 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2333), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2334), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2335), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2336), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2323) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3704 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2323), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2324), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N407) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3703 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n461), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n429), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2967), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2960) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3702 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2952), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2953), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2954), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2955), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2951) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3701 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2960), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2961), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2962), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2963), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2950) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3700 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2950), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2951), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N339) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3699 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n462), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n430), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2322), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2315) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3698 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2307), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2308), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2309), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2310), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2306) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3697 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2315), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2316), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2317), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2318), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2305) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3696 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2305), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2306), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N408) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3695 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n462), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n430), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2949), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2942) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3694 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2934), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2935), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2936), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2937), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2933) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3693 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2942), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2943), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2944), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2945), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2932) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3692 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2932), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2933), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N340) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3691 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n463), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n431), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2304), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2297) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3690 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2289), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2290), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2291), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2292), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2288) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3689 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2297), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2298), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2299), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2300), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2287) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3688 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2287), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2288), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N409) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3687 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n463), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n431), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2931), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2924) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3686 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2916), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2917), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2918), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2919), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2915) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3685 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2924), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2925), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2926), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2927), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2914) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3684 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2914), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2915), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N341) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3683 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n464), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n432), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2286), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2279) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3682 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2271), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2272), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2273), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2274), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2270) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3681 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2279), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2280), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2281), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2282), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2269) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3680 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2270), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N410) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3679 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n464), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n432), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2913), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2906) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3678 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2898), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2899), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2900), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2901), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2897) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3677 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2906), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2907), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2908), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2909), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2896) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3676 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2896), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2897), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N342) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3675 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n465), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n433), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2268), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2261) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3674 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2254), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2255), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2256), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2252) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3673 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2262), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2263), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2264), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2251) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3672 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2252), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N411) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3671 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n465), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n433), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2895), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2888) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3670 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2880), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2881), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2882), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2883), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2879) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3669 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2888), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2889), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2890), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2891), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2878) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3668 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2878), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2879), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N343) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3667 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n466), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n434), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2250), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2243) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3666 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2235), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2236), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2237), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2238), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2234) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3665 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2244), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2245), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2246), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2233) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3664 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2233), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2234), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N412) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3663 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n466), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n434), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2877), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2870) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3662 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2862), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2863), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2864), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2865), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2861) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3661 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2870), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2871), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2872), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2873), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2860) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3660 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2860), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2861), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N344) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3659 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n467), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n435), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2232), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2225) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3658 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2217), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2218), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2219), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2220), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2216) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3657 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2225), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2226), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2227), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2228), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2215) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3656 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2215), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2216), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N413) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3655 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n467), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n435), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2859), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2852) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3654 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2844), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2845), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2846), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2847), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2843) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3653 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2853), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2854), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2855), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2842) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3652 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2842), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2843), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N345) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3651 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n468), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n436), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2214), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2207) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3650 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2199), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2200), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2201), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2202), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2198) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3649 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2207), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2208), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2209), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2210), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2197) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3648 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2197), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2198), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N414) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3647 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n468), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n436), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2841), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2834) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3646 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2826), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2827), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2828), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2829), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2825) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3645 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2834), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2835), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2836), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2837), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2824) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3644 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2825), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N346) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3643 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n469), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n437), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2196), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2189) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3642 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2181), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2182), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2183), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2184), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2180) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3641 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2189), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2190), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2191), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2192), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2179) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3640 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2179), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2180), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N415) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3639 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n469), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n437), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2823), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2816) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3638 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2808), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2809), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2810), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2811), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2807) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3637 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2816), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2817), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2818), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2819), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2806) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3636 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2806), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2807), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N347) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3635 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n470), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n438), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2178), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2171) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3634 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2163), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2164), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2165), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2166), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2162) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3633 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2171), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2172), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2173), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2174), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2161) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3632 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2161), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2162), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N416) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3631 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n470), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n438), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2805), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2798) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3630 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2790), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2791), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2792), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2793), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2789) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3629 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2799), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2800), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2801), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2788) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3628 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2788), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2789), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N348) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3627 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n471), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n439), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2153) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3626 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2145), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2146), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2147), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2148), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2144) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3625 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2153), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2154), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2155), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2143) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3624 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2143), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2144), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N417) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3623 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n471), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n439), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2787), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2780) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3622 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2772), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2773), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2774), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2775), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2771) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3621 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2780), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2781), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2782), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2783), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2770) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3620 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2771), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N349) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3619 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n472), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n440), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2142), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2135) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3618 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2127), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2128), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2129), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2130), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2126) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3617 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2135), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2136), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2137), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2138), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2125) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3616 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2125), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2126), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N418) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3615 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n472), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n440), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2769), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2762) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3614 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2754), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2755), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2756), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2757), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2753) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3613 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2762), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2763), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2764), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2765), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2752) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3612 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2752), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2753), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N350) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3611 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n473), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n441), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2124), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2117) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3610 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2109), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2110), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2111), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2112), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2108) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3609 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2117), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2118), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2119), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2120), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2107) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3608 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2107), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2108), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N419) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3607 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n473), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n441), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2751), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2744) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3606 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2736), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2737), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2738), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2739), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2735) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3605 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2745), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2746), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2747), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2734) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3604 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2734), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2735), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N351) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3603 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n474), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n442), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2106), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2099) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3602 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2091), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2092), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2093), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2094), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2090) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3601 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2099), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2100), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2101), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2102), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2089) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3600 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2089), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2090), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N420) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3599 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n474), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n442), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2733), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2726) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3598 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2718), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2719), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2720), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2721), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2717) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3597 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2726), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2727), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2728), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2729), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2716) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3596 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2717), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N352) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3595 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n475), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n443), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2088), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2081) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3594 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2073), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2074), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2075), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2076), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2072) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3593 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2081), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2082), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2083), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2084), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2071) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3592 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2071), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2072), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N421) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3591 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n475), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n443), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2715), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2708) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3590 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2700), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2701), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2702), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2703), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2699) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3589 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2708), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2709), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2710), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2711), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2698) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3588 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2698), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2699), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N353) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3587 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n476), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n444), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2070), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2063) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3586 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2055), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2056), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2057), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2058), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2054) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3585 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2063), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2064), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2065), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2066), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2053) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3584 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2053), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2054), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N422) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3583 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n476), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n444), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2697), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2690) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3582 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2682), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2683), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2684), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2685), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2681) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3581 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2690), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2691), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2692), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2693), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2680) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3580 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2680), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2681), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N354) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3579 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n477), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n445), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2052), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2045) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3578 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2037), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2038), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2039), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2040), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2036) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3577 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2045), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2046), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2047), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2048), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2035) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3576 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2035), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2036), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N423) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3575 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n477), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n445), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2679), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2672) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3574 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2664), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2665), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2666), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2667), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2663) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3573 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2672), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2673), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2674), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2675), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2662) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3572 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2662), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2663), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N355) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3571 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n478), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n446), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2034), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2027) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3570 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2019), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2020), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2021), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2022), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2018) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3569 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2027), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2028), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2029), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2030), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2017) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3568 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2017), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2018), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N424) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3567 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n478), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n446), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2661), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2654) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3566 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2646), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2647), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2648), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2649), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2645) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3565 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2654), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2655), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2656), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2657), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2644) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3564 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2644), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2645), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N356) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3563 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n479), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n447), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2016), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2009) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3562 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2001), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2002), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2003), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2004), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2000) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3561 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2009), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2010), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2011), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2012), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1999) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3560 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1999), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2000), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N425) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3559 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n479), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n447), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2643), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2636) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3558 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2628), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2629), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2630), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2631), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2627) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3557 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2636), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2637), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2638), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2639), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2626) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3556 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2626), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2627), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N357) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3555 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n480), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n448), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1998), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1991) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3554 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1983), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1984), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1985), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1986), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1982) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3553 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1991), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1992), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1993), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1994), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1981) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3552 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1981), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1982), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N426) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3551 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n480), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n448), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2625), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2618) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3550 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2610), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2611), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2612), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2613), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2609) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3549 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2618), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2619), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2620), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2621), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2608) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3548 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2608), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2609), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N358) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3547 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n481), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n449), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1977), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1955) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3546 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1929), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1930), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1931), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1932), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1928) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3545 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1955), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1956), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1957), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1958), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1927) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3544 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1927), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1928), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N427) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3543 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n481), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n449), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2604), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2582) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3542 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2556), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2557), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2558), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2559), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2555) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3541 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2582), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2583), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n2584), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n2585), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2554) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3540 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2554), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2555), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_N359) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3539 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__31_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2540) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3538 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1026), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n994), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2540), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2523) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3537 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__31_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3167) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3536 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1026), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n994), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3167), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3150) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3535 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__30_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2512) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3534 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1027), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n995), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2512), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2505) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3533 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__30_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3139) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3532 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1027), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n995), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3139), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3132) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3531 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__29_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2494) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3530 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1028), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n996), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2494), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2487) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3529 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__29_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3121) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3528 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1028), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n996), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3121), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3114) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3527 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__28_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2476) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3526 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1029), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n997), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2476), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2469) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3525 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__28_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3103) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3524 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1029), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n997), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3103), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3096) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3523 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__27_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2458) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3522 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1030), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n998), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2458), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2451) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3521 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__27_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3085) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3520 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1030), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n998), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3085), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3078) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3519 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__26_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2440) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3518 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1031), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n999), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2440), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2433) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3517 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__26_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3067) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3516 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1031), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n999), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3067), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3060) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3515 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__25_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2422) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3514 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1032), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1000), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2422), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2415) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3513 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__25_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3049) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3512 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1032), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1000), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3049), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3042) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3511 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__24_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2404) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3510 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1033), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1001), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2404), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2397) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3509 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__24_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3031) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3508 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1033), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1001), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3031), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3024) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3507 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__23_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2386) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3506 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1034), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1002), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2386), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2379) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3505 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__23_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3013) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3504 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1034), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1002), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3013), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3006) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3503 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__22_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2368) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3502 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1035), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1003), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2368), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2361) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3501 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__22_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2995) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3500 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1035), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1003), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2995), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2988) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3499 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__21_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2350) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3498 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1036), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1004), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2350), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2343) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3497 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__21_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2977) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3496 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1036), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1004), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2977), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2970) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3495 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__20_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2332) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3494 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1037), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1005), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2332), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2325) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3493 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__20_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2959) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3492 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1037), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1005), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2959), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2952) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3491 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__19_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2314) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3490 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1038), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1006), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2314), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2307) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3489 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__19_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2941) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3488 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1038), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1006), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2941), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2934) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3487 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__18_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2296) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3486 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1039), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1007), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2296), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2289) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3485 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__18_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2923) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3484 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1039), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1007), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2923), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2916) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3483 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__17_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2278) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3482 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1040), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1008), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2278), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2271) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3481 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__17_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2905) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3480 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1040), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1008), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2905), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2898) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3479 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__16_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2260) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3478 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1041), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1009), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2260), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2253) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3477 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__16_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2887) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3476 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1041), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1009), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2887), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2880) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3475 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__15_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2242) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3474 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1042), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1010), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2242), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2235) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3473 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__15_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2869) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3472 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1042), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1010), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2869), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2862) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3471 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__14_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2224) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3470 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1043), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1011), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2224), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2217) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3469 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__14_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2851) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3468 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1043), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1011), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2851), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2844) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3467 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__13_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2206) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3466 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1044), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1012), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2206), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2199) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3465 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__13_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2833) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3464 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1044), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1012), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2833), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2826) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3463 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__12_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2188) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3462 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1045), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1013), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2188), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2181) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3461 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__12_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2815) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3460 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1045), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1013), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2815), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2808) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3459 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__11_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2170) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3458 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1046), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1014), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2170), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2163) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3457 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__11_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2797) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3456 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1046), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1014), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2797), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2790) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3455 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__10_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2152) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3454 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1047), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1015), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2152), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2145) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3453 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__10_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2779) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3452 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1047), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1015), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2779), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2772) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3451 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__9_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2134) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3450 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1048), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1016), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2134), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2127) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3449 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__9_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2761) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3448 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1048), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1016), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2761), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2754) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3447 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__8_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2116) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3446 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1049), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1017), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2116), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2109) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3445 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__8_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2743) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3444 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1049), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1017), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2743), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2736) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3443 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__7_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2098) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3442 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1050), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1018), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2098), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2091) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3441 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__7_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2725) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3440 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1050), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1018), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2725), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2718) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3439 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__6_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2080) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3438 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1051), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1019), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2080), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2073) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3437 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__6_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2707) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3436 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1051), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1019), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2707), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2700) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3435 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__5_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2062) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3434 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1052), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1020), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2062), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2055) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3433 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__5_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2689) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3432 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1052), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1020), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2689), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2682) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3431 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__4_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2044) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3430 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1053), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1021), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2044), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2037) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3429 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__4_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2671) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3428 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1053), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1021), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2671), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2664) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3427 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__3_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2026) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3426 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1054), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1022), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2026), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2019) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3425 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__3_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2653) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3424 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1054), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1022), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2653), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2646) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3423 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__2_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2008) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3422 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1055), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1023), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2008), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2001) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3421 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__2_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2635) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3420 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1055), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1023), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2635), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2628) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3419 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__1_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1990) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3418 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1056), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1024), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1990), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1983) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3417 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__1_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2617) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3416 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1056), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1024), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2617), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2610) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3415 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__0_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1951) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3414 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1057), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1025), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1951), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1929) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3413 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__0_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2578) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3412 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1057), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1025), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2578), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2556) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3411 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2550) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3410 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n322), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n290), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2550), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2542) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3409 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2537) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3408 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n962), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n930), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2537), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2524) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3407 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3177) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3406 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n322), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n290), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3177), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3169) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3405 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3164) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3404 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n962), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n930), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3164), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3151) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3403 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2519) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3402 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n323), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n291), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2519), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2514) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3401 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2511) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3400 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n963), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n931), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2511), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2506) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3399 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3146) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3398 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n323), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n291), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3146), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3141) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3397 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3138) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3396 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n963), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n931), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3138), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3133) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3395 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2501) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3394 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n324), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n292), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2501), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2496) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3393 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2493) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3392 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n964), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n932), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2493), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2488) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3391 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3128) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3390 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n324), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n292), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3128), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3123) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3389 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3120) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3388 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n964), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n932), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3120), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3115) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3387 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2483) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3386 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n325), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n293), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2483), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2478) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3385 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2475) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3384 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n965), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n933), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2475), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2470) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3383 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3110) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3382 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n325), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n293), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3110), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3105) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3381 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3102) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3380 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n965), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n933), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3102), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3097) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3379 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2465) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3378 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n326), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n294), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2465), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2460) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3377 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2457) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3376 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n966), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n934), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2457), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2452) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3375 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3092) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3374 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n326), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n294), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3092), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3087) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3373 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3084) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3372 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n966), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n934), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3084), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3079) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3371 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2447) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3370 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n327), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n295), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2447), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2442) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3369 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2439) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3368 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n967), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n935), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2439), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2434) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3367 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3074) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3366 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n327), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n295), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3074), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3069) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3365 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3066) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3364 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n967), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n935), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3066), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3061) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3363 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2429) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3362 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n328), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n296), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2429), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2424) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3361 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2421) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3360 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n968), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n936), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2421), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2416) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3359 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3056) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3358 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n328), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n296), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3056), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3051) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3357 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3048) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3356 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n968), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n936), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3048), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3043) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3355 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2411) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3354 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n329), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n297), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2411), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2406) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3353 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2403) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3352 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n969), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n937), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2403), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2398) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3351 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3038) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3350 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n329), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n297), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3038), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3033) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3349 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3030) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3348 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n969), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n937), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3030), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3025) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3347 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2393) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3346 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n330), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n298), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2393), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2388) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3345 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2385) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3344 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n970), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n938), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2385), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2380) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3343 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3020) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3342 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n330), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n298), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3020), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3015) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3341 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3012) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3340 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n970), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n938), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3012), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3007) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3339 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2375) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3338 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n331), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n299), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2375), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2370) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3337 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2367) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3336 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n971), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n939), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2367), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2362) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3335 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3002) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3334 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n331), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n299), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3002), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2997) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3333 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2994) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3332 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n971), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n939), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2994), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2989) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3331 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2357) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3330 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n332), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n300), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2357), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2352) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3329 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2349) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3328 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n972), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n940), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2349), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2344) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3327 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2984) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3326 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n332), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n300), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2984), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2979) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3325 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2976) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3324 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n972), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n940), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2976), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2971) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3323 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2339) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3322 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n333), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n301), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2339), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2334) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3321 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2331) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3320 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n973), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n941), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2331), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2326) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3319 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2966) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3318 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n333), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n301), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2966), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2961) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3317 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2958) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3316 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n973), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n941), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2958), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2953) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3315 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2321) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3314 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n334), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n302), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2321), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2316) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3313 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2313) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3312 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n974), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n942), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2313), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2308) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3311 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2948) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3310 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n334), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n302), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2948), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2943) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3309 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2940) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3308 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n974), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n942), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2940), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2935) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3307 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2303) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3306 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n335), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n303), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2303), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2298) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3305 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2295) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3304 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n975), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n943), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2295), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2290) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3303 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2930) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3302 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n335), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n303), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2930), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2925) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3301 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2922) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3300 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n975), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n943), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2922), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2917) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3299 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2285) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3298 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n336), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n304), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2285), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2280) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3297 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2277) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3296 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n976), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n944), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2277), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2272) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3295 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2912) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3294 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n336), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n304), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2912), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2907) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3293 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2904) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3292 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n976), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n944), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2904), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2899) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3291 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2267) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3290 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n337), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n305), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2267), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2262) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3289 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2259) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3288 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n977), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n945), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2259), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2254) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3287 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2894) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3286 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n337), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n305), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2894), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2889) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3285 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2886) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3284 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n977), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n945), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2886), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2881) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3283 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2249) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3282 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n338), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n306), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2249), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2244) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3281 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2241) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3280 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n978), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n946), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2241), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2236) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3279 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2876) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3278 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n338), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n306), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2876), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2871) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3277 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2868) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3276 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n978), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n946), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2868), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2863) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3275 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2231) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3274 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n339), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n307), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2231), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2226) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3273 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2223) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3272 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n979), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n947), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2223), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2218) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3271 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2858) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3270 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n339), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n307), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2858), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2853) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3269 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2850) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3268 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n979), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n947), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2850), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2845) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3267 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2213) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3266 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n340), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n308), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2213), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2208) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3265 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2205) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3264 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n980), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n948), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2205), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2200) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3263 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2840) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3262 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n340), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n308), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2840), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2835) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3261 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2832) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3260 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n980), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n948), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2832), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2827) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3259 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2195) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3258 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n341), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n309), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2195), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2190) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3257 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2187) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3256 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n981), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n949), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2187), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2182) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3255 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2822) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3254 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n341), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n309), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2822), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2817) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3253 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2814) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3252 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n981), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n949), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2814), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2809) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3251 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2177) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3250 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n342), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n310), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2177), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2172) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3249 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2169) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3248 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n982), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n950), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2169), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2164) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3247 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2804) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3246 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n342), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n310), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2804), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2799) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3245 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2796) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3244 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n982), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n950), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2796), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2791) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3243 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2159) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3242 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n343), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n311), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2154) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3241 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2151) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3240 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n983), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n951), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2151), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2146) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3239 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2786) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3238 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n343), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n311), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2786), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2781) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3237 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2778) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3236 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n983), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n951), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2778), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2773) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3235 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2141) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3234 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n344), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n312), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2141), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2136) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3233 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2133) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3232 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n984), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n952), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2133), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2128) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3231 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2768) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3230 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n344), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n312), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2768), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2763) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3229 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2760) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3228 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n984), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n952), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2760), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2755) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3227 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2123) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3226 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n345), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n313), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2123), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2118) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3225 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2115) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3224 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n985), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n953), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2115), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2110) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3223 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2750) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3222 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n345), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n313), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2750), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2745) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3221 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2742) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3220 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n985), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n953), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2742), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2737) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3219 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2105) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3218 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n346), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n314), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2105), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2100) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3217 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2097) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3216 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n986), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n954), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2097), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2092) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3215 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2732) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3214 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n346), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n314), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2732), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2727) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3213 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2724) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3212 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n986), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n954), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2724), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2719) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3211 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2087) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3210 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n347), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n315), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2087), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2082) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3209 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2079) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3208 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n987), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n955), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2079), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2074) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3207 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2714) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3206 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n347), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n315), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2714), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2709) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3205 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2706) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3204 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n987), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n955), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2706), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2701) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3203 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2069) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3202 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n348), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n316), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2069), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2064) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3201 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2061) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3200 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n988), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n956), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2061), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2056) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3199 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2696) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3198 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n348), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n316), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2696), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2691) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3197 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2688) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3196 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n988), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n956), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2688), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2683) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3195 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2051) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3194 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n349), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n317), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2051), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2046) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3193 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2043) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3192 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n989), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n957), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2043), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2038) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3191 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2678) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3190 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n349), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n317), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2678), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2673) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3189 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2670) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3188 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n989), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n957), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2670), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2665) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3187 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2033) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3186 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n350), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n318), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2033), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2028) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3185 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2025) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3184 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n990), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n958), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2025), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2020) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3183 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2660) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3182 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n350), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n318), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2660), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2655) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3181 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2652) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3180 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n990), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n958), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2652), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2647) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3179 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2015) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3178 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n351), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n319), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2015), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2010) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3177 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2007) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3176 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n991), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n959), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2007), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2002) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3175 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2642) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3174 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n351), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n319), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2642), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2637) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3173 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2634) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3172 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n991), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n959), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2634), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2629) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3171 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1997) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3170 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n352), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n320), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1997), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1992) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3169 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1989) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3168 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n992), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n960), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1989), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1984) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3167 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2624) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3166 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n352), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n320), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2624), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2619) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3165 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2616) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3164 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n992), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n960), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2616), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2611) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3163 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1972) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3162 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n353), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n321), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1972), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1956) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3161 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1946) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3160 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n993), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n961), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1946), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1930) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3159 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2599) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3158 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n353), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n321), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2599), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2583) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3157 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2573) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3156 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n993), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n961), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2573), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2557) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3155 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__31_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2547) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3154 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n162), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n130), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2547), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2543) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3153 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__31_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2534) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3152 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n738), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n706), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2534), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2525) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3151 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__31_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3174) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3150 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n162), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n130), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3174), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3170) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3149 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__31_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3161) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3148 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n738), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n706), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3161), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3152) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3147 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__30_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2518) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3146 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n163), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n131), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2518), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2515) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3145 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__30_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2510) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3144 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n707), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2510), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2507) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3143 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__30_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3145) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3142 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n163), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n131), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3145), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3142) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3141 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__30_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3137) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3140 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n707), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3137), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3134) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3139 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__29_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2500) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3138 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n164), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n132), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2500), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2497) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3137 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__29_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2492) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3136 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n708), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2492), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2489) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3135 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__29_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3127) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3134 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n164), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n132), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3127), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3124) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3133 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__29_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3119) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3132 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n708), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3119), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3116) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3131 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__28_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2482) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3130 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n165), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n133), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2482), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2479) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3129 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__28_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2474) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3128 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n709), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2474), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2471) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3127 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__28_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3109) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3126 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n165), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n133), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3109), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3106) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3125 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__28_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3101) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3124 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n709), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3101), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3098) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3123 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__27_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2464) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3122 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n166), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n134), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2464), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2461) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3121 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__27_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2456) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3120 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n742), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n710), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2456), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2453) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3119 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__27_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3091) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3118 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n166), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n134), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3091), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3088) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3117 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__27_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3083) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3116 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n742), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n710), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3083), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3080) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3115 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__26_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2446) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3114 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n167), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n135), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2446), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2443) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3113 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__26_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2438) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3112 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n743), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n711), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2438), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2435) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3111 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__26_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3073) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3110 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n167), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n135), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3073), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3070) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3109 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__26_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3065) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3108 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n743), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n711), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3065), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3062) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3107 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__25_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2428) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3106 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n168), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n136), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2428), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2425) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3105 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__25_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2420) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3104 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n744), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n712), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2420), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2417) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3103 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__25_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3055) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3102 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n168), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n136), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3055), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3052) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3101 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__25_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3047) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3100 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n744), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n712), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3047), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3044) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3099 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__24_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2410) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3098 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n169), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n137), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2410), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2407) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3097 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__24_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2402) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3096 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n745), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n713), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2402), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2399) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3095 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__24_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3037) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3094 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n169), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n137), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3037), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3034) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3093 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__24_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3029) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3092 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n745), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n713), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3029), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3026) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3091 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__23_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2392) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3090 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n170), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n138), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2392), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2389) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3089 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__23_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2384) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3088 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n746), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n714), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2384), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2381) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3087 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__23_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3019) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3086 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n170), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n138), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3019), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3016) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3085 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__23_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3011) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3084 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n746), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n714), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3011), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3008) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3083 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__22_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2374) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3082 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n171), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n139), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2374), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2371) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3081 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__22_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2366) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3080 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n747), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n715), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2366), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2363) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3079 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__22_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3001) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3078 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n171), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n139), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3001), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2998) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3077 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__22_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2993) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3076 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n747), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n715), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2993), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2990) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3075 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__21_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2356) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3074 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n172), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n140), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2356), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2353) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3073 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__21_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2348) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3072 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n748), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n716), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2348), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2345) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3071 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__21_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2983) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3070 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n172), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n140), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2983), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2980) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3069 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__21_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2975) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3068 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n748), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n716), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2975), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2972) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3067 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__20_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2338) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3066 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n173), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n141), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2338), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2335) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3065 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__20_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2330) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3064 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n749), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n717), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2330), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2327) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3063 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__20_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2965) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3062 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n173), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n141), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2965), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2962) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3061 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__20_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2957) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3060 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n749), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n717), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2957), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2954) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3059 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__19_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2320) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3058 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n174), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n142), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2320), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2317) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3057 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__19_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2312) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3056 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n750), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n718), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2312), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2309) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3055 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__19_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2947) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3054 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n174), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n142), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2947), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2944) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3053 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__19_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2939) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3052 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n750), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n718), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2939), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2936) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3051 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__18_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2302) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3050 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n175), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n143), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2302), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2299) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3049 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__18_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2294) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3048 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n751), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n719), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2294), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2291) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3047 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__18_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2929) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3046 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n175), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n143), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2929), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2926) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3045 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__18_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2921) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3044 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n751), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n719), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2921), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2918) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3043 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__17_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2284) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3042 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n176), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n144), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2284), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2281) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3041 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__17_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2276) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3040 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n752), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n720), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2276), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2273) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3039 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__17_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2911) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3038 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n176), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n144), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2911), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2908) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3037 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__17_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2903) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3036 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n752), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n720), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2903), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2900) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3035 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__16_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2266) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3034 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n177), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n145), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2266), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2263) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3033 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__16_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2258) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3032 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n753), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n721), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2258), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2255) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3031 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__16_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2893) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3030 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n177), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n145), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2893), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2890) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3029 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__16_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2885) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3028 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n753), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n721), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2885), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2882) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3027 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__15_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2248) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3026 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n178), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n146), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2248), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2245) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3025 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__15_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2240) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3024 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n722), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2240), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2237) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3023 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__15_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2875) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3022 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n178), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n146), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2875), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2872) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3021 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__15_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2867) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3020 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n722), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2867), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2864) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3019 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__14_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2230) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3018 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n179), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n147), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2230), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2227) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3017 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__14_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2222) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3016 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n723), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2222), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2219) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3015 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__14_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2857) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3014 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n179), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n147), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2857), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2854) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3013 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__14_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2849) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3012 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n723), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2849), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2846) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3011 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__13_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2212) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3010 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n180), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n148), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2212), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2209) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3009 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__13_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2204) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3008 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2204), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2201) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3007 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__13_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2839) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3006 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n180), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n148), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2839), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2836) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3005 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__13_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2831) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3004 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2831), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2828) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3003 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__12_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2194) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3002 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n181), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n149), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2194), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2191) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3001 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__12_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2186) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3000 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n757), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2186), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2183) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2999 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__12_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2821) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2998 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n181), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n149), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2821), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2818) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2997 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__12_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2813) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2996 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n757), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n725), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2813), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2810) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2995 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__11_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2176) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2994 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n182), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n150), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2176), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2173) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2993 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__11_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2168) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2992 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n758), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2168), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2165) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2991 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__11_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2803) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2990 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n182), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n150), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2803), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2800) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2989 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__11_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2795) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2988 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n758), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n726), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2795), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2792) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2987 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__10_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2158) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2986 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n183), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n151), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2158), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2155) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2985 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__10_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2150) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2984 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n759), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n727), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2150), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2147) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2983 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__10_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2785) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2982 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n183), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n151), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2785), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2782) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2981 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__10_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2777) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2980 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n759), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n727), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2777), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2774) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2979 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__9_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2140) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2978 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n184), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n152), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2140), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2137) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2977 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__9_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2132) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2976 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n760), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n728), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2132), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2129) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2975 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__9_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2767) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2974 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n184), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n152), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2767), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2764) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2973 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__9_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2759) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2972 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n760), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n728), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2759), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2756) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2971 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__8_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2122) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2970 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n185), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n153), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2122), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2119) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2969 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__8_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2114) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2968 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n761), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n729), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2114), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2111) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2967 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__8_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2749) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2966 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n185), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n153), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2749), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2746) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2965 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__8_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2741) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2964 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n761), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n729), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2741), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2738) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2963 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__7_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2104) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2962 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n186), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n154), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2104), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2101) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2961 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__7_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2096) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2960 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n762), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n730), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2096), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2093) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2959 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__7_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2731) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2958 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n186), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n154), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2731), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2728) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2957 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__7_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2723) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2956 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n762), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n730), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2723), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2720) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2955 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__6_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2086) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2954 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n187), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n155), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2086), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2083) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2953 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__6_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2078) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2952 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n763), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n731), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2078), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2075) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2951 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__6_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2713) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2950 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n187), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n155), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2713), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2710) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2949 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__6_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2705) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2948 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n763), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n731), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2705), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2702) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2947 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__5_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2068) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2946 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n188), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n156), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2068), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2065) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2945 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__5_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2060) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2944 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n764), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n732), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2060), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2057) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2943 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__5_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2695) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2942 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n188), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n156), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2695), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2692) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2941 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__5_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2687) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2940 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n764), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n732), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2687), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2684) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2939 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__4_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2050) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2938 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n189), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n157), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2050), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2047) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2937 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__4_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2042) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2936 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n765), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n733), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2042), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2039) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2935 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__4_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2677) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2934 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n189), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n157), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2677), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2674) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2933 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__4_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2669) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2932 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n765), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n733), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2669), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2666) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2931 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__3_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2032) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2930 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n190), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n158), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2032), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2029) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2929 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__3_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2024) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2928 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n734), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2024), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2021) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2927 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__3_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2659) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2926 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n190), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n158), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2659), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2656) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2925 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__3_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2651) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2924 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n766), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n734), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2651), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2648) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2923 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__2_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2014) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2922 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n191), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n159), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2014), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2011) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2921 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__2_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2006) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2920 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n735), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2006), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2003) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2919 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__2_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2641) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2918 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n191), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n159), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2641), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2638) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2917 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__2_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2633) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2916 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n767), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n735), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2633), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2630) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2915 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__1_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1996) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2914 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n192), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n160), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1996), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1993) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2913 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__1_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1988) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2912 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n736), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1988), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1985) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2911 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__1_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2623) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2910 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n192), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n160), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2623), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2620) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2909 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__1_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2615) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2908 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n768), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n736), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2615), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2612) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2907 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__0_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1966) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2906 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n193), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n161), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1966), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1957) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2905 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__0_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1940) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2904 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n769), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n737), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1940), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1931) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2903 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__0_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2593) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2902 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n193), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n161), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2593), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2584) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2901 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__0_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2567) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2900 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n769), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n737), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2567), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2558) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2899 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2545) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2898 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n34), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2545), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2544) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2897 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2527) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2896 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n610), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n578), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2527), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2526) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2895 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3172) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2894 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n34), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3172), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3171) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2893 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3154) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2892 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n610), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n578), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3154), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3153) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2891 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2517) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2890 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n35), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2517), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2516) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2889 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2509) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2888 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n611), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n579), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2509), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2508) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2887 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3144) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2886 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n35), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3144), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3143) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2885 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3136) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2884 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n611), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n579), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3136), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3135) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2883 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2499) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2882 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n36), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2499), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2498) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2881 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2491) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2880 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n612), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n580), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2491), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2490) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2879 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3126) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2878 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n36), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3126), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3125) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2877 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3118) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2876 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n612), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n580), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3118), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3117) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2875 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2481) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2874 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n37), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n5), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2481), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2480) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2873 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2473) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2872 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n613), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n581), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2473), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2472) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2871 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3108) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2870 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n37), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n5), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3108), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3107) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2869 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3100) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2868 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n613), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n581), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3100), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3099) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2867 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2463) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2866 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n38), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n6), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2463), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2462) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2865 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2455) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2864 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n614), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n582), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2455), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2454) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2863 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3090) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2862 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n38), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n6), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3090), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3089) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2861 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3082) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2860 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n614), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n582), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3082), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3081) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2859 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2445) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2858 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n39), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n7), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2445), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2444) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2857 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2437) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2856 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n615), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n583), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2437), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2436) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2855 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3072) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2854 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n39), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n7), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3072), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3071) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2853 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3064) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2852 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n615), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n583), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3064), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3063) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2851 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2427) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2850 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n40), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n8), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2427), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2426) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2849 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2419) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2848 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n616), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n584), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2419), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2418) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2847 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3054) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2846 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n40), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n8), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3054), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3053) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2845 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3046) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2844 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n616), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n584), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3046), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3045) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2843 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2409) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2842 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n41), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n9), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2409), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2408) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2841 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2401) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2840 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n617), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n585), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2401), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2400) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2839 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3036) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2838 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n41), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n9), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3036), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3035) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2837 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3028) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2836 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n617), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n585), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3028), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3027) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2835 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2391) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2834 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n42), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n10), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2391), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2390) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2833 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2383) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2832 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n618), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n586), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2383), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2382) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2831 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3018) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2830 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n42), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n10), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3018), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3017) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2829 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3010) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2828 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n618), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n586), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3010), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3009) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2827 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2373) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2826 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n43), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n11), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2373), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2372) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2825 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2365) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2824 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n619), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n587), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2365), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2364) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2823 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3000) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2822 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n43), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n11), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3000), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2999) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2821 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2992) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2820 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n619), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n587), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2992), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2991) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2819 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2355) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2818 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n44), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n12), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2355), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2354) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2817 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2347) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2816 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n620), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n588), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2347), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2346) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2815 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2982) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2814 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n44), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n12), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2982), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2981) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2813 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2974) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2812 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n620), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n588), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2974), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2973) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2811 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2337) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2810 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n45), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n13), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2337), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2336) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2809 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2329) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2808 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n621), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n589), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2329), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2328) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2807 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2964) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2806 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n45), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n13), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2964), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2963) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2805 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2956) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2804 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n621), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n589), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2956), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2955) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2803 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2319) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2802 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n46), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n14), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2319), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2318) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2801 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2311) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2800 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n622), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n590), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2311), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2310) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2799 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2946) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2798 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n46), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n14), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2946), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2945) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2797 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2938) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2796 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n622), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n590), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2938), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2937) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2795 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2301) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2794 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n47), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n15), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2301), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2300) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2793 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2293) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2792 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n623), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n591), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2293), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2292) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2791 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2928) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2790 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n47), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n15), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2928), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2927) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2789 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2920) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2788 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n623), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n591), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2920), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2919) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2787 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2283) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2786 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n48), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n16), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2283), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2282) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2785 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2275) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2784 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n624), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n592), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2275), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2274) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2783 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2910) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2782 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n48), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n16), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2910), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2909) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2781 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2902) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2780 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n624), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n592), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2902), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2901) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2779 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2265) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2778 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n49), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n17), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2265), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2264) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2777 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2257) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2776 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n625), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n593), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2257), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2256) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2775 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2892) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2774 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n49), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n17), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2892), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2891) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2773 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2884) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2772 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n625), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n593), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2884), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2883) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2771 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2247) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2770 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n50), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n18), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2247), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2246) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2769 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2239) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2768 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n626), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n594), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2239), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2238) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2767 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2874) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2766 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n50), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n18), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2874), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2873) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2765 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2866) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2764 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n626), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n594), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2866), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2865) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2763 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2229) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2762 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n51), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n19), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2229), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2228) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2761 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2221) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2760 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n627), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n595), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2221), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2220) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2759 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2856) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2758 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n51), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n19), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2856), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2855) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2757 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2848) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2756 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n627), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n595), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2848), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2847) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2755 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2211) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2754 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n52), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n20), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2211), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2210) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2753 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2203) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2752 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n628), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n596), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2203), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2202) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2751 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2838) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2750 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n52), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n20), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2838), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2837) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2749 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2830) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2748 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n628), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n596), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2830), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2829) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2747 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2193) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2746 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n53), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n21), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2193), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2192) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2745 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2185) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2744 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n629), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n597), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2185), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2184) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2743 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2820) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2742 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n53), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n21), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2820), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2819) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2741 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2812) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2740 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n629), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n597), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2812), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2811) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2739 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2175) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2738 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n54), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n22), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2175), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2174) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2737 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2167) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2736 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n630), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n598), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2167), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2166) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2735 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2802) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2734 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n54), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n22), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2802), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2801) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2733 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2794) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2732 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n630), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n598), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2794), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2793) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2731 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2157) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2730 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n55), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n23), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2156) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2729 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2149) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2728 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n631), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n599), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2149), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2148) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2727 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2784) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2726 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n55), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n23), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2784), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2783) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2725 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2776) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2724 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n631), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n599), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2776), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2775) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2723 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2139) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2722 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n56), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n24), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2139), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2138) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2721 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2131) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2720 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n632), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n600), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2131), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2130) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2719 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2766) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2718 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n56), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n24), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2766), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2765) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2717 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2758) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2716 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n632), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n600), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2758), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2757) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2715 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2121) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2714 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n57), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n25), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2121), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2120) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2713 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2113) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2712 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n633), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n601), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2113), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2112) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2711 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2748) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2710 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n57), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n25), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2748), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2747) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2709 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2740) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2708 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n633), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n601), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2740), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2739) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2707 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2103) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2706 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n58), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n26), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2103), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2102) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2705 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2095) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2704 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n634), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n602), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2095), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2094) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2703 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2730) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2702 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n58), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n26), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2730), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2729) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2701 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2722) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2700 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n634), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n602), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2722), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2721) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2699 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2085) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2698 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n59), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n27), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2085), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2084) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2697 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2077) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2696 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n635), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n603), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2077), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2076) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2695 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2712) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2694 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n59), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n27), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2712), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2711) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2693 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2704) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2692 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n635), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n603), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2704), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2703) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2691 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2067) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2690 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n60), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n28), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2067), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2066) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2689 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2059) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2688 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n636), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n604), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2059), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2058) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2687 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2694) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2686 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n60), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n28), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2694), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2693) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2685 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2686) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2684 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n636), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n604), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2686), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2685) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2683 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2049) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2682 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n61), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n29), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2049), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2048) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2681 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2041) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2680 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n637), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n605), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2041), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2040) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2679 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2676) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2678 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n61), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n29), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2676), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2675) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2677 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2668) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2676 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n637), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n605), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2668), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2667) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2675 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2031) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2674 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n62), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n30), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2031), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2030) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2673 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2023) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2672 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n638), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n606), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2023), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2022) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2671 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2658) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2670 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n62), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n30), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2658), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2657) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2669 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2650) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2668 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n638), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n606), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2650), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2649) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2667 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2013) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2666 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n63), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n31), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2013), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2012) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2665 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2005) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2664 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n639), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n607), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2005), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2004) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2663 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2640) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2662 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n63), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n31), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2640), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2639) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2661 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2632) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2660 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n639), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n607), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2632), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2631) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2659 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1995) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2658 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n64), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n32), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1995), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1994) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2657 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1987) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2656 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n640), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n608), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1987), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1986) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2655 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2622) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2654 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n64), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n32), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2622), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2621) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2653 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2614) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2652 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n640), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n608), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2614), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2613) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2651 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1961) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2650 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n65), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n33), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1961), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1958) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2649 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1935) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2648 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n641), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n609), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1935), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1932) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2647 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2588) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2646 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n65), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n33), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2588), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2585) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2645 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2562) );
  OAI221_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2644 ( .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n641), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n609), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747), .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2562), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2559) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2643 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__31_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2553) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2642 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__31_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__31_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3180) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2641 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__30_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2520) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2640 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__30_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__30_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3147) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2639 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__29_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2502) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2638 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__29_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__29_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3129) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2637 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__28_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2484) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2636 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__28_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__28_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3111) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2635 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__27_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2466) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2634 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__27_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__27_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3093) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2633 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__26_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2448) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2632 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__26_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__26_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3075) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2631 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__25_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2430) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2630 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__25_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__25_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3057) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2629 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__24_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2412) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2628 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__24_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__24_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3039) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2627 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__23_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2394) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2626 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__23_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__23_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3021) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2625 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__22_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2376) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2624 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__22_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__22_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3003) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2623 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__21_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2358) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2622 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__21_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__21_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2985) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2621 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__20_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2340) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2620 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__20_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__20_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2967) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2619 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__19_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2322) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2618 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__19_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__19_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2949) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2617 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__18_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2304) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2616 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__18_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__18_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2931) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2615 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__17_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2286) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2614 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__17_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__17_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2913) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2613 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__16_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2268) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2612 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__16_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__16_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2895) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2611 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__15_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2250) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2610 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__15_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__15_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2877) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2609 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__14_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2232) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2608 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__14_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__14_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2859) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2607 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__13_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2214) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2606 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__13_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__13_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2841) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2605 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__12_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2196) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2604 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__12_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__12_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2823) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2603 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__11_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2178) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2602 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__11_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__11_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2805) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2601 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__10_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2160) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2600 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__10_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__10_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2787) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2599 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__9_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2142) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2598 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__9_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__9_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2769) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2597 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__8_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2124) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2596 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__8_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__8_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2751) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2595 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__7_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2106) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2594 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__7_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__7_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2733) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2593 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__6_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2088) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2592 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__6_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__6_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2715) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2591 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__5_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2070) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2590 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__5_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__5_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2697) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2589 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__4_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2052) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2588 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__4_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__4_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2679) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2587 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__3_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2034) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2586 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__3_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__3_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2661) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2585 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__2_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2016) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2584 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__2_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__2_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2643) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2583 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__1_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1998) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2582 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__1_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__1_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2625) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2581 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__0_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1977) );
  AOI222_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2580 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__0_), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__0_), .C1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203), .C2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2604) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2579 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[23]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4225), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1261) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2578 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1261), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1130) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2577 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[22]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4225), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1260) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2576 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1260), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1131) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2575 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[21]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4225), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1259) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2574 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1259), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1132) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2573 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[20]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4225), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1258) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2572 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1258), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1133) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2571 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[19]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4224), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1257) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2570 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1257), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1134) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2569 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[18]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4224), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1256) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2568 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1256), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1135) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2567 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[17]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4224), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1255) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2566 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1255), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1136) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2565 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[16]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4224), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1254) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2564 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1254), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1137) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2563 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[15]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4224), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1253) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2562 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1253), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1138) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2561 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[14]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4223), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1252) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2560 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1252), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1139) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2559 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[13]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4223), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1251) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2558 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1251), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1140) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2557 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219), .A2(
        dp_wr_data_id_i[12]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4223), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1250) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2556 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1250), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1141) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2555 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[11]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4223), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1249) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2554 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1249), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1142) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2553 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[10]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4223), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1248) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2552 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1248), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1143) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2551 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[9]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4222), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1247) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2550 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1247), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1144) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2549 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[8]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4222), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1246) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2548 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1246), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1145) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2547 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[7]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4222), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1245) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2546 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1245), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1146) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2545 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[6]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4222), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1244) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2544 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1244), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1147) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2543 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[5]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4222), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1243) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2542 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1243), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1148) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2541 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[4]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4221), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1242) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2540 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1242), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1149) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2539 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[3]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4221), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1241) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2538 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1241), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1150) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2537 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[2]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4221), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1240) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2536 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1240), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1151) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2535 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[1]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4221), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1239) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2534 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1239), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1152) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2533 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218), .A2(
        dp_wr_data_id_i[0]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4221), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1237) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2532 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1237), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1153) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2531 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220), .A2(dp_n12), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4227), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1269) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2530 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1269), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1122) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2529 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220), .A2(dp_n10), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4227), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1268) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2528 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1268), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1123) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2527 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220), .A2(
        dp_wr_data_id_i[29]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4226), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1267) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2526 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1267), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1124) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2525 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220), .A2(
        dp_wr_data_id_i[28]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4226), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1266) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2524 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1266), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1125) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2523 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220), .A2(dp_n8), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4226), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1265) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2522 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1265), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1126) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2521 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220), .A2(dp_n6), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4226), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1264) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2520 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1264), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1127) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2519 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220), .A2(
        dp_wr_data_id_i[25]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4226), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1263) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2518 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1263), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1128) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2517 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4220), .A2(
        dp_wr_data_id_i[24]), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4225), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1262) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2516 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1262), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1129) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2515 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4020), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1677) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2514 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1677), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n490) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2513 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4020), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1676) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2512 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1676), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n491) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2511 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4020), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1675) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2510 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1675), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n492) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2509 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4020), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1674) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2508 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1674), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n493) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2507 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4019), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1673) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2506 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1673), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n494) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2505 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4019), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1672) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2504 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1672), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n495) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2503 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4019), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1671) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2502 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1671), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n496) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2501 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4019), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1670) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2500 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1670), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n497) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2499 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4019), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1669) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2498 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1669), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n498) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2497 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4018), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1668) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2496 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1668), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n499) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2495 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4018), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1667) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2494 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1667), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n500) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2493 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4018), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1666) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2492 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1666), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n501) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2491 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4018), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1665) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2490 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1665), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n502) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2489 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4018), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1664) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2488 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1664), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n503) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2487 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4017), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1663) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2486 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1663), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n504) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2485 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4017), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1662) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2484 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1662), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n505) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2483 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4017), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1661) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2482 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1661), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n506) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2481 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4017), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1660) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2480 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1660), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n507) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2479 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4017), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1659) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2478 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1659), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n508) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2477 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4016), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1658) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2476 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1658), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n509) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2475 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4016), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1657) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2474 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1657), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n510) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2473 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4016), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1656) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2472 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1656), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n511) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2471 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4016), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1655) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2470 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1655), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n512) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2469 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4016), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1653) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2468 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1653), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n513) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2467 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4022), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1685) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2466 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1685), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n482) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2465 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4022), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1684) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2464 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1684), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n483) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2463 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4021), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1683) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2462 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1683), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n484) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2461 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4021), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1682) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2460 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1682), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n485) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2459 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4021), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1681) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2458 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1681), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n486) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2457 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4021), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1680) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2456 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1680), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n487) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2455 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4021), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1679) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2454 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1679), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n488) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2453 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4020), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1678) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2452 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1678), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n489) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2451 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4151), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1374) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2450 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1374), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n906) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2449 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4151), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1373) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2448 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1373), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n907) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2447 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4151), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1372) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2446 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1372), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n908) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2445 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4151), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1371) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2444 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1371), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n909) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2443 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4150), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1370) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2442 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1370), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n910) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2441 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4150), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1369) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2440 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1369), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n911) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2439 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4150), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1368) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2438 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1368), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n912) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2437 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4150), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1367) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2436 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1367), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n913) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2435 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4150), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1366) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2434 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1366), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n914) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2433 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4149), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1365) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2432 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1365), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n915) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2431 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4149), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1364) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2430 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1364), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n916) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2429 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4149), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1363) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2428 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1363), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n917) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2427 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4149), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1362) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2426 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1362), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n918) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2425 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4149), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1361) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2424 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1361), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n919) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2423 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4148), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1360) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2422 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1360), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n920) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2421 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4148), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1359) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2420 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1359), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n921) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2419 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4148), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1358) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2418 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1358), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n922) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2417 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4148), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1357) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2416 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1357), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n923) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2415 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4148), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1356) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2414 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1356), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n924) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2413 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4147), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1355) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2412 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1355), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n925) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2411 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4147), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1354) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2410 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1354), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n926) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2409 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4147), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1353) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2408 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1353), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n927) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2407 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4147), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1352) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2406 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1352), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n928) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2405 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4147), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1350) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2404 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1350), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n929) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2403 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3989), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1713) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2402 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1713), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n394) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2401 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3989), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1712) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2400 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1712), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n395) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2399 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3989), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1711) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2398 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1711), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n396) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2397 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3989), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1710) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2396 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1710), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n397) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2395 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3988), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1709) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2394 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1709), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n398) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2393 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3988), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1708) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2392 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1708), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n399) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2391 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3988), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1707) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2390 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1707), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n400) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2389 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3988), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1706) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2388 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1706), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n401) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2387 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3988), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1705) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2386 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1705), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n402) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2385 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3987), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1704) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2384 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1704), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n403) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2383 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3987), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1703) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2382 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1703), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n404) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2381 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3987), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1702) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2380 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1702), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n405) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2379 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3987), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1701) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2378 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1701), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n406) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2377 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3987), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1700) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2376 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1700), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n407) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2375 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3986), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1699) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2374 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1699), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n408) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2373 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3986), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1698) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2372 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1698), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n409) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2371 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3986), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1697) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2370 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1697), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n410) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2369 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3986), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1696) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2368 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1696), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n411) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2367 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3986), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1695) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2366 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1695), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n412) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2365 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3985), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1694) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2364 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1694), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n413) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2363 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3985), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1693) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2362 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1693), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n414) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2361 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3985), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1692) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2360 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1692), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n415) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2359 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3985), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1691) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2358 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1691), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n416) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2357 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3985), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1689) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2356 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1689), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n417) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2355 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4153), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1382) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2354 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1382), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n898) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2353 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4153), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1381) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2352 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1381), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n899) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2351 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4152), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1380) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2350 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1380), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n900) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2349 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4152), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1379) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2348 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1379), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n901) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2347 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4152), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1378) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2346 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1378), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n902) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2345 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4152), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1377) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2344 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1377), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n903) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2343 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4152), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1376) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2342 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1376), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n904) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2341 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4151), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1375) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2340 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1375), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n905) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2339 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3991), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1721) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2338 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1721), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n386) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2337 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3991), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1720) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2336 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1720), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n387) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2335 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3990), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1719) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2334 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1719), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n388) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2333 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3990), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1718) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2332 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1718), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n389) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2331 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3990), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1717) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2330 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1717), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n390) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2329 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3990), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1716) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2328 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1716), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n391) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2327 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3990), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1715) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2326 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1715), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n392) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2325 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3989), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1714) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2324 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1714), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n393) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2323 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3929), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1848) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2322 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1848), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n202) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2321 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3929), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1847) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2320 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1847), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n203) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2319 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3929), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1846) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2318 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1846), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n204) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2317 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3929), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1845) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2316 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1845), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n205) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2315 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3928), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1844) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2314 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1844), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n206) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2313 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3928), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1843) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2312 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1843), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n207) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2311 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3928), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1842) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2310 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1842), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n208) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2309 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3928), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1841) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2308 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1841), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n209) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2307 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3928), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1840) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2306 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1840), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n210) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2305 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3927), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1839) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2304 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1839), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n211) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2303 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3927), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1838) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2302 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1838), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n212) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2301 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3927), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1837) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2300 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1837), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n213) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2299 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3927), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1836) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2298 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1836), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n214) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2297 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3927), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1835) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2296 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1835), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n215) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2295 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3926), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1834) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2294 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1834), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n216) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2293 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3926), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1833) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2292 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1833), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n217) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2291 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3926), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1832) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2290 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1832), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n218) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2289 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3926), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1831) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2288 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1831), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n219) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2287 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3926), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1830) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2286 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1830), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n220) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2285 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3925), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1829) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2284 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1829), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n221) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2283 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3925), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1828) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2282 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1828), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n222) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2281 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3925), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1827) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2280 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1827), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n223) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2279 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3925), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1826) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2278 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1826), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n224) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2277 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3925), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1824) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2276 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1824), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n225) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2275 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3938), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1814) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2274 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1814), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n234) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2273 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3938), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1813) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2272 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1813), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n235) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2271 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3938), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1812) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2270 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1812), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n236) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2269 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3938), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1811) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2268 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1811), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n237) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2267 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3937), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1810) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2266 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1810), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n238) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2265 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3937), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1809) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2264 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1809), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n239) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2263 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3937), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1808) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2262 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1808), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n240) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2261 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3937), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1807) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2260 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1807), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n241) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2259 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3937), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1806) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2258 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1806), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n242) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2257 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3936), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1805) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2256 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1805), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n243) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2255 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3936), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1804) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2254 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1804), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n244) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2253 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3936), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1803) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2252 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1803), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n245) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2251 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3936), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1802) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2250 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1802), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n246) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2249 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3936), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1801) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2248 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1801), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n247) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2247 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3935), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1800) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2246 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1800), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n248) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2245 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3935), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1799) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2244 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1799), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n249) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2243 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3935), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1798) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2242 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1798), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n250) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2241 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3935), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1797) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2240 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1797), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n251) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2239 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3935), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1796) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2238 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1796), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n252) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2237 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3934), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1795) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2236 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1795), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n253) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2235 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3934), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1794) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2234 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1794), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n254) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2233 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3934), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1793) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2232 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1793), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n255) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2231 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3934), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1792) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2230 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1792), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n256) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2229 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3934), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1790) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2228 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1790), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n257) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2227 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4071), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1576) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2226 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1576), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n650) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2225 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4071), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1575) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2224 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1575), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n651) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2223 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4071), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1574) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2222 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1574), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n652) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2221 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4071), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1573) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2220 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1573), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n653) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2219 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4070), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1572) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2218 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1572), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n654) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2217 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4070), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1571) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2216 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1571), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n655) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2215 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4070), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1570) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2214 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1570), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n656) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2213 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4070), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1569) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2212 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1569), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n657) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2211 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4070), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1568) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2210 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1568), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n658) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2209 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4069), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1567) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2208 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1567), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n659) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2207 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4069), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1566) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2206 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1566), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n660) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2205 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4069), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1565) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2204 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1565), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n661) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2203 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4069), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1564) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2202 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1564), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n662) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2201 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4069), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1563) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2200 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1563), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n663) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2199 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4068), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1562) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2198 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1562), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n664) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2197 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4068), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1561) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2196 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1561), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n665) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2195 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4068), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1560) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2194 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1560), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n666) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2193 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4068), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1559) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2192 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1559), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n667) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2191 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4068), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1558) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2190 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1558), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n668) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2189 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4067), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1557) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2188 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1557), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n669) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2187 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4067), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1556) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2186 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1556), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n670) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2185 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4067), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1555) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2184 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1555), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n671) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2183 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4067), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1554) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2182 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1554), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n672) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2181 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4067), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1552) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2180 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1552), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n673) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2179 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4080), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1543) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2178 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1543), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n682) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2177 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4080), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1542) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2176 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1542), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n683) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2175 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4080), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1541) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2174 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1541), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n684) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2173 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4080), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1540) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2172 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1540), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n685) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2171 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4079), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1539) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2170 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1539), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n686) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2169 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4079), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1538) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2168 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1538), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n687) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2167 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4079), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1537) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2166 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1537), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n688) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2165 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4079), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1536) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2164 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1536), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n689) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2163 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4079), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1535) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2162 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1535), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n690) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2161 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4078), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1534) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2160 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1534), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n691) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2159 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4078), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1533) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2158 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n692) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2157 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4078), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1532) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2156 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n693) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2155 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4078), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1531) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2154 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1531), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n694) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2153 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4078), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1530) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2152 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n695) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2151 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4077), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1529) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2150 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n696) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2149 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4077), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1528) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2148 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1528), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n697) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2147 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4077), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1527) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2146 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1527), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n698) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2145 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4077), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1526) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2144 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1526), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n699) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2143 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4077), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1525) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2142 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1525), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n700) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2141 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4076), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1524) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2140 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1524), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n701) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2139 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4076), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1523) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2138 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1523), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n702) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2137 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4076), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1522) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2136 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1522), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n703) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2135 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4076), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1521) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2134 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1521), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n704) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2133 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4076), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1519) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2132 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1519), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n705) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2131 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3931), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1856) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2130 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1856), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n194) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2129 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3931), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1855) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2128 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1855), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n195) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2127 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3930), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1854) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2126 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1854), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n196) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2125 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3930), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1853) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2124 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1853), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n197) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2123 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3930), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1852) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2122 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1852), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n198) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2121 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3930), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1851) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2120 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1851), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n199) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2119 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3930), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1850) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2118 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1850), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n200) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2117 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3929), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1849) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2116 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1849), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n201) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2115 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3940), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1822) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2114 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1822), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n226) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2113 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3940), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1821) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2112 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1821), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n227) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2111 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3939), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1820) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2110 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1820), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n228) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2109 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3939), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1819) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2108 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1819), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n229) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2107 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3939), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1818) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2106 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1818), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n230) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2105 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3939), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1817) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2104 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1817), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n231) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2103 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3939), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1816) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2102 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1816), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n232) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2101 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3938), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1815) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2100 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1815), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n233) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2099 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4073), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1584) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2098 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1584), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n642) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2097 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4073), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1583) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2096 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1583), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n643) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2095 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4072), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1582) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2094 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1582), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n644) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2093 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4072), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1581) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2092 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1581), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n645) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2091 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4072), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1580) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2090 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1580), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n646) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2089 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4072), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1579) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2088 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1579), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n647) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2087 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4072), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1578) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2086 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1578), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n648) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2085 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4071), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1577) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2084 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1577), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n649) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2083 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4082), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1551) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2082 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1551), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n674) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2081 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4082), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1550) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2080 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1550), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n675) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2079 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4081), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1549) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2078 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1549), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n676) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2077 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4081), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1548) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2076 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1548), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n677) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2075 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4081), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1547) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2074 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1547), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n678) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2073 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4081), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1546) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2072 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1546), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n679) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2071 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4081), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1545) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2070 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1545), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n680) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2069 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4080), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1544) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2068 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1544), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n681) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2067 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3948), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1781) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2066 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1781), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n266) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2065 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3948), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1780) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2064 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1780), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n267) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2063 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3948), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1779) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2062 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1779), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n268) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2061 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3948), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1778) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2060 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1778), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n269) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2059 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3947), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1777) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2058 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1777), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n270) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2057 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3947), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1776) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2056 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1776), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n271) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2055 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3947), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1775) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2054 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1775), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n272) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2053 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3947), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1774) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2052 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1774), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n273) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2051 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3947), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1773) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2050 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1773), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n274) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2049 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3946), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1772) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2048 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1772), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n275) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2047 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3946), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1771) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2046 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1771), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n276) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2045 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3946), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1770) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2044 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1770), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n277) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2043 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3946), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1769) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2042 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1769), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n278) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2041 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3946), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1768) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2040 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1768), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n279) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2039 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3945), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1767) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2038 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1767), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n280) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2037 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3945), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1766) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2036 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1766), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n281) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2035 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3945), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1765) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2034 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1765), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n282) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2033 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3945), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1764) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2032 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1764), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n283) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2031 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3945), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1763) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2030 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1763), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n284) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2029 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3944), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1762) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2028 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1762), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n285) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2027 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3944), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1761) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2026 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1761), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n286) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2025 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3944), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1760) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2024 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1760), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n287) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2023 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3944), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1759) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2022 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1759), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n288) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2021 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3944), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1757) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2020 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1757), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n289) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2019 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4030), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1644) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2018 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1644), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n522) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2017 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4030), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1643) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2016 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1643), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n523) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2015 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4030), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1642) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2014 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1642), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n524) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2013 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4030), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1641) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2012 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1641), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n525) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2011 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4029), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1640) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2010 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1640), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n526) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2009 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4029), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1639) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2008 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1639), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n527) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2007 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4029), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1638) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2006 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1638), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n528) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2005 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4029), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1637) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2004 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1637), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n529) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2003 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4029), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1636) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2002 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1636), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n530) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2001 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4028), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1635) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2000 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1635), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n531) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1999 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4028), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1634) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1998 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1634), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n532) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1997 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4028), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1633) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1996 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1633), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n533) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1995 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4028), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1632) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1994 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1632), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n534) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1993 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4028), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1631) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1992 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1631), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n535) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1991 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4027), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1630) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1990 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1630), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n536) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1989 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4027), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1629) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1988 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1629), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n537) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1987 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4027), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1628) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1986 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1628), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n538) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1985 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4027), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1627) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1984 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1627), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n539) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1983 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4027), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1626) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1982 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1626), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n540) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1981 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4026), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1625) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1980 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1625), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n541) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1979 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4026), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1624) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1978 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1624), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n542) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1977 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4026), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1623) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1976 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1623), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n543) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1975 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4026), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1622) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1974 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1622), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n544) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1973 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4026), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1620) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1972 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1620), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n545) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1971 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4112), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1507) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1970 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1507), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n778) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1969 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4112), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1506) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1968 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1506), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n779) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1967 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4112), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1505) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1966 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1505), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n780) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1965 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4112), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1504) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1964 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1504), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n781) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1963 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4111), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1503) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1962 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1503), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n782) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1961 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4111), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1502) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1960 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1502), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n783) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1959 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4111), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1501) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1958 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1501), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n784) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1957 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4111), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1500) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1956 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1500), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n785) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1955 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4111), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1499) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1954 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1499), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n786) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1953 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4110), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1498) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1952 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1498), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n787) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1951 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4110), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1497) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1950 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1497), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n788) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1949 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4110), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1496) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1948 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1496), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n789) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1947 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4110), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1495) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1946 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1495), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n790) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1945 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4110), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1494) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1944 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1494), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n791) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1943 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4109), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1493) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1942 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1493), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n792) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1941 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4109), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1492) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1940 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1492), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n793) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1939 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4109), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1491) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1938 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1491), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n794) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1937 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4109), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1490) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1936 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1490), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n795) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1935 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4109), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1489) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1934 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1489), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n796) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1933 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4108), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1488) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1932 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1488), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n797) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1931 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4108), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1487) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1930 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1487), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n798) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1929 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4108), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1486) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1928 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1486), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n799) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1927 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4108), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1485) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1926 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1485), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n800) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1925 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4108), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1483) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1924 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1483), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n801) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1923 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3888), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1916) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1922 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1916), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n74) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1921 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3888), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1915) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1920 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1915), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n75) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1919 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3888), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1914) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1918 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1914), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n76) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1917 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3888), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1913) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1916 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1913), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n77) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1915 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3887), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1912) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1914 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1912), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n78) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1913 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3887), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1911) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1912 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1911), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n79) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1911 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3887), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1910) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1910 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1910), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n80) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1909 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3887), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1909) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1908 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1909), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n81) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1907 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3887), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1908) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1906 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1908), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n82) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1905 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3886), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1907) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1904 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1907), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n83) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1903 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3886), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1906) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1902 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1906), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n84) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1901 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3886), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1905) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1900 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1905), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n85) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1899 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3886), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1904) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1898 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1904), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n86) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1897 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3886), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1903) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1896 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1903), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n87) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1895 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3885), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1902) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1894 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1902), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n88) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1893 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3885), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1901) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1892 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1901), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n89) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1891 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3885), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1900) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1890 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1900), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n90) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1889 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3885), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1899) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1888 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1899), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n91) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1887 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3885), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1898) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1886 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1898), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n92) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1885 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3884), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1897) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1884 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1897), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n93) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1883 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3884), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1896) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1882 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1896), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n94) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1881 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3884), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1895) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1880 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1895), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n95) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1879 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3884), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1894) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1878 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1894), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n96) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1877 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3884), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1892) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1876 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1892), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n97) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1875 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3898), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1883) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1874 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1883), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n106) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1873 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3898), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1882) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1872 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1882), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n107) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1871 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3898), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1881) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1870 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1881), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n108) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1869 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3898), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1880) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1868 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1880), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n109) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1867 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3897), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1879) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1866 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1879), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n110) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1865 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3897), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1878) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1864 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1878), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n111) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1863 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3897), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1877) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1862 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1877), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n112) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1861 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3897), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1876) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1860 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1876), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n113) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1859 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3897), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1875) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1858 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1875), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n114) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1857 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3896), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1874) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1856 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1874), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n115) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1855 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3896), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1873) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1854 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1873), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n116) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1853 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3896), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1872) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1852 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1872), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n117) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1851 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3896), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1871) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1850 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1871), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n118) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1849 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3896), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1870) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1848 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1870), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n119) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1847 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3895), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1869) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1846 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1869), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n120) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1845 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3895), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1868) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1844 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1868), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n121) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1843 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3895), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1867) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1842 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1867), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n122) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1841 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3895), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1866) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1840 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1866), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n123) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1839 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3895), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1865) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1838 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1865), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n124) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1837 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3894), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1864) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1836 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1864), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n125) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1835 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3894), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1863) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1834 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1863), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n126) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1833 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3894), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1862) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1832 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1862), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n127) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1831 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3894), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1861) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1830 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1861), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n128) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1829 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3894), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1859) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1828 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1859), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n129) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1827 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3980), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1746) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1826 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1746), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n362) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1825 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3980), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1745) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1824 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1745), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n363) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1823 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3980), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1744) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1822 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1744), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n364) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1821 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3980), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1743) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1820 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1743), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n365) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1819 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3979), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1742) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1818 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1742), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n366) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1817 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3979), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1741) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1816 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1741), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n367) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1815 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3979), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1740) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1814 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1740), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n368) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1813 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3979), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1739) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1812 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1739), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n369) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1811 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3979), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1738) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1810 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1738), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n370) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1809 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3978), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1737) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1808 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1737), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n371) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1807 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3978), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1736) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1806 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1736), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n372) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1805 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3978), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1735) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1804 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1735), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n373) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1803 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3978), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1734) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1802 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1734), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n374) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1801 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3978), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1733) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1800 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1733), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n375) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1799 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3977), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1732) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1798 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1732), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n376) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1797 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3977), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1731) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1796 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1731), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n377) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1795 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3977), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1730) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1794 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1730), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n378) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1793 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3977), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1729) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1792 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1729), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n379) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1791 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3977), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1728) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1790 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1728), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n380) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1789 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3976), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1727) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1788 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1727), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n381) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1787 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3976), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1726) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1786 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1726), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n382) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1785 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3976), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1725) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1784 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1725), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n383) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1783 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3976), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1724) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1782 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1724), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n384) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1781 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3976), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1722) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1780 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1722), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n385) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1779 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4132), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1441) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1778 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1441), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n842) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1777 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4132), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1440) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1776 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1440), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n843) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1775 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4132), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1439) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1774 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1439), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n844) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1773 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4132), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1438) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1772 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1438), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n845) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1771 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4131), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1437) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1770 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1437), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n846) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1769 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4131), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1436) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1768 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1436), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n847) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1767 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4131), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1435) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1766 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1435), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n848) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1765 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4131), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1434) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1764 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1434), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n849) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1763 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4131), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1433) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1762 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1433), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n850) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1761 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4130), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1432) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1760 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1432), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n851) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1759 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4130), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1431) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1758 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1431), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n852) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1757 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4130), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1430) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1756 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1430), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n853) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1755 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4130), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1429) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1754 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1429), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n854) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1753 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4130), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1428) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1752 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1428), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n855) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1751 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4129), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1427) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1750 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1427), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n856) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1749 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4129), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1426) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1748 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1426), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n857) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1747 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4129), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1425) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1746 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1425), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n858) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1745 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4129), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1424) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1744 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1424), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n859) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1743 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4129), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1423) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1742 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1423), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n860) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1741 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4128), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1422) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1740 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1422), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n861) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1739 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4128), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1421) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1738 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1421), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n862) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1737 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4128), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1420) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1736 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1420), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n863) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1735 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4128), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1419) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1734 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1419), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n864) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1733 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4128), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1417) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1732 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1417), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n865) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1731 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4142), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1408) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1730 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1408), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n874) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1729 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4142), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1407) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1728 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1407), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n875) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1727 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4142), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1406) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1726 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1406), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n876) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1725 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4142), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1405) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1724 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1405), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n877) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1723 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4141), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1404) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1722 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1404), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n878) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1721 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4141), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1403) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1720 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1403), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n879) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1719 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4141), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1402) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1718 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1402), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n880) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1717 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4141), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1401) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1716 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1401), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n881) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1715 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4141), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1400) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1714 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1400), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n882) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1713 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4140), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1399) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1712 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1399), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n883) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1711 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4140), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1398) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1710 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1398), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n884) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1709 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4140), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1397) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1708 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1397), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n885) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1707 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4140), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1396) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1706 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1396), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n886) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1705 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4140), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1395) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1704 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1395), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n887) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1703 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4139), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1394) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1702 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1394), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n888) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1701 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4139), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1393) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1700 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1393), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n889) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1699 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4139), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1392) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1698 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1392), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n890) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1697 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4139), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1391) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1696 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1391), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n891) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1695 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4139), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1390) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1694 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1390), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n892) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1693 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4138), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1389) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1692 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1389), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n893) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1691 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4138), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1388) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1690 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1388), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n894) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1689 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4138), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1387) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1688 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1387), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n895) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1687 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4138), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1386) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1686 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1386), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n896) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1685 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4138), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1384) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1684 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1384), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n897) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1683 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4040), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1611) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1682 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1611), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n554) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1681 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4040), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1610) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1680 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1610), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n555) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1679 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4040), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1609) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1678 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1609), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n556) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1677 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4040), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1608) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1676 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1608), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n557) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1675 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4039), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1607) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1674 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1607), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n558) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1673 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4039), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1606) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1672 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1606), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n559) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1671 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4039), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1605) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1670 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1605), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n560) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1669 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4039), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1604) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1668 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1604), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n561) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1667 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4039), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1603) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1666 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1603), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n562) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1665 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4038), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1602) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1664 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1602), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n563) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1663 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4038), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1601) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1662 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1601), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n564) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1661 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4038), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1600) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1660 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1600), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n565) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1659 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4038), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1599) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1658 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1599), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n566) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1657 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4038), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1598) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1656 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1598), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n567) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1655 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4037), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1597) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1654 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1597), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n568) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1653 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4037), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1596) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1652 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1596), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n569) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1651 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4037), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1595) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1650 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1595), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n570) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1649 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4037), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1594) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1648 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1594), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n571) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1647 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4037), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1593) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1646 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1593), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n572) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1645 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4036), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1592) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1644 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1592), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n573) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1643 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4036), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1591) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1642 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1591), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n574) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1641 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4036), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1590) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1640 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1590), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n575) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1639 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4036), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1589) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1638 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1589), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n576) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1637 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4036), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1587) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1636 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1587), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n577) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1635 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4122), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1474) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1634 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1474), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n810) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1633 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4122), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1473) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1632 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1473), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n811) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1631 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4122), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1472) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1630 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1472), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n812) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1629 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4122), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1471) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1628 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1471), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n813) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1627 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4121), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1470) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1626 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1470), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n814) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1625 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4121), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1469) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1624 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1469), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n815) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1623 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4121), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1468) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1622 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1468), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n816) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1621 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4121), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1467) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1620 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1467), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n817) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1619 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4121), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1466) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1618 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1466), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n818) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1617 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4120), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1465) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1616 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1465), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n819) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1615 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4120), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1464) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1614 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1464), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n820) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1613 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4120), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1463) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1612 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1463), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n821) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1611 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4120), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1462) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1610 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1462), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n822) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1609 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4120), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1461) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1608 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1461), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n823) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1607 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4119), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1460) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1606 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1460), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n824) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1605 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4119), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1459) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1604 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1459), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n825) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1603 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4119), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1458) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1602 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1458), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n826) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1601 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4119), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1457) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1600 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1457), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n827) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1599 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4119), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1456) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1598 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1456), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n828) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1597 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4118), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1455) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1596 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1455), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n829) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1595 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4118), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1454) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1594 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1454), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n830) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1593 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4118), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1453) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1592 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1453), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n831) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1591 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4118), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1452) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1590 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1452), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n832) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1589 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4118), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1450) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1588 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1450), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n833) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1587 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4215), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1296) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1586 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1296), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1098) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1585 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4215), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1295) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1584 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1295), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1099) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1583 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4215), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1294) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1582 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1294), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1100) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1581 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4215), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1293) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1580 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1293), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1101) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1579 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4214), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1292) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1578 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1292), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1102) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1577 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4214), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1291) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1576 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1291), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1103) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1575 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4214), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1290) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1574 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1290), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1104) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1573 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4214), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1289) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1572 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1289), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1105) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1571 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4214), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1288) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1570 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1288), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1106) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1569 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4213), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1287) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1568 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1287), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1107) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1567 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4213), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1286) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1566 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1286), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1108) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1565 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4213), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1285) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1564 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1285), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1109) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1563 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4213), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1284) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1562 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1284), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1110) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1561 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4213), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1283) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1560 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1283), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1111) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1559 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4212), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1282) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1558 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1282), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1112) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1557 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4212), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1281) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1556 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1281), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1113) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1555 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4212), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1280) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1554 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1280), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1114) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1553 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4212), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1279) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1552 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1279), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1115) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1551 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4212), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1278) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1550 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1278), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1116) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1549 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4211), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1277) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1548 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1277), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1117) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1547 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4211), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1276) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1546 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1276), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1118) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1545 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4211), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1275) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1544 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1275), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1119) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1543 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4211), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1274) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1542 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1274), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1120) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1541 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4211), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1272) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1540 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1272), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1121) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1539 ( .A1(
        dp_wr_data_id_i[23]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4205), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__23_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1330) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1538 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1330), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1066) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1537 ( .A1(
        dp_wr_data_id_i[22]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4205), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__22_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1329) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1536 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1329), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1067) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1535 ( .A1(
        dp_wr_data_id_i[21]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4205), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__21_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1328) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1534 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1328), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1068) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1533 ( .A1(
        dp_wr_data_id_i[20]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4205), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__20_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1327) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1532 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1327), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1069) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1531 ( .A1(
        dp_wr_data_id_i[19]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4204), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__19_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1326) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1530 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1326), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1070) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1529 ( .A1(
        dp_wr_data_id_i[18]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4204), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__18_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1325) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1528 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1325), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1071) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1527 ( .A1(
        dp_wr_data_id_i[17]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4204), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__17_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1324) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1526 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1324), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1072) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1525 ( .A1(
        dp_wr_data_id_i[16]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4204), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__16_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1323) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1524 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1323), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1073) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1523 ( .A1(
        dp_wr_data_id_i[15]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4204), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__15_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1322) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1522 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1322), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1074) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1521 ( .A1(
        dp_wr_data_id_i[14]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4203), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__14_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1321) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1520 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1321), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1075) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1519 ( .A1(
        dp_wr_data_id_i[13]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4203), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__13_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1320) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1518 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1320), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1076) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1517 ( .A1(
        dp_wr_data_id_i[12]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4203), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__12_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1319) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1516 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1319), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1077) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1515 ( .A1(
        dp_wr_data_id_i[11]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4203), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__11_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1318) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1514 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1318), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1078) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1513 ( .A1(
        dp_wr_data_id_i[10]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4203), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__10_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1317) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1512 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1317), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1079) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1511 ( .A1(
        dp_wr_data_id_i[9]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4202), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__9_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1316) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1510 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1316), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1080) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1509 ( .A1(
        dp_wr_data_id_i[8]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4202), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__8_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1315) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1508 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1315), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1081) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1507 ( .A1(
        dp_wr_data_id_i[7]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4202), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__7_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1314) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1506 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1314), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1082) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1505 ( .A1(
        dp_wr_data_id_i[6]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4202), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__6_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1313) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1504 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1313), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1083) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1503 ( .A1(
        dp_wr_data_id_i[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4202), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__5_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1312) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1502 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1312), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1084) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1501 ( .A1(
        dp_wr_data_id_i[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4201), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__4_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1311) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1500 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1311), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1085) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1499 ( .A1(
        dp_wr_data_id_i[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4201), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__3_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1310) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1498 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1310), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1086) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1497 ( .A1(
        dp_wr_data_id_i[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4201), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__2_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1309) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1496 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1309), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1087) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1495 ( .A1(
        dp_wr_data_id_i[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4201), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__1_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1308) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1494 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1308), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1088) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1493 ( .A1(
        dp_wr_data_id_i[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4201), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__0_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1306) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1492 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1306), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1089) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1491 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3950), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1789) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1490 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1789), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n258) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1489 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3950), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1788) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1488 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1788), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n259) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1487 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3949), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1787) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1486 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1787), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n260) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1485 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3949), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1786) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1484 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1786), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n261) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1483 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3949), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1785) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1482 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1785), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n262) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1481 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3949), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1784) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1480 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1784), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n263) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1479 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3949), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1783) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1478 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1783), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n264) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1477 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3943), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3948), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1782) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1476 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1782), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n265) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1475 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4032), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1652) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1474 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1652), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n514) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1473 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4032), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1651) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1472 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1651), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n515) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1471 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4031), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1650) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1470 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1650), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n516) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1469 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4031), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1649) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1468 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1649), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n517) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1467 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4031), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1648) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1466 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1648), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n518) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1465 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4031), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1647) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1464 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1647), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n519) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1463 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4031), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1646) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1462 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1646), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n520) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1461 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4025), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4030), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1645) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1460 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1645), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n521) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1459 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4114), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1515) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1458 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1515), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n770) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1457 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4114), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1514) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1456 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1514), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n771) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1455 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4113), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1513) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1454 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1513), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n772) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1453 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4113), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1512) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1452 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1512), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n773) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1451 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4113), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1511) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1450 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1511), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n774) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1449 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4113), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1510) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1448 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1510), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n775) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1447 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4113), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1509) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1446 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1509), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n776) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1445 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4107), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4112), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1508) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1444 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1508), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n777) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1443 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3890), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1924) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1442 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1924), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n66) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1441 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3890), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1923) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1440 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1923), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n67) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1439 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3889), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1922) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1438 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1922), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n68) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1437 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3889), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1921) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1436 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1921), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n69) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1435 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3889), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1920) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1434 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1920), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n70) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1433 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3889), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1919) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1432 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1919), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n71) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1431 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3889), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1918) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1430 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1918), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n72) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1429 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3883), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3888), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1917) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1428 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1917), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n73) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1427 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3900), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1891) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1426 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1891), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n98) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1425 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3900), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1890) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1424 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1890), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n99) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1423 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3899), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1889) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1422 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1889), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n100) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1421 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3899), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1888) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1420 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1888), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n101) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1419 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3899), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1887) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1418 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1887), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n102) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1417 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3899), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1886) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1416 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1886), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n103) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1415 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3899), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1885) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1414 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1885), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n104) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1413 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3893), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3898), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1884) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1412 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1884), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n105) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1411 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3982), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1754) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1410 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1754), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n354) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1409 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3982), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1753) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1408 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1753), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n355) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1407 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3981), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1752) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1406 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1752), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n356) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1405 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3981), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1751) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1404 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1751), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n357) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1403 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3981), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1750) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1402 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1750), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n358) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1401 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3981), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1749) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1400 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1749), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n359) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1399 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3981), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1748) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1398 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1748), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n360) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1397 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3975), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3980), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1747) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1396 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1747), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n361) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1395 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4134), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1449) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1394 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1449), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n834) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1393 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4134), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1448) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1392 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1448), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n835) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1391 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4133), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1447) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1390 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1447), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n836) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1389 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4133), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1446) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1388 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1446), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n837) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1387 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4133), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1445) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1386 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1445), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n838) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1385 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4133), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1444) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1384 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1444), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n839) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1383 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4133), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1443) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1382 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1443), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n840) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1381 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4127), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4132), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1442) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1380 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1442), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n841) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1379 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4144), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1416) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1378 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1416), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n866) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1377 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4144), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1415) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1376 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1415), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n867) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1375 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4143), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1414) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1374 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1414), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n868) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1373 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4143), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1413) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1372 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1413), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n869) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1371 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4143), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1412) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1370 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1412), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n870) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1369 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4143), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1411) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1368 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1411), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n871) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1367 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4143), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1410) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1366 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1410), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n872) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1365 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4137), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4142), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1409) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1364 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1409), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n873) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1363 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4042), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1619) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1362 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1619), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n546) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1361 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4042), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1618) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1360 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1618), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n547) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1359 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4041), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1617) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1358 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1617), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n548) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1357 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4041), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1616) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1356 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1616), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n549) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1355 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4041), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1615) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1354 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1615), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n550) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1353 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4041), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1614) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1352 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1614), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n551) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1351 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4041), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1613) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1350 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1613), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n552) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1349 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4035), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4040), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1612) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1348 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1612), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n553) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1347 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4124), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1482) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1346 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1482), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n802) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1345 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4124), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1481) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1344 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1481), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n803) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1343 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4123), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1480) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1342 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1480), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n804) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1341 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4123), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1479) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1340 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1479), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n805) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1339 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4123), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1478) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1338 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1478), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n806) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1337 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4123), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1477) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1336 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1477), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n807) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1335 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4123), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1476) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1334 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1476), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n808) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1333 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4117), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4122), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1475) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1332 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1475), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n809) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1331 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4217), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1304) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1330 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1304), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1090) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1329 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4217), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1303) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1328 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1303), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1091) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1327 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4216), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1302) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1326 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1302), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1092) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1325 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4216), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1301) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1324 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1301), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1093) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1323 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4216), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1300) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1322 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1300), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1094) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1321 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4216), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1299) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1320 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1299), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1095) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1319 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4216), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1298) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1318 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1298), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1096) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1317 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4210), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4215), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1297) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1316 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1297), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1097) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1315 ( .A1(dp_n12), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__31_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1338) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1314 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1338), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1058) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1313 ( .A1(dp_n10), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4207), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__30_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1337) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1312 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1337), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1059) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1311 ( .A1(
        dp_wr_data_id_i[29]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__29_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1336) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1310 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1336), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1060) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1309 ( .A1(
        dp_wr_data_id_i[28]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__28_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1335) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1308 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1335), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1061) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1307 ( .A1(dp_n8), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__27_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1334) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1306 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1334), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1062) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1305 ( .A1(dp_n6), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__26_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1333) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1304 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1333), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1063) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1303 ( .A1(
        dp_wr_data_id_i[25]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4206), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__25_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1332) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1302 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1332), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1064) );
  AOI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1301 ( .A1(
        dp_wr_data_id_i[24]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4200), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4205), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__24_), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1331) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1300 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1331), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1065) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1299 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4178), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n994), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3244) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1298 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4178), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n995), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3243) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1297 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4178), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n996), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3242) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1296 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4178), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n997), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3241) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1295 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4179), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n998), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3240) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1294 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4179), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n999), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3239) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1293 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4179), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1000), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3238) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1292 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4179), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1001), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3237) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1291 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4180), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1002), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3236) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1290 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4180), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1003), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3235) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1289 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4180), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1004), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3234) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1288 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4180), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1005), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3233) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1287 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4181), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1006), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3232) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1286 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4181), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1007), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3231) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1285 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4181), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1008), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3230) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1284 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4181), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1009), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3229) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1283 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4182), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1010), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3228) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1282 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4182), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1011), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3227) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1281 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4182), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1012), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3226) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1280 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4182), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1013), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3225) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1279 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4183), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1014), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3224) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1278 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4183), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1015), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3223) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1277 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4183), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1016), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3222) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1276 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4183), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1017), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3221) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1275 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4184), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1018), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3220) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1274 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4184), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1019), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3219) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1273 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4184), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1020), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3218) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1272 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4184), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1021), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3217) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1271 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4185), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1022), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3216) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1270 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4185), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1023), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3215) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1269 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4185), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1024), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3214) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1268 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4185), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1025), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3213) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1267 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4173), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n986), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3252) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1266 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4173), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n987), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3251) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1265 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4173), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n988), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3250) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1264 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4173), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n989), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3249) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1263 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4174), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n990), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3248) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1262 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4174), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n991), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3247) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1261 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4174), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n992), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3246) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1260 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4174), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n993), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3245) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1259 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4162), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n954), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3284) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1258 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4162), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n955), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3283) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1257 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4162), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n956), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3282) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1256 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4162), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n957), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3281) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1255 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4163), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n958), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3280) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1254 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4163), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n959), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3279) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1253 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4163), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n960), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3278) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1252 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4163), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n961), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3277) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1251 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4167), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n962), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3276) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1250 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4167), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n963), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3275) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1249 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4167), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n964), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3274) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1248 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4167), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n965), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3273) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1247 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4168), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n966), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3272) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1246 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4168), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n967), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3271) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1245 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4168), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n968), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3270) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1244 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4168), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n969), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3269) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1243 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4169), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n970), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3268) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1242 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4169), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n971), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3267) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1241 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4169), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n972), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3266) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1240 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4169), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n973), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3265) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1239 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4170), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n974), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3264) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1238 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4170), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n975), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3263) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1237 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4170), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n976), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3262) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1236 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4170), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n977), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3261) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1235 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4171), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n978), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3260) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1234 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4171), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n979), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3259) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1233 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4171), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n980), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3258) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1232 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4171), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n981), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3257) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1231 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4172), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n982), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3256) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1230 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4172), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n983), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3255) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1229 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4172), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n984), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3254) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1228 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4172), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n985), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3253) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1227 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4156), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n930), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3308) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1226 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4156), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n931), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3307) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1225 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4156), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n932), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3306) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1224 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4156), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n933), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3305) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1223 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4157), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n934), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3304) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1222 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4157), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n935), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3303) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1221 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4157), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n936), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3302) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1220 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4157), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n937), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3301) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1219 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4158), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n938), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3300) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1218 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4158), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n939), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3299) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1217 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4158), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n940), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3298) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1216 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4158), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n941), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3297) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1215 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4159), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n942), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3296) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1214 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4159), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n943), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3295) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1213 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4159), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n944), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3294) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1212 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4159), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n945), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3293) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1211 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4160), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n946), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3292) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1210 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4160), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n947), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3291) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1209 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4160), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n948), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3290) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1208 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4160), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n949), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3289) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1207 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4161), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n950), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3288) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1206 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4161), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n951), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3287) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1205 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4161), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n952), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3286) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1204 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4161), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n953), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3285) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1203 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4011), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n474), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3444) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1202 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4011), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n475), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3443) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1201 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4011), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n476), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3442) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1200 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4011), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n477), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3441) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1199 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4012), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n478), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3440) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1198 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4012), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n479), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3439) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1197 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4012), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n480), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3438) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1196 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4012), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n481), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3437) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1195 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4000), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n442), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3476) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1194 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4000), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n443), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3475) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1193 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4000), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n444), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3474) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1192 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4000), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n445), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3473) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1191 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4001), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n446), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3472) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1190 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4001), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n447), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3471) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1189 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4001), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n448), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3470) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1188 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4001), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n449), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3469) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1187 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4005), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n450), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3468) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1186 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4005), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n451), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3467) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1185 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4005), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n452), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3466) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1184 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4005), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n453), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3465) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1183 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4006), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n454), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3464) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1182 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4006), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n455), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3463) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1181 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4006), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n456), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3462) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1180 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4006), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n457), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3461) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1179 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4007), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n458), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3460) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1178 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4007), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n459), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3459) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1177 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4007), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n460), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3458) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1176 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4007), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n461), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3457) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1175 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4008), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n462), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3456) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1174 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4008), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n463), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3455) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1173 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4008), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n464), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3454) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1172 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4008), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n465), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3453) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1171 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4009), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n466), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3452) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1170 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4009), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n467), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3451) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1169 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4009), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n468), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3450) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1168 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4009), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n469), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3449) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1167 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4010), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n470), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3448) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1166 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4010), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n471), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3447) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1165 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4010), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n472), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3446) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1164 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4010), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n473), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3445) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1163 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3994), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n418), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3500) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1162 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3994), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n419), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3499) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1161 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3994), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n420), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3498) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1160 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3994), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n421), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3497) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1159 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3995), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n422), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3496) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1158 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3995), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n423), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3495) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1157 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3995), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n424), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3494) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1156 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3995), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n425), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3493) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1155 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3996), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n426), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3492) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1154 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3996), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n427), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3491) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1153 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3996), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n428), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3490) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1152 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3996), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n429), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3489) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1151 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3997), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n430), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3488) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1150 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3997), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n431), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3487) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1149 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3997), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n432), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3486) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1148 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3997), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n433), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3485) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1147 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3998), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n434), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3484) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1146 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3998), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n435), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3483) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1145 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3998), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n436), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3482) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1144 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3998), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n437), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3481) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1143 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3999), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n438), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3480) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1142 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3999), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n439), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3479) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1141 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3999), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n440), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3478) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1140 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3999), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n441), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3477) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1139 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3909), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n154), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3604) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1138 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3909), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n155), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3603) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1137 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3909), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3602) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1136 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3909), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3601) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1135 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3910), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n158), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3600) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1134 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3910), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3599) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1133 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3910), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3598) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1132 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3910), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n161), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3597) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1131 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3920), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n186), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3572) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1130 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3920), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n187), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3571) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1129 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3920), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n188), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3570) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1128 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3920), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n189), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3569) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1127 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3921), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n190), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3568) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1126 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3921), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n191), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3567) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1125 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3921), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n192), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3566) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1124 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3921), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n193), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3565) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1123 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3903), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n130), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3628) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1122 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3903), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n131), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3627) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1121 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3903), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n132), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3626) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1120 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3903), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n133), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3625) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1119 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3904), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n134), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3624) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1118 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3904), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n135), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3623) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1117 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3904), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n136), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3622) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1116 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3904), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n137), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3621) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1115 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3905), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n138), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3620) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1114 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3905), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n139), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3619) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1113 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3905), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n140), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3618) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1112 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3905), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n141), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3617) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1111 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3906), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n142), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3616) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1110 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3906), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n143), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3615) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1109 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3906), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n144), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3614) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1108 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3906), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n145), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3613) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1107 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3907), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n146), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3612) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1106 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3907), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n147), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3611) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1105 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3907), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n148), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3610) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1104 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3907), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n149), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3609) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1103 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3908), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n150), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3608) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1102 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3908), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n151), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3607) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1101 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3908), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n152), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3606) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1100 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3908), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n153), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3605) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1099 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3914), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n162), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3596) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1098 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3914), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n163), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3595) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1097 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3914), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n164), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3594) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1096 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3914), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n165), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3593) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1095 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3915), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n166), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3592) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1094 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3915), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n167), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3591) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1093 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3915), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n168), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3590) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1092 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3915), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n169), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3589) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1091 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3916), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n170), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3588) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1090 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3916), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n171), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3587) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1089 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3916), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n172), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3586) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1088 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3916), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n173), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3585) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1087 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3917), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n174), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3584) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1086 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3917), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n175), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3583) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1085 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3917), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n176), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3582) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1084 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3917), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n177), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3581) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1083 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3918), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n178), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3580) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1082 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3918), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n179), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3579) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1081 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3918), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n180), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3578) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1080 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3918), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n181), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3577) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1079 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3919), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n182), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3576) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1078 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3919), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n183), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3575) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1077 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3919), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n184), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3574) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1076 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3919), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n185), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3573) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1075 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4091), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n730), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3348) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1074 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4091), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n731), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3347) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1073 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4091), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n732), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3346) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1072 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4091), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n733), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3345) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1071 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4092), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n734), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3344) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1070 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4092), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n735), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3343) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1069 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4092), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n736), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3342) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1068 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4092), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n737), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3341) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1067 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4102), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n762), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3316) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1066 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4102), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n763), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3315) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1065 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4102), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n764), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3314) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1064 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4102), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n765), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3313) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1063 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4103), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n766), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3312) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1062 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4103), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n767), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3311) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1061 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4103), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n768), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3310) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1060 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4103), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n769), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3309) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1059 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4085), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n706), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3372) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1058 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4085), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n707), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3371) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1057 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4085), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n708), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3370) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1056 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4085), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n709), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3369) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1055 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4086), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n710), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3368) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1054 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4086), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n711), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3367) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1053 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4086), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n712), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3366) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1052 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4086), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n713), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3365) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1051 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4087), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n714), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3364) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1050 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4087), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n715), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3363) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1049 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4087), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n716), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3362) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1048 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4087), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n717), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3361) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1047 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4088), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n718), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3360) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1046 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4088), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n719), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3359) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1045 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4088), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n720), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3358) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1044 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4088), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n721), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3357) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1043 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4089), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n722), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3356) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1042 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4089), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n723), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3355) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1041 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4089), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n724), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3354) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1040 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4089), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n725), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3353) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1039 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4090), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n726), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3352) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1038 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4090), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n727), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3351) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1037 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4090), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n728), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3350) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1036 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4090), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n729), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3349) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1035 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4096), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n738), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3340) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1034 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4096), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n739), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3339) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1033 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4096), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n740), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3338) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1032 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4096), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n741), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3337) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1031 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4097), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n742), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3336) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1030 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4097), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n743), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3335) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1029 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4097), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n744), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3334) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1028 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4097), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n745), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3333) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1027 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4098), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n746), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3332) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1026 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4098), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n747), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3331) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1025 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4098), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n748), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3330) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1024 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4098), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n749), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3329) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1023 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4099), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n750), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3328) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1022 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4099), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n751), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3327) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1021 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4099), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n752), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3326) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1020 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4099), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n753), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3325) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1019 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4100), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n754), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3324) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1018 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4100), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n755), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3323) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1017 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4100), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n756), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3322) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1016 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4100), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n757), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3321) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1015 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4101), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n758), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3320) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1014 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4101), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n759), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3319) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1013 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4101), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n760), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3318) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1012 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4101), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n761), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3317) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1011 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3867), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n26), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3668) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1010 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3867), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n27), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3667) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1009 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3867), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n28), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3666) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1008 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3867), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n29), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3665) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1007 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3868), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n30), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3664) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1006 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3868), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n31), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3663) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1005 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3868), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n32), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3662) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1004 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3868), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n33), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3661) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1003 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3970), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n346), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3508) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1002 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3970), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n347), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3507) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1001 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3970), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n348), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3506) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U1000 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3970), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n349), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3505) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U999 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3971), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n350), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3504) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U998 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3971), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n351), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3503) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U997 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3971), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n352), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3502) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U996 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3971), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n353), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3501) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U995 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4051), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n602), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3412) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U994 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4051), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n603), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3411) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U993 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4051), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n604), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3410) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U992 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4051), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n605), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3409) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U991 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4052), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n606), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3408) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U990 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4052), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n607), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3407) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U989 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4052), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n608), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3406) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U988 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4052), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n609), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3405) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U987 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4062), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n634), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3380) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U986 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4062), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n635), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3379) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U985 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4062), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n636), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3378) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U984 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4062), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n637), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3377) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U983 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4063), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n638), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3376) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U982 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4063), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n639), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3375) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U981 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4063), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n640), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3374) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U980 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4063), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n641), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3373) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U979 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3878), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n58), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3636) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U978 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3878), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n59), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3635) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U977 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3878), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n60), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3634) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U976 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3878), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n61), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3633) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U975 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3879), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n62), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3632) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U974 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3879), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n63), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3631) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U973 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3879), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n64), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3630) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U972 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3879), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n65), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3629) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U971 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3959), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n314), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3540) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U970 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3959), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n315), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3539) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U969 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3959), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n316), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3538) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U968 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3959), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n317), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3537) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U967 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3960), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n318), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3536) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U966 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3960), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n319), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3535) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U965 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3960), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n320), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3534) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U964 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3960), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n321), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3533) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U963 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4245), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4195), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1050), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3188) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U962 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4244), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4195), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1051), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3187) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U961 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4243), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4195), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1052), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3186) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U960 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4242), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4195), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1053), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3185) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U959 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4241), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4196), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1054), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3184) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U958 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4240), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4196), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1055), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3183) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U957 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4239), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4196), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1056), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3182) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U956 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4238), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4196), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1057), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3181) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U955 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3861), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3692) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U954 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3861), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3691) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U953 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3861), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3690) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U952 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3861), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n5), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3689) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U951 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3862), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n6), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3688) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U950 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3862), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n7), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3687) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U949 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3862), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n8), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3686) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U948 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3862), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n9), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3685) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U947 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3863), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n10), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3684) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U946 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3863), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n11), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3683) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U945 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3863), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n12), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3682) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U944 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3863), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n13), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3681) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U943 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3864), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n14), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3680) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U942 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3864), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n15), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3679) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U941 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3864), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n16), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3678) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U940 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3864), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n17), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3677) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U939 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3865), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n18), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3676) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U938 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3865), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n19), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3675) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U937 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3865), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n20), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3674) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U936 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3865), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n21), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3673) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U935 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3866), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n22), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3672) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U934 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3866), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n23), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3671) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U933 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3866), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n24), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3670) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U932 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3866), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n25), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3669) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U931 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3964), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n322), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3532) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U930 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3964), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n323), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3531) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U929 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3964), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n324), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3530) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U928 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3964), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n325), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3529) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U927 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3965), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n326), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3528) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U926 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3965), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n327), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3527) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U925 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3965), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n328), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3526) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U924 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3965), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n329), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3525) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U923 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3966), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n330), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3524) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U922 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3966), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n331), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3523) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U921 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3966), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n332), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3522) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U920 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3966), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n333), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3521) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U919 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3967), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n334), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3520) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U918 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3967), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n335), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3519) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U917 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3967), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n336), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3518) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U916 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3967), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n337), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3517) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U915 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3968), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n338), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3516) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U914 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3968), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n339), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3515) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U913 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3968), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n340), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3514) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U912 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3968), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n341), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3513) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U911 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3969), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n342), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3512) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U910 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3969), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n343), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3511) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U909 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3969), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n344), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3510) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U908 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3969), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n345), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3509) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U907 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4045), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n578), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3436) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U906 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4045), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n579), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3435) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U905 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4045), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n580), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3434) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U904 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4045), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n581), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3433) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U903 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4046), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n582), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3432) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U902 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4046), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n583), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3431) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U901 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4046), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n584), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3430) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U900 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4046), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n585), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3429) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U899 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4047), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n586), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3428) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U898 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4047), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n587), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3427) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U897 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4047), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n588), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3426) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U896 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4047), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n589), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3425) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U895 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4048), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n590), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3424) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U894 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4048), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n591), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3423) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U893 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4048), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n592), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3422) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U892 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4048), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n593), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3421) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U891 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4049), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n594), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3420) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U890 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4049), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n595), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3419) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U889 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4049), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n596), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3418) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U888 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4049), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n597), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3417) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U887 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4050), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n598), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3416) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U886 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4050), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n599), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3415) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U885 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4050), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n600), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3414) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U884 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4050), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n601), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3413) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U883 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4056), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n610), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3404) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U882 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4056), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n611), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3403) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U881 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4056), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n612), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3402) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U880 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4056), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n613), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3401) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U879 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4057), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n614), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3400) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U878 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4057), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n615), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3399) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U877 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4057), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n616), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3398) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U876 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4057), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n617), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3397) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U875 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4058), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n618), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3396) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U874 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4058), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n619), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3395) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U873 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4058), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n620), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3394) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U872 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4058), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n621), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3393) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U871 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4059), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n622), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3392) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U870 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4059), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n623), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3391) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U869 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4059), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n624), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3390) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U868 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4059), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n625), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3389) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U867 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4060), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n626), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3388) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U866 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4060), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n627), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3387) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U865 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4060), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n628), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3386) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U864 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4060), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n629), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3385) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U863 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4061), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n630), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3384) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U862 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4061), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n631), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3383) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U861 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4061), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n632), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3382) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U860 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4061), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n633), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3381) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U859 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3872), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n34), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3660) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U858 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3872), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n35), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3659) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U857 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3872), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n36), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3658) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U856 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3872), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n37), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3657) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U855 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3873), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n38), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3656) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U854 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3873), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n39), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3655) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U853 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3873), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n40), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3654) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U852 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3873), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n41), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3653) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U851 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3874), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n42), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3652) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U850 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3874), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n43), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3651) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U849 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3874), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n44), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3650) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U848 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3874), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n45), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3649) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U847 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3875), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n46), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3648) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U846 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3875), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n47), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3647) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U845 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3875), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n48), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3646) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U844 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3875), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n49), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3645) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U843 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3876), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n50), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3644) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U842 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3876), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n51), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3643) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U841 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3876), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n52), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3642) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U840 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3876), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n53), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3641) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U839 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3877), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n54), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3640) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U838 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3877), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n55), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3639) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U837 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3877), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n56), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3638) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U836 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3877), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n57), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3637) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U835 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3953), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n290), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3564) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U834 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3953), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n291), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3563) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U833 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3953), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n292), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3562) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U832 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3953), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n293), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3561) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U831 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3954), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n294), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3560) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U830 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3954), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n295), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3559) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U829 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3954), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n296), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3558) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U828 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3954), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n297), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3557) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U827 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3955), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n298), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3556) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U826 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3955), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n299), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3555) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U825 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3955), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n300), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3554) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U824 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3955), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n301), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3553) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U823 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3956), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n302), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3552) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U822 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3956), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n303), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3551) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U821 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3956), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n304), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3550) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U820 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3956), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n305), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3549) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U819 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3957), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n306), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3548) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U818 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3957), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n307), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3547) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U817 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3957), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n308), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3546) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U816 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3957), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n309), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3545) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U815 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3958), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n310), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3544) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U814 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3958), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n311), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3543) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U813 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3958), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n312), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3542) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U812 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3958), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n313), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3541) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U811 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4189), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1026), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3212) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U810 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4189), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1027), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3211) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U809 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4189), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1028), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3210) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U808 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4189), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1029), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3209) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U807 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4190), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1030), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3208) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U806 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4190), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1031), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3207) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U805 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4190), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1032), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3206) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U804 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4190), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1033), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3205) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U803 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4191), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1034), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3204) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U802 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4191), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1035), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3203) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U801 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4191), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1036), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3202) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U800 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4191), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1037), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3201) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U799 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4192), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1038), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3200) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U798 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4192), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1039), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3199) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U797 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4192), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1040), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3198) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U796 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4192), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1041), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3197) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U795 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4193), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1042), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3196) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U794 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4193), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1043), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3195) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U793 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4193), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1044), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3194) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U792 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4193), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1045), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3193) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U791 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4194), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1046), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3192) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U790 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4194), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1047), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3191) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U789 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4247), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4194), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1048), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3190) );
  OAI22_X1 dp_id_stage_regfile_DataPath_Physical_RF_U788 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4246), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188), .B1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4194), .B2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1049), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3189) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U787 ( .A(
        dp_id_stage_regfile_DataPath_addr_rd2_p[3]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1201) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U786 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_N429), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U785 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_N428), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U784 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_N429), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U783 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_N428), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U782 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_N429), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U781 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_N428), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U780 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4234), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[3]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2536) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U779 ( .A(
        dp_id_stage_regfile_DataPath_addr_rd2_p[0]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4270) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U778 ( .A(
        dp_id_stage_regfile_DataPath_addr_rd2_p[1]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4236) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U777 ( .A1(
        dp_id_stage_regfile_DataPath_addr_rd2_p[0]), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[1]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529) );
  NOR3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U776 ( .A1(
        dp_id_stage_regfile_DataPath_addr_rd2_p[3]), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[4]), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n4235), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2548) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U775 ( .A(
        dp_id_stage_regfile_DataPath_mux_wr_out[3]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1192) );
  AND4_X2 dp_id_stage_regfile_DataPath_Physical_RF_U774 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[3]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1342), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1191), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1190), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686) );
  AND4_X2 dp_id_stage_regfile_DataPath_Physical_RF_U773 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[4]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1342), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1192), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1190), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517) );
  AND4_X2 dp_id_stage_regfile_DataPath_Physical_RF_U772 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1342), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1192), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1191), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1190), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823) );
  AND4_X2 dp_id_stage_regfile_DataPath_Physical_RF_U771 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[4]), .A2(
        dp_id_stage_regfile_DataPath_mux_wr_out[3]), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1342), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1190), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U770 ( .A(
        dp_id_stage_regfile_DataPath_addr_rd2_p[4]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4234) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U769 ( .A(
        dp_id_stage_regfile_DataPath_mux_rd_out[4]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1195) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U768 ( .A(
        dp_id_stage_regfile_DataPath_mux_rd_out[3]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1196) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U767 ( .A(
        dp_id_stage_regfile_DataPath_mux_rd_out[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1197) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U766 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2531), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1980) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U765 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2551), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1973) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U764 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2549), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1968) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U763 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2539), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1947) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U762 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2535), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1941) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U761 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2528), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1937) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U760 ( .A1(
        dp_id_stage_regfile_DataPath_addr_rd2_p[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1953) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U759 ( .A1(
        dp_id_stage_regfile_DataPath_mux_rd_out[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2580) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U758 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2531), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1979) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U757 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2535), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1943) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U756 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2535), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1942) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U755 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2528), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1936) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U754 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1954) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U753 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1952) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U752 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2581) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U751 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2579) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U750 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2548), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1969) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U749 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2548), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1967) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U748 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2546), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1963) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U747 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2546), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1962) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U746 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2551), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1976) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U745 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2549), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1971) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U744 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2539), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1945) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U743 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2551), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1975) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U742 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2549), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1970) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U741 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2539), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1944) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U740 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2528), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1939) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U739 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2531), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1934) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U738 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2536), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4235), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2531) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U737 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3179), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3178) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U736 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3163), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3155) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U735 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2536), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2528) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U734 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1195), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[3]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3163) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U733 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1196), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[4]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3179) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U732 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1949) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U731 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2576) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U730 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1201), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[4]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2552) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U729 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4234), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1201), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2538) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U728 ( .A1(
        dp_id_stage_regfile_DataPath_mux_rd_out[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3165), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3166) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U727 ( .A(
        dp_id_stage_regfile_DataPath_mux_rd_out[0]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1199) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U726 ( .A(
        dp_id_stage_regfile_DataPath_mux_rd_out[1]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1198) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U725 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2548), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1964) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U724 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2548), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1965) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U723 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2546), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1959) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U722 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2546), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2529), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1960) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U721 ( .A1(
        dp_id_stage_regfile_DataPath_mux_rd_out[0]), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[1]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U720 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4236), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4270), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533) );
  NOR3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U719 ( .A1(
        dp_id_stage_regfile_DataPath_mux_rd_out[3]), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[4]), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1197), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3175) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U718 ( .A(
        dp_id_stage_regfile_DataPath_mux_wr_out[0]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1194) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U717 ( .A(
        dp_id_stage_regfile_DataPath_mux_wr_out[4]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1191) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U716 ( .A(
        dp_id_stage_regfile_DataPath_mux_wr_out[1]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1193) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U715 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1344), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1654) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U714 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1383), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1690) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U713 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1347), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1825) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U712 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1344), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1791) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U711 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1383), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1553) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U710 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1349), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1520) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U709 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1383), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1351) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U708 ( .A(
        dp_id_stage_regfile_DataPath_mux_wr_out[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1190) );
  AND3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U707 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[1]), .A2(
        dp_id_stage_regfile_DataPath_mux_wr_out[0]), .A3(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1344) );
  AND3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U706 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1194), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1193), .A3(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1383) );
  AND3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U705 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[1]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1194), .A3(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1347) );
  AND3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U704 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[0]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1193), .A3(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1349) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U703 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1341), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1758) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U702 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1341), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1621) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U701 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1341), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1484) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U700 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1305), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1893) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U699 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1270), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1860) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U698 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1270), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1723) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U697 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1305), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1418) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U696 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1270), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1385) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U695 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1339), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1588) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U694 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1339), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1451) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U693 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1270), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1271), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1238) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U692 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1305), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1271), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1273) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U691 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1339), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1271), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1307) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U690 ( .A(dp_n12), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4269) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U689 ( .A(dp_n10), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4268) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U688 ( .A(
        dp_wr_data_id_i[29]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4267) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U687 ( .A(
        dp_wr_data_id_i[28]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4266) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U686 ( .A(dp_n8), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4265) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U685 ( .A(dp_n6), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4264) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U684 ( .A(
        dp_wr_data_id_i[25]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4263) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U683 ( .A(
        dp_wr_data_id_i[24]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4262) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U682 ( .A(
        dp_wr_data_id_i[23]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4261) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U681 ( .A(
        dp_wr_data_id_i[22]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4260) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U680 ( .A(
        dp_wr_data_id_i[21]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4259) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U679 ( .A(
        dp_wr_data_id_i[20]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4258) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U678 ( .A(
        dp_wr_data_id_i[19]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4257) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U677 ( .A(
        dp_wr_data_id_i[18]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4256) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U676 ( .A(
        dp_wr_data_id_i[17]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4255) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U675 ( .A(
        dp_wr_data_id_i[16]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4254) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U674 ( .A(
        dp_wr_data_id_i[15]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4253) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U673 ( .A(
        dp_wr_data_id_i[14]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4252) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U672 ( .A(
        dp_wr_data_id_i[13]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4251) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U671 ( .A(
        dp_wr_data_id_i[12]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4250) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U670 ( .A(
        dp_wr_data_id_i[11]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4249) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U669 ( .A(
        dp_wr_data_id_i[10]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4248) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U668 ( .A(dp_wr_data_id_i[9]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4247) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U667 ( .A(dp_wr_data_id_i[8]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4246) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U666 ( .A(dp_wr_data_id_i[7]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4245) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U665 ( .A(dp_wr_data_id_i[6]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4244) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U664 ( .A(dp_wr_data_id_i[5]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4243) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U663 ( .A(dp_wr_data_id_i[4]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4242) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U662 ( .A(dp_wr_data_id_i[3]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4241) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U661 ( .A(dp_wr_data_id_i[2]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4240) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U660 ( .A(dp_wr_data_id_i[1]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4239) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U659 ( .A(dp_wr_data_id_i[0]), .ZN(dp_id_stage_regfile_DataPath_Physical_RF_n4238) );
  NOR3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U658 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1194), .A2(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1193), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1270) );
  NOR3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U657 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[1]), .A2(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]), .A3(
        dp_id_stage_regfile_DataPath_mux_wr_out[0]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1341) );
  NOR3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U656 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[0]), .A2(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1193), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1305) );
  NOR3_X1 dp_id_stage_regfile_DataPath_Physical_RF_U655 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[1]), .A2(
        dp_id_stage_regfile_DataPath_mux_wr_out[2]), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1194), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1339) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U654 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1173) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U653 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1172) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U652 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2538), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4235), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2535) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U651 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3165), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1197), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3162) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U650 ( .A(
        dp_id_stage_regfile_DataPath_addr_rd2_p[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4235) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U649 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3158), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2607) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U648 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3178), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2600) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U647 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3176), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2595) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U646 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3166), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2574) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U645 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3162), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2568) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U644 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3155), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2564) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U643 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2551), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1978) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U642 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2549), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1974) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U641 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2535), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1948) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U640 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3178), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2605) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U639 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3158), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2606) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U638 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3162), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2570) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U637 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3162), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2569) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U636 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3155), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2563) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U635 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3175), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2596) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U634 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3175), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2594) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U633 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3173), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2590) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U632 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3173), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2589) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U631 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2539), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1950) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U630 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2528), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1938) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U629 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2531), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2533), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1933) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U628 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3166), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2577) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U627 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3155), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2565) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U626 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3178), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2603) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U625 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3176), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2598) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U624 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3166), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2572) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U623 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3178), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2602) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U622 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3176), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2597) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U621 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3166), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2571) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U620 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3155), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2566) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U619 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3158), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2561) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U618 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2552), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n4235), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2549) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U617 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3179), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1197), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3176) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U616 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3163), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1197), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3158) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U615 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n2552), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[2]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2551) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U614 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1195), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1196), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3165) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U613 ( .A1(
        dp_id_stage_regfile_DataPath_addr_rd2_p[2]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n2538), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2539) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U612 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3175), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2591) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U611 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3175), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2592) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U610 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1980), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3753) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U609 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1969), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3780) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U608 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1954), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3807) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U607 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1943), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3834) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U606 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2581), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3699) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U605 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1937), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3849) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U604 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1963), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3795) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U603 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1979), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3756) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U602 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1968), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3783) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U601 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1953), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3810) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U600 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1942), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3837) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U599 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2580), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3702) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U598 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1975), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3765) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U597 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1970), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3777) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U596 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1964), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3792) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U595 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1959), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3804) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U594 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1949), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3819) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U593 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1944), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3831) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U592 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2576), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3711) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U591 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1973), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3771) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U590 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1947), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3825) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U589 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1936), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3852) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U588 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1962), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3798) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U587 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1967), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3786) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U586 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1952), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3813) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U585 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1941), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3840) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U584 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2579), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3705) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U583 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3173), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2586) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U582 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3173), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3156), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2587) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U581 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1976), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3762) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U580 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1971), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3774) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U579 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1965), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3789) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U578 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1960), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3801) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U577 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1945), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3828) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U576 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1939), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3843) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U575 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1934), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3855) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U574 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1980), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3752) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U573 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1969), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3779) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U572 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1954), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3806) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U571 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1943), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3833) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U570 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2581), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3698) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U569 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1980), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3751) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U568 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1969), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3778) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U567 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1954), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3805) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U566 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1943), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3832) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U565 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2581), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3697) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U564 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1963), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3794) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U563 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1937), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3848) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U562 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1963), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3793) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U561 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1937), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3847) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U560 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1979), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3755) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U559 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1968), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3782) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U558 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1953), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3809) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U557 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1942), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3836) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U556 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2580), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3701) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U555 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1979), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3754) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U554 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1968), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3781) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U553 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1953), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3808) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U552 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1942), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3835) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U551 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2580), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3700) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U550 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1975), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3763) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U549 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1970), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3775) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U548 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1964), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3790) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U547 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1959), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3802) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U546 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1949), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3817) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U545 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1944), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3829) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U544 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2576), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3709) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U543 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1975), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3764) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U542 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1970), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3776) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U541 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1964), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3791) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U540 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1959), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3803) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U539 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1949), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3818) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U538 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1944), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3830) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U537 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2576), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3710) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U536 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1973), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3769) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U535 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1962), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3796) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U534 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1947), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3823) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U533 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1936), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3850) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U532 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1973), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3770) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U531 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1962), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3797) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U530 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1947), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3824) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U529 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1936), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3851) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U528 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1967), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3784) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U527 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1952), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3811) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U526 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1941), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3838) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U525 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2579), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3703) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U524 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1967), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3785) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U523 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1952), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3812) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U522 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1941), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3839) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U521 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2579), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3704) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U520 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1976), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3760) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U519 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1971), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3772) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U518 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1965), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3787) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U517 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1960), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3799) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U516 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1945), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3826) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U515 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1939), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3841) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U514 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1934), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3853) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U513 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1976), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3761) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U512 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1971), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3773) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U511 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1965), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3788) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U510 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1960), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3800) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U509 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1945), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3827) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U508 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1939), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3842) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U507 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1934), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3854) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U506 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1198), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1199), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U505 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1654), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4022) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U504 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1690), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3991) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U503 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1825), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3931) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U502 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1791), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3940) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U501 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1553), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4073) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U500 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1520), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4082) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U499 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1238), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4227) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U498 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1273), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4217) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U497 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1307), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4207) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U496 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1351), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4153) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U495 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1758), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3950) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U494 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1621), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4032) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U493 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1484), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4114) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U492 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1893), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3890) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U491 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1860), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3900) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U490 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1723), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3982) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U489 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1418), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4134) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U488 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1385), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4144) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U487 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1588), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4042) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U486 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1451), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4124) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U485 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1654), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4021) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U484 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1654), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4020) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U483 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1654), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4019) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U482 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1654), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4018) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U481 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1654), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4017) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U480 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1654), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4016) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U479 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1351), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4152) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U478 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1351), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4151) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U477 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1351), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4150) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U476 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1351), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4149) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U475 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1351), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4148) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U474 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1351), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4147) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U473 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1690), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3990) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U472 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1690), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3989) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U471 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1690), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3988) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U470 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1690), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3987) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U469 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1690), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3986) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U468 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1690), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3985) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U467 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1173), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1169) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U466 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1172), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1170) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U465 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1172), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1171) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U464 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3176), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2601) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U463 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3162), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2575) );
  NAND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U462 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n3158), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n3160), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2560) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U461 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2607), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1205) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U460 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2596), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1232) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U459 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2570), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3726) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U458 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1974), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3768) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U457 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1948), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3822) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U456 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2564), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3741) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U455 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2590), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1755) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U454 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2606), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1208) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U453 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2595), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1235) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U452 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2569), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3729) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U451 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1938), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3846) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U450 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1933), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3858) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U449 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2602), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1217) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U448 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2597), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1229) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U447 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2591), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1586) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U446 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2586), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3696) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U445 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2571), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3723) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U444 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2565), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3738) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U443 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2600), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1223) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U442 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2574), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3717) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U441 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2563), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3744) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U440 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2589), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1858) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U439 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1978), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3759) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U438 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2605), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1211) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U437 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2594), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1343) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U436 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2568), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3732) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U435 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1950), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3816) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U434 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2603), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1214) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U433 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2598), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1226) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U432 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2592), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1516) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U431 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2587), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3693) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U430 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2577), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3708) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U429 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2572), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3720) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U428 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2566), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3735) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U427 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2561), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3747) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U426 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2607), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1204) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U425 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2596), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1231) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U424 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2570), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3725) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U423 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2607), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1203) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U422 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2596), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1230) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U421 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2570), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3724) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U420 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1974), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3767) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U419 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1948), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3821) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U418 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2590), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1688) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U417 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2564), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3740) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U416 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1974), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3766) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U415 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1948), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3820) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U414 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2590), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1687) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U413 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2564), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3739) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U412 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2606), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1207) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U411 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2595), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1234) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U410 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2569), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3728) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U409 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2606), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1206) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U408 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2595), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1233) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U407 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2569), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3727) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U406 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1938), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3844) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U405 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1933), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3856) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U404 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2602), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1215) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U403 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2597), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1227) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U402 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2591), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1518) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U401 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2586), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3694) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U400 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2571), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3721) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U399 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2565), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3736) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U398 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1938), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3845) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U397 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1933), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3857) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U396 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2602), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1216) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U395 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2597), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1228) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U394 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2591), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1585) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U393 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2586), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3695) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U392 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2571), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3722) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U391 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2565), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3737) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U390 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2600), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1221) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U389 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2589), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1756) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U388 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2574), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3715) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U387 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2563), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3742) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U386 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2600), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1222) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U385 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2589), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1857) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U384 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2574), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3716) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U383 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2563), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3743) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U382 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1978), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3757) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U381 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2605), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1209) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U380 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2594), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1236) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U379 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2568), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3730) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U378 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1978), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3758) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U377 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2605), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1210) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U376 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2594), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1340) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U375 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2568), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3731) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U374 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1950), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3814) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U373 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2603), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1212) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U372 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2598), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1224) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U371 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2592), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1346) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U370 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2587), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1925) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U369 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2577), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3706) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U368 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2572), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3718) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U367 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2566), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3733) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U366 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2561), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3745) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U365 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1950), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3815) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U364 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2603), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1213) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U363 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2598), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1225) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U362 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2592), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1348) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U361 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2587), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1926) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U360 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2577), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3707) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U359 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2572), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3719) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U358 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2566), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3734) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U357 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2561), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3746) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U356 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1161), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4178) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U355 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1161), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4179) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U354 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1161), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4180) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U353 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1161), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4181) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U352 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1161), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4182) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U351 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1161), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4183) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U350 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4178), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4184) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U349 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4179), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4185) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U348 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1160), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4167) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U347 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1160), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4168) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U346 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1160), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4169) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U345 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1160), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4170) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U344 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1160), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4171) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U343 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1160), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4172) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U342 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1159), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4156) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U341 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1159), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4157) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U340 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1159), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4158) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U339 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1159), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4159) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U338 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1159), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4160) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U337 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1159), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4161) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U336 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4167), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4173) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U335 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4168), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4174) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U334 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4156), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4162) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U333 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4157), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4163) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U332 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1158), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4005) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U331 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1158), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4006) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U330 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1158), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4007) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U329 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1158), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4008) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U328 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1158), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4009) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U327 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1158), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4010) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U326 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1157), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3994) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U325 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1157), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3995) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U324 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1157), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3996) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U323 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1157), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3997) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U322 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1157), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3998) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U321 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1157), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3999) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U320 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4005), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4011) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U319 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4006), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4012) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U318 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3994), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4000) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U317 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3995), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4001) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U316 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1156), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3903) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U315 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1156), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3904) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U314 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1156), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3905) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U313 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1156), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3906) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U312 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1156), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3907) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U311 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1156), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3908) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U310 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1155), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3914) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U309 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1155), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3915) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U308 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1155), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3916) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U307 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1155), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3917) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U306 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1155), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3918) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U305 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1155), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3919) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U304 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3903), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3909) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U303 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3904), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3910) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U302 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3914), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3920) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U301 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3915), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3921) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U300 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1154), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4085) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U299 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1154), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4086) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U298 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1154), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4087) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U297 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1154), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4088) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U296 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1154), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4089) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U295 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1154), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4090) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U294 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4096) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U293 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4097) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U292 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4098) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U291 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4099) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U290 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4100) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U289 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4101) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U288 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4085), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4091) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U287 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4086), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4092) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U286 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4096), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4102) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U285 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4097), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4103) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U284 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3864), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3861) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U283 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3865), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3862) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U282 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3866), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3863) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U281 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1168), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3864) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U280 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1168), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3865) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U279 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1168), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3866) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U278 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3967), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3964) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U277 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3968), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3965) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U276 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3969), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3966) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U275 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1167), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3967) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U274 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1167), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3968) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U273 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1167), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3969) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U272 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4048), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4045) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U271 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4049), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4046) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U270 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4050), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4047) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U269 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1166), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4048) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U268 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1166), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4049) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U267 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1166), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4050) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U266 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4059), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4056) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U265 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4060), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4057) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U264 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4061), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4058) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U263 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1165), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4059) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U262 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1165), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4060) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U261 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1165), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4061) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U260 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3875), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3872) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U259 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3876), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3873) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U258 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3877), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3874) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U257 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1164), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3875) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U256 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1164), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3876) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U255 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1164), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3877) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U254 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3956), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3953) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U253 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3957), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3954) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U252 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3958), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3955) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U251 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1163), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3956) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U250 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1163), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3957) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U249 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1163), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3958) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U248 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4192), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4189) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U247 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4193), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4190) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U246 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4194), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4191) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U245 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1162), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4192) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U244 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1162), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4193) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U243 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1162), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4194) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U242 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1161), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4186) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U241 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1160), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4175) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U240 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1159), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4164) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U239 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1158), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4013) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U238 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1157), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4002) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U237 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1156), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3911) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U236 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1155), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3922) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U235 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1154), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4093) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U234 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4104) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U233 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1168), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3869) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U232 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1167), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3972) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U231 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1166), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4053) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U230 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1165), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4064) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U229 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1164), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3880) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U228 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1163), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3961) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U227 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1162), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4197) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U226 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4227), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4219) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U225 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4227), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4218) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U224 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4022), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4015) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U223 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4022), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4014) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U222 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4153), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4146) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U221 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4153), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4145) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U220 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3991), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3984) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U219 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3991), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3983) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U218 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3931), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3924) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U217 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3931), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3923) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U216 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3940), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3933) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U215 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3940), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3932) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U214 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4073), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4066) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U213 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4073), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4065) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U212 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4082), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4075) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U211 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4082), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4074) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U210 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3950), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3942) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U209 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3950), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3941) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U208 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4032), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4024) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U207 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4032), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4023) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U206 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4114), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4106) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U205 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4114), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4105) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U204 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3890), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3882) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U203 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3890), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3881) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U202 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3900), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3892) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U201 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3900), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3891) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U200 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3982), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3974) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U199 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3982), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3973) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U198 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4134), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4126) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U197 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4134), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4125) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U196 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4144), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4136) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U195 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4144), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4135) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U194 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4042), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4034) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U193 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4042), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4033) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U192 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4124), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4116) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U191 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4124), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4115) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U190 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4217), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4209) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U189 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4217), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4208) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U188 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4207), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4199) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U187 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4207), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4198) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U186 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1169), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1189) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U185 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1170), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1200) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U184 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1171), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1202) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U183 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2601), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1220) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U182 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2575), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3714) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U181 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2560), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3750) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U180 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2601), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1219) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U179 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2575), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3713) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U178 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2601), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n1218) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U177 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2575), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3712) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U176 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2560), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3748) );
  BUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U175 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n2560), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3749) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U174 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4186), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4176) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U173 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4186), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4177) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U172 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4175), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4165) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U171 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4175), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4166) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U170 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4164), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4154) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U169 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4164), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4155) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U168 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4013), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4003) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U167 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4013), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4004) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U166 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4002), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3992) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U165 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4002), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3993) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U164 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3911), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3901) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U163 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3911), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3902) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U162 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3922), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3912) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U161 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3922), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3913) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U160 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4093), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4083) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U159 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4093), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4084) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U158 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4104), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4094) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U157 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4104), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4095) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U156 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3869), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3859) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U155 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3869), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3860) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U154 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3972), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3962) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U153 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3972), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3963) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U152 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4053), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4043) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U151 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4053), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4044) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U150 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4064), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4054) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U149 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4064), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4055) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U148 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3880), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3870) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U147 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3880), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3871) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U146 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3961), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3951) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U145 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n3961), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3952) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U144 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4197), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4187) );
  INV_X1 dp_id_stage_regfile_DataPath_Physical_RF_U143 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n4197), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4188) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U142 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4236), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[0]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2532) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U141 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n4270), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[1]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2530) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U140 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1198), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[0]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3159) );
  NOR2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U139 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1199), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[1]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3157) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U138 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1825), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3930) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U137 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1825), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3929) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U136 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1825), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3928) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U135 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1825), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3927) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U134 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1825), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3926) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U133 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1825), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3925) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U132 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1791), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3939) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U131 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1791), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3938) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U130 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1791), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3937) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U129 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1791), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3936) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U128 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1791), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3935) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U127 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1791), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3934) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U126 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1553), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4072) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U125 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1553), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4071) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U124 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1553), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4070) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U123 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1553), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4069) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U122 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1553), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4068) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U121 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1553), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4067) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U120 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1520), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4081) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U119 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1520), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4080) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U118 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1520), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4079) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U117 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1520), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4078) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U116 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1520), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4077) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U115 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1520), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4076) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U114 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1758), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3949) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U113 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1758), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3948) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U112 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1758), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3947) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U111 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1758), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3946) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U110 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1758), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3945) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U109 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1758), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3944) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U108 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1621), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4031) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U107 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1621), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4030) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U106 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1621), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4029) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U105 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1621), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4028) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U104 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1621), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4027) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U103 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1621), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4026) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U102 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1484), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4113) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U101 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1484), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4112) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U100 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1484), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4111) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U99 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1484), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4110) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U98 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1484), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4109) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U97 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1484), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4108) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U96 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1893), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3889) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U95 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1893), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3888) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U94 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1893), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3887) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U93 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1893), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3886) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U92 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1893), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3885) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U91 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1893), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3884) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U90 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1860), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3899) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U89 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1860), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3898) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U88 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1860), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3897) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U87 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1860), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3896) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U86 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1860), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3895) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U85 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1860), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3894) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U84 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1723), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3981) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U83 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1723), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3980) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U82 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1723), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3979) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U81 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1723), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3978) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U80 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1723), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3977) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U79 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1723), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3976) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U78 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1418), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4133) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U77 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1418), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4132) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U76 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1418), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4131) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U75 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1418), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4130) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U74 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1418), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4129) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U73 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1418), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4128) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U72 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1385), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4143) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U71 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1385), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4142) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U70 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1385), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4141) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U69 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1385), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4140) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U68 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1385), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4139) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U67 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1385), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4138) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U66 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1588), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4041) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U65 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1588), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4040) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U64 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1588), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4039) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U63 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1588), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4038) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U62 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1588), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4037) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U61 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1588), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4036) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U60 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1451), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4123) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U59 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1451), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4122) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U58 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1451), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4121) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U57 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1451), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4120) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U56 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1451), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4119) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U55 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1451), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4118) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U54 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1273), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4216) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U53 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1273), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4215) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U52 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1273), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4214) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U51 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1273), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4213) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U50 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1273), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4212) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U49 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1273), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4211) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U48 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1307), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4204) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U47 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1307), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4203) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U46 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1307), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4202) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U45 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1307), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4201) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U44 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1238), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4226) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U43 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1238), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4225) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U42 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1238), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4224) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U41 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1238), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4223) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U40 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1238), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4222) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U39 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1238), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4221) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U38 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1307), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4205) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U37 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1307), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4206) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U36 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1168), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3867) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U35 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1168), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3868) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U34 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1167), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3970) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U33 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1167), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3971) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U32 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1166), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4051) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U31 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1166), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4052) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U30 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1165), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4062) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U29 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1165), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4063) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U28 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1164), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3878) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U27 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1164), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3879) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U26 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1163), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3959) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U25 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1163), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n3960) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U24 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1162), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4195) );
  CLKBUF_X1 dp_id_stage_regfile_DataPath_Physical_RF_U23 ( .A(
        dp_id_stage_regfile_DataPath_Physical_RF_n1162), .Z(
        dp_id_stage_regfile_DataPath_Physical_RF_n4196) );
  INV_X32 dp_id_stage_regfile_DataPath_Physical_RF_U22 ( .A(
        dp_id_stage_regfile_rst_rf), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U21 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1341), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1168) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U20 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1305), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1167) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U19 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1305), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1166) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U18 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1270), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1165) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U17 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1339), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1164) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U16 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1339), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1163) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U15 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1341), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1271), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1162) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U14 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1344), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1161) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U13 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1347), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1160) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U12 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1349), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1345), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1159) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U11 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1347), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1158) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U10 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1686), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1349), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1157) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U9 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1383), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1156) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U8 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1823), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1349), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1155) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U7 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1347), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1154) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U6 ( .A1(
        dp_id_stage_regfile_DataPath_Physical_RF_n1517), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1344), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U5 ( .A1(
        dp_id_stage_regfile_DataPath_addr_rd2_p[2]), .A2(
        dp_id_stage_regfile_DataPath_addr_rd2_p[3]), .A3(
        dp_id_stage_regfile_DataPath_addr_rd2_p[4]), .A4(
        dp_id_stage_regfile_DataPath_addr_rd2_p[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2546) );
  NOR4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U4 ( .A1(
        dp_id_stage_regfile_DataPath_mux_rd_out[2]), .A2(
        dp_id_stage_regfile_DataPath_mux_rd_out[3]), .A3(
        dp_id_stage_regfile_DataPath_mux_rd_out[4]), .A4(
        dp_id_stage_regfile_DataPath_mux_rd_out[5]), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3173) );
  AND4_X1 dp_id_stage_regfile_DataPath_Physical_RF_U3 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_out[5]), .A2(
        dp_id_stage_regfile_DataPath_Physical_RF_n1342), .A3(
        dp_id_stage_regfile_DataPath_Physical_RF_n1192), .A4(
        dp_id_stage_regfile_DataPath_Physical_RF_n1191), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1271) );
  AND2_X1 dp_id_stage_regfile_DataPath_Physical_RF_U2 ( .A1(
        dp_id_stage_regfile_DataPath_mux_wr_control_out), .A2(
        dp_id_stage_regfile_DataPath_mux_en_control_out), .ZN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1342) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1089), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1079), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1078), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1077), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1076), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1075), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1074), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1073), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1121), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1111), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1110), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1109), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1108), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1107), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1106), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1105), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1088), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1087), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1086), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1085), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1084), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1083), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1082), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1081), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1080), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1072), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1071), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1070), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1069), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1068), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1067), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1066), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1120), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1119), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1118), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1117), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1116), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1115), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1114), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1113), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1112), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1104), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1103), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1102), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1101), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1100), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1099), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1098), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1153), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1152), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1151), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1150), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1149), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1148), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1147), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1146), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1145), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1144), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1143), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1142), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1141), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1140), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1139), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1138), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1137), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1136), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1135), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1134), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1133), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1132), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1131), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1130), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n577), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n567), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n566), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n565), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n564), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n563), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n562), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n561), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n833), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n823), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n822), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n821), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n820), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n819), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n818), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n817), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n97), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n87), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n86), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n85), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n84), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n83), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n82), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n81), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n129), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n119), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n118), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n117), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n116), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n115), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n114), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n113), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n385), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n375), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n374), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n373), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n372), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n371), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n370), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n369), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n865), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n855), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n854), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n853), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n852), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n851), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n850), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n849), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n897), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n887), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n886), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n885), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n884), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n883), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n882), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n881), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n576), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n575), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n574), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n573), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n572), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n571), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n570), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n569), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n568), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n560), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n559), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n558), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n557), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n556), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n555), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n554), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n832), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n831), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n830), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n829), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n828), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n827), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n826), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n825), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n824), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n816), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n815), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n814), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n813), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n812), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n811), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n810), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n96), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n95), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n94), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n93), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n92), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n91), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n90), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n89), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n88), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n80), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n79), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n78), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n77), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n76), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n75), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n74), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n128), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n127), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n126), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n125), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n124), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n123), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n122), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n121), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n120), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n112), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n111), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n110), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n109), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n108), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n107), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n106), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n384), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n383), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n382), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n381), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n380), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n379), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n378), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n377), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n376), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n368), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n367), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n366), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n365), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n364), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n363), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n362), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n864), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n863), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n862), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n861), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n860), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n859), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n858), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n857), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n856), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n848), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n847), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n846), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n845), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n844), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n843), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n842), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n896), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n895), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n894), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n893), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n892), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n891), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n890), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n889), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n888), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n880), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n879), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n878), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n877), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n876), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n875), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n874), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1063), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1062), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1059), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1058), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1095), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1094), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1091), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1090), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1127), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1126), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1123), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1122), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1065), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1064), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1061), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1060), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1097), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1096), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1093), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1092), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n551), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n550), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n547), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n546), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n807), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n806), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n803), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n802), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n71), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n70), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n67), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n66), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n103), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n102), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n99), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n98), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n359), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n358), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n355), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n354), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n839), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n838), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n835), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n834), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n871), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n870), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n867), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n866), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1129), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1128), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1125), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n1124), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n289), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n279), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n278), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n277), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n276), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n275), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n274), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n273), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n545), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n535), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n534), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n533), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n532), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n531), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n530), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n529), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n801), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n791), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n790), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n789), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n788), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n787), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n786), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n785), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n288), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n287), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n286), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n285), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n284), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n283), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n282), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n281), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n280), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n272), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n271), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n270), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n269), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n268), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n267), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n266), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n544), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n543), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n542), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n541), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n540), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n539), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n538), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n537), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n536), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n528), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n527), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n526), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n525), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n524), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n523), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n522), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n800), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n799), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n798), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n797), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n796), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n795), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n794), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n793), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n792), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n784), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n783), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n782), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n781), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n780), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n779), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n778), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n553), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n552), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n549), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n548), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n809), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n808), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n805), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n804), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n73), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n72), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n69), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n68), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n105), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n104), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n101), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n100), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n361), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n360), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n357), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n356), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n841), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n840), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n837), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n836), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n873), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n872), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n869), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n868), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n263), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n262), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n259), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n258), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n519), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n518), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n515), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n514), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n775), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n774), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n771), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n770), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n265), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n264), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n261), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n260), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n521), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n520), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n517), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n516), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n777), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n776), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n773), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n772), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n417), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n407), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n406), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n405), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n404), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n403), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n402), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n401), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n416), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n415), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n414), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n413), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n412), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n411), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n410), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n409), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n408), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n400), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n399), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n398), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n397), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n396), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n395), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n394), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n929), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n919), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n918), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n917), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n916), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n915), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n914), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n913), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n928), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n927), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n926), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n925), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n924), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n923), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n922), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n921), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n920), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n912), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n911), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n910), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n909), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n908), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n907), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n906), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n673), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n663), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n662), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n661), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n660), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n659), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n658), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n657), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n705), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n695), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n694), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n693), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n692), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n691), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n690), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n689), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n672), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n671), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n670), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n669), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n668), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n667), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n666), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n665), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n664), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n656), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n655), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n654), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n653), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n652), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n651), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n650), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n704), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n703), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n702), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n701), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n700), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n699), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n698), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n697), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n696), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n688), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n687), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n686), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n685), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n684), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n683), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n682), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n225), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n215), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n214), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n213), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n212), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n211), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n210), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n209), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n224), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n223), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n222), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n221), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n220), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n219), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n218), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n217), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n216), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n208), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n207), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n206), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n205), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n204), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n203), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n202), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n257), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n247), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n246), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n245), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n244), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n243), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n242), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n241), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n256), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n255), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n254), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n253), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n252), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n251), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n250), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n249), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n248), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n240), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n239), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n238), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n237), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n236), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n235), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n234), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n391), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n390), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n387), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n386), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n903), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n902), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n899), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n898), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n647), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n646), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n643), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n642), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n679), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n678), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n675), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n674), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n199), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n198), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n195), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n194), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n231), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n230), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n227), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n226), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n393), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n392), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n389), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n388), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n905), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n904), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n901), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n900), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n649), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n648), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n645), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n644), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n681), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n680), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n677), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n676), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n201), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n200), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n197), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n196), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n233), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n232), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n229), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n228), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n513), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__0_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n503), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__10_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n502), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__11_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n501), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__12_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n500), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__13_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n499), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__14_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n498), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__15_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n497), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__16_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n512), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__1_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n511), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__2_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n510), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__3_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n509), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__4_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n508), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__5_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n507), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__6_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n506), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__7_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n505), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__8_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n504), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__9_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n496), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__17_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n495), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__18_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n494), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__19_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n493), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__20_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n492), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__21_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n491), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__22_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n490), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__23_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n487), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__26_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n486), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__27_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n483), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__30_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n482), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__31_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n489), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__24_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n488), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__25_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n485), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__28_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n484), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .Q(
        dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15__29_) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3508), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n346) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3406), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n608) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3407), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n607) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3408), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n606) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3409), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n605) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3410), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n604) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3411), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n603) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3412), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n602) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3374), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n640) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3375), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n639) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3376), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n638) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3377), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n637) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3378), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n636) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3379), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n635) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3380), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n634) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3207), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1031) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3208), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1030) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3211), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1027) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3212), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1026) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3191), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1047) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3192), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1046) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3193), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1045) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3194), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1044) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3195), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1043) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3196), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1042) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3197), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1041) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3189), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1049) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3190), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1048) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3198), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1040) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3199), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1039) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3200), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1038) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3201), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1037) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3202), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1036) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3203), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1035) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3204), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1034) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3205), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1033) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3206), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1032) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3209), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1029) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3210), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1028) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3687), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n7) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3688), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n6) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3691), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n3) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3692), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n2) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3671), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n23) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3672), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n22) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3673), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n21) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3674), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n20) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3675), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n19) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3676), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n18) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3677), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n17) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3669), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n25) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3670), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n24) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3678), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n16) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3679), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n15) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3680), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n14) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3681), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n13) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3682), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n12) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3683), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n11) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3684), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n10) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3685), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n9) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3686), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n8) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3689), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n5) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3690), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3181), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1057) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3182), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1056) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3183), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1055) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3184), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1054) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3185), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1053) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3186), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1052) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3187), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1051) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3188), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1050) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3661), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n33) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3662), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n32) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3663), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n31) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3664), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n30) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3665), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n29) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3666), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n28) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3667), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n27) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3668), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n26) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3367), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n711) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3368), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n710) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3371), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n707) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3372), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n706) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3335), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n743) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3336), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n742) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3339), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n739) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3340), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n738) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3351), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n727) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3352), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n726) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3353), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n725) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3354), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n724) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3355), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n723) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3356), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n722) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3357), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n721) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3319), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n759) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3320), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n758) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3321), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n757) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3322), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n756) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3323), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n755) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3324), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n754) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3325), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n753) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3349), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n729) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3350), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n728) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3358), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n720) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3359), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n719) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3360), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n718) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3361), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n717) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3362), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n716) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3363), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n715) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3364), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n714) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3365), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n713) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3366), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n712) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3369), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n709) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3370), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n708) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3317), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n761) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3318), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n760) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3326), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n752) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3327), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n751) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3328), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n750) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3329), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n749) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3330), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n748) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3331), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n747) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3332), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n746) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3333), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n745) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3334), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n744) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3337), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n741) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3338), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n740) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3463), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n455) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3464), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n454) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3467), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n451) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3468), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n450) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3623), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n135) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3624), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n134) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3627), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n131) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3628), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n130) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3591), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n167) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3592), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n166) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3595), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n163) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3596), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n162) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3495), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n423) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3496), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n422) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3499), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n419) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3500), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n418) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3271), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n967) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3272), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n966) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3275), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n963) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3276), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n962) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3303), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n935) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3304), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n934) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3307), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n931) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3308), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n930) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3447), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n471) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3448), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n470) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3449), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n469) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3450), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n468) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3451), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n467) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3452), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n466) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3453), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n465) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3445), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n473) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3446), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n472) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3454), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n464) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3455), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n463) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3456), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n462) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3457), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n461) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3458), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n460) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3459), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n459) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3460), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n458) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3461), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n457) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3462), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n456) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3465), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n453) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3466), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n452) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3607), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n151) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3608), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n150) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3609), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n149) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3610), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n148) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3611), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n147) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3612), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n146) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3613), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n145) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3575), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n183) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3576), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n182) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3577), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n181) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3578), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n180) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3579), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n179) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3580), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n178) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3581), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n177) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3479), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n439) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3480), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n438) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3481), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n437) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3482), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n436) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3483), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n435) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3484), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n434) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3485), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n433) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3605), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n153) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3606), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n152) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3614), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n144) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3615), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n143) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3616), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n142) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3617), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n141) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3618), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n140) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3619), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n139) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3620), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n138) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3621), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n137) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3622), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n136) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3625), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n133) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3626), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n132) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3573), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n185) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3574), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n184) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3582), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n176) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3583), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n175) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3584), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n174) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3585), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n173) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3586), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n172) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3587), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n171) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3588), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n170) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3589), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n169) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3590), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n168) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3593), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n165) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3594), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n164) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3477), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n441) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3478), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n440) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3486), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n432) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3487), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n431) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3488), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n430) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3489), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n429) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3490), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n428) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3491), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n427) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3492), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n426) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3493), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n425) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3494), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n424) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3497), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n421) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3498), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n420) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3255), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n983) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3256), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n982) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3257), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n981) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3258), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n980) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3259), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n979) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3260), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n978) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3261), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n977) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3253), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n985) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3254), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n984) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3262), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n976) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3263), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n975) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3264), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n974) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3265), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n973) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3266), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n972) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3267), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n971) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3268), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n970) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3269), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n969) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3270), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n968) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3273), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n965) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3274), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n964) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3287), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n951) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3288), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n950) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3289), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n949) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3290), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n948) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3291), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n947) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3292), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n946) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3293), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n945) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3285), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n953) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3286), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n952) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3294), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n944) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3295), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n943) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3296), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n942) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3297), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n941) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3298), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n940) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3299), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n939) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3300), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n938) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3301), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n937) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3302), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n936) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3305), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n933) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3306), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n932) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3341), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n737) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3309), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n769) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3342), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n736) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3343), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n735) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3344), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n734) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3345), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n733) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3346), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n732) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3347), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n731) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3348), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n730) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3310), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n768) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3311), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n767) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3312), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n766) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3313), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n765) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3314), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n764) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3315), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n763) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3316), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n762) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3437), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n481) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3438), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n480) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3439), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n479) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3440), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n478) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3441), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n477) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3442), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n476) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3443), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n475) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3444), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n474) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3597), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n161) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3565), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n193) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3469), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n449) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3598), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n160) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3599), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n159) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3600), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n158) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3601), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n157) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3602), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n156) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3603), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n155) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3604), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n154) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3566), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n192) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3567), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n191) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3568), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n190) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3569), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n189) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3570), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n188) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3571), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n187) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3572), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n186) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3470), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n448) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3471), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n447) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3472), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n446) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3473), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n445) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3474), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n444) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3475), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n443) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3476), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n442) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3245), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n993) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3246), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n992) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3247), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n991) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3248), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n990) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3249), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n989) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3250), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n988) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3251), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n987) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3252), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n986) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3277), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n961) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3278), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n960) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3279), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n959) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3280), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n958) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3281), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n957) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3282), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n956) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3283), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n955) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3284), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n954) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3239), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n999) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3240), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n998) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3243), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n995) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3244), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n994) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3223), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1015) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3224), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1014) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3225), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1013) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3226), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1012) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3227), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1011) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3228), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1010) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3229), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1009) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3221), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1017) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3222), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1016) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3230), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1008) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3231), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1007) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3232), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1006) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3233), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1005) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3234), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1004) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3235), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1003) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3236), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1002) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3237), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1001) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3238), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1000) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3241), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n997) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3242), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n996) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3213), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1025) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3214), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1024) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3215), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1023) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3216), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1022) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3217), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1021) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3218), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1020) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3219), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1019) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3220), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n4237), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1018) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_0_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N359), .Q(
        dp_id_stage_out1_i[0]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_0_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N427), .Q(
        dp_id_stage_out2_i[0]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_1_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N358), .Q(
        dp_id_stage_out1_i[1]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_1_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N426), .Q(
        dp_id_stage_out2_i[1]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_2_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N357), .Q(
        dp_id_stage_out1_i[2]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_2_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N425), .Q(
        dp_id_stage_out2_i[2]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_3_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N356), .Q(
        dp_id_stage_out1_i[3]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_3_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N424), .Q(
        dp_id_stage_out2_i[3]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_4_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N355), .Q(
        dp_id_stage_out1_i[4]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_4_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N423), .Q(
        dp_id_stage_out2_i[4]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_5_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N354), .Q(
        dp_id_stage_out1_i[5]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_5_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N422), .Q(
        dp_id_stage_out2_i[5]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_6_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N353), .Q(
        dp_id_stage_out1_i[6]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_6_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N421), .Q(
        dp_id_stage_out2_i[6]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_7_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N352), .Q(
        dp_id_stage_out1_i[7]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_7_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N420), .Q(
        dp_id_stage_out2_i[7]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_8_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N351), .Q(
        dp_id_stage_out1_i[8]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_8_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N419), .Q(
        dp_id_stage_out2_i[8]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_9_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4233), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N350), .Q(
        dp_id_stage_out1_i[9]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_9_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4230), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N418), .Q(
        dp_id_stage_out2_i[9]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_10_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N349), .Q(
        dp_id_stage_out1_i[10]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_10_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N417), .Q(
        dp_id_stage_out2_i[10]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_11_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N348), .Q(
        dp_id_stage_out1_i[11]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_11_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N416), .Q(
        dp_id_stage_out2_i[11]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_12_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N347), .Q(
        dp_id_stage_out1_i[12]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_12_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N415), .Q(
        dp_id_stage_out2_i[12]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_13_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N346), .Q(
        dp_id_stage_out1_i[13]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_13_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N414), .Q(
        dp_id_stage_out2_i[13]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_14_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N345), .Q(
        dp_id_stage_out1_i[14]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_14_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N413), .Q(
        dp_id_stage_out2_i[14]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_15_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N344), .Q(
        dp_id_stage_out1_i[15]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_15_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N412), .Q(
        dp_id_stage_out2_i[15]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_16_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N343), .Q(
        dp_id_stage_out1_i[16]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_16_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N411), .Q(
        dp_id_stage_out2_i[16]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_17_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N342), .Q(
        dp_id_stage_out1_i[17]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_17_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N410), .Q(
        dp_id_stage_out2_i[17]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_18_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N341), .Q(
        dp_id_stage_out1_i[18]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_18_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N409), .Q(
        dp_id_stage_out2_i[18]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_19_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N340), .Q(
        dp_id_stage_out1_i[19]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_19_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N408), .Q(
        dp_id_stage_out2_i[19]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_20_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4232), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N339), .Q(
        dp_id_stage_out1_i[20]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_20_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4229), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N407), .Q(
        dp_id_stage_out2_i[20]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_21_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N338), .Q(
        dp_id_stage_out1_i[21]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_21_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N406), .Q(
        dp_id_stage_out2_i[21]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_22_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N337), .Q(
        dp_id_stage_out1_i[22]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_22_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N405), .Q(
        dp_id_stage_out2_i[22]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_23_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N336), .Q(
        dp_id_stage_out1_i[23]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_23_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N404), .Q(
        dp_id_stage_out2_i[23]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_24_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N335), .Q(
        dp_id_stage_out1_i[24]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_24_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N403), .Q(
        dp_id_stage_out2_i[24]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_25_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N334), .Q(
        dp_id_stage_out1_i[25]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_25_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N402), .Q(
        dp_id_stage_out2_i[25]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_26_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N333), .Q(
        dp_id_stage_out1_i[26]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_26_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N401), .Q(
        dp_id_stage_out2_i[26]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_27_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N332), .Q(
        dp_id_stage_out1_i[27]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_27_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N400), .Q(
        dp_id_stage_out2_i[27]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_28_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N331), .Q(
        dp_id_stage_out1_i[28]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_28_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N399), .Q(
        dp_id_stage_out2_i[28]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_29_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N330), .Q(
        dp_id_stage_out1_i[29]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_29_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N398), .Q(
        dp_id_stage_out2_i[29]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_30_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N329), .Q(
        dp_id_stage_out1_i[30]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_30_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N397), .Q(
        dp_id_stage_out2_i[30]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_31_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4231), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N328), .Q(
        dp_id_stage_out1_i[31]) );
  DLH_X1 dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_31_ ( .G(
        dp_id_stage_regfile_DataPath_Physical_RF_n4228), .D(
        dp_id_stage_regfile_DataPath_Physical_RF_N396), .Q(
        dp_id_stage_out2_i[31]) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3373), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1171), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n641) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3381), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n633) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3382), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n632) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3383), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n631) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3384), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n630) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3385), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n629) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3386), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n628) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3387), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n627) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3388), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1174), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n626) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3389), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n625) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3390), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n624) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3391), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n623) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3392), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n622) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3393), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n621) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3394), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n620) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3395), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n619) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3396), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n618) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3397), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n617) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3398), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n616) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3399), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n615) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3400), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1175), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n614) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3401), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1176), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n613) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3402), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1176), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n612) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3403), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1176), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n611) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3404), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1176), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n610) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3405), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1176), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n609) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3413), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n601) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3414), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n600) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3415), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n599) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3416), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n598) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3417), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n597) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3418), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n596) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3419), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n595) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3420), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n594) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3421), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n593) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3422), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n592) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3423), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n591) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3424), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1177), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n590) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3425), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n589) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3426), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n588) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3427), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n587) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3428), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n586) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3429), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n585) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3430), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n584) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3431), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n583) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3432), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n582) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3433), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n581) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3434), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n580) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3435), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n579) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3436), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1178), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n578) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3501), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1179), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n353) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3502), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1179), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n352) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3503), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1179), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n351) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3504), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1179), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n350) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3505), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n349) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3506), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n348) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3507), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n347) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3509), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n345) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3510), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n344) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3511), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n343) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3512), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n342) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3513), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n341) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3514), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n340) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3515), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n339) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3516), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1180), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n338) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3517), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n337) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3518), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n336) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3519), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n335) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3520), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n334) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3521), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n333) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3522), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n332) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3523), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n331) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3524), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n330) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3525), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n329) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3526), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n328) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3527), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n327) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3528), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1181), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n326) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3529), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n325) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3530), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n324) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3531), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n323) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3532), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n322) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3533), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n321) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3534), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n320) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3535), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n319) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3536), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n318) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3537), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n317) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3538), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n316) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3539), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n315) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3540), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1182), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n314) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3541), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n313) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3542), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n312) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3543), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n311) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3544), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n310) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3545), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n309) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3546), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n308) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3547), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n307) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3548), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n306) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3549), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n305) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3550), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n304) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3551), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n303) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3552), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1183), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n302) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3553), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n301) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3554), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n300) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3555), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n299) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3556), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n298) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3557), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n297) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3558), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n296) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3559), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n295) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3560), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n294) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3561), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n293) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3562), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n292) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3563), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n291) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3564), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1184), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n290) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__0_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3629), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1185), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n65) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__1_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3630), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1185), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n64) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__2_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3631), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1185), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n63) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__3_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3632), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1185), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n62) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__4_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3633), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n61) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__5_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3634), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n60) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__6_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3635), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n59) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__7_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3636), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n58) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__8_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3637), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n57) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__9_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3638), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n56) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__10_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3639), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n55) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__11_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3640), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n54) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__12_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3641), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n53) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__13_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3642), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n52) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__14_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3643), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n51) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__15_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3644), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1186), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n50) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__16_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3645), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n49) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__17_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3646), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n48) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__18_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3647), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n47) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__19_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3648), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n46) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__20_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3649), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n45) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__21_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3650), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n44) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__22_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3651), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n43) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__23_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3652), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n42) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__24_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3653), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n41) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__25_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3654), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n40) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__26_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3655), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n39) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__27_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3656), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1187), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n38) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__28_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3657), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1188), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n37) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__29_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3658), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1188), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n36) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__30_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3659), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1188), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n35) );
  DFFR_X1 dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1__31_ ( .D(
        dp_id_stage_regfile_DataPath_Physical_RF_n3660), .CK(CLK), .RN(
        dp_id_stage_regfile_DataPath_Physical_RF_n1188), .QN(
        dp_id_stage_regfile_DataPath_Physical_RF_n34) );
  NOR4_X1 dp_ex_stage_U11 ( .A1(dp_rf_out1_ex_i[1]), .A2(dp_rf_out1_ex_i[19]), 
        .A3(dp_rf_out1_ex_i[18]), .A4(dp_rf_out1_ex_i[17]), .ZN(dp_ex_stage_n5) );
  NOR4_X1 dp_ex_stage_U10 ( .A1(dp_rf_out1_ex_i[16]), .A2(dp_rf_out1_ex_i[15]), 
        .A3(dp_rf_out1_ex_i[14]), .A4(dp_rf_out1_ex_i[13]), .ZN(dp_ex_stage_n4) );
  NOR4_X1 dp_ex_stage_U9 ( .A1(dp_rf_out1_ex_i[12]), .A2(dp_rf_out1_ex_i[11]), 
        .A3(dp_rf_out1_ex_i[10]), .A4(dp_rf_out1_ex_i[0]), .ZN(dp_ex_stage_n3)
         );
  NAND4_X1 dp_ex_stage_U8 ( .A1(dp_ex_stage_n3), .A2(dp_ex_stage_n4), .A3(
        dp_ex_stage_n5), .A4(dp_ex_stage_n6), .ZN(dp_ex_stage_n2) );
  NAND4_X1 dp_ex_stage_U7 ( .A1(dp_ex_stage_n7), .A2(dp_ex_stage_n8), .A3(
        dp_ex_stage_n9), .A4(dp_ex_stage_n10), .ZN(dp_ex_stage_n1) );
  OR2_X1 dp_ex_stage_U6 ( .A1(dp_ex_stage_n1), .A2(dp_ex_stage_n2), .ZN(
        dp_branch_t_ex_o) );
  NOR4_X1 dp_ex_stage_U5 ( .A1(dp_rf_out1_ex_i[27]), .A2(dp_rf_out1_ex_i[26]), 
        .A3(dp_rf_out1_ex_i[25]), .A4(dp_rf_out1_ex_i[24]), .ZN(dp_ex_stage_n7) );
  NOR4_X1 dp_ex_stage_U4 ( .A1(dp_rf_out1_ex_i[30]), .A2(dp_rf_out1_ex_i[2]), 
        .A3(dp_rf_out1_ex_i[29]), .A4(dp_rf_out1_ex_i[28]), .ZN(dp_ex_stage_n8) );
  NOR4_X1 dp_ex_stage_U3 ( .A1(dp_rf_out1_ex_i[5]), .A2(dp_rf_out1_ex_i[4]), 
        .A3(dp_rf_out1_ex_i[3]), .A4(dp_rf_out1_ex_i[31]), .ZN(dp_ex_stage_n9)
         );
  NOR4_X1 dp_ex_stage_U2 ( .A1(dp_rf_out1_ex_i[9]), .A2(dp_rf_out1_ex_i[8]), 
        .A3(dp_rf_out1_ex_i[7]), .A4(dp_rf_out1_ex_i[6]), .ZN(dp_ex_stage_n10)
         );
  NOR4_X1 dp_ex_stage_U1 ( .A1(dp_rf_out1_ex_i[23]), .A2(dp_rf_out1_ex_i[22]), 
        .A3(dp_rf_out1_ex_i[21]), .A4(dp_rf_out1_ex_i[20]), .ZN(dp_ex_stage_n6) );
  MUX2_X1 dp_ex_stage_muxA_U40 ( .A(dp_rf_out1_ex_i[31]), .B(dp_npc_ex_i[31]), 
        .S(dp_ex_stage_muxA_n2), .Z(dp_ex_stage_muxA_out[31]) );
  MUX2_X1 dp_ex_stage_muxA_U39 ( .A(dp_rf_out1_ex_i[30]), .B(dp_npc_ex_i[30]), 
        .S(dp_ex_stage_muxA_n3), .Z(dp_ex_stage_muxA_out[30]) );
  MUX2_X1 dp_ex_stage_muxA_U38 ( .A(dp_rf_out1_ex_i[29]), .B(dp_npc_ex_i[29]), 
        .S(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_out[29]) );
  MUX2_X1 dp_ex_stage_muxA_U37 ( .A(dp_rf_out1_ex_i[28]), .B(dp_npc_ex_i[28]), 
        .S(dp_ex_stage_muxA_n2), .Z(dp_ex_stage_muxA_out[28]) );
  MUX2_X1 dp_ex_stage_muxA_U36 ( .A(dp_rf_out1_ex_i[27]), .B(dp_npc_ex_i[27]), 
        .S(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_out[27]) );
  MUX2_X1 dp_ex_stage_muxA_U35 ( .A(dp_rf_out1_ex_i[26]), .B(dp_npc_ex_i[26]), 
        .S(dp_ex_stage_muxA_n3), .Z(dp_ex_stage_muxA_out[26]) );
  MUX2_X1 dp_ex_stage_muxA_U34 ( .A(dp_rf_out1_ex_i[25]), .B(dp_npc_ex_i[25]), 
        .S(dp_ex_stage_muxA_n3), .Z(dp_ex_stage_muxA_out[25]) );
  MUX2_X1 dp_ex_stage_muxA_U33 ( .A(dp_rf_out1_ex_i[24]), .B(dp_npc_ex_i[24]), 
        .S(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_out[24]) );
  MUX2_X1 dp_ex_stage_muxA_U32 ( .A(dp_rf_out1_ex_i[23]), .B(dp_npc_ex_i[23]), 
        .S(dp_ex_stage_muxA_n6), .Z(dp_ex_stage_muxA_out[23]) );
  MUX2_X1 dp_ex_stage_muxA_U31 ( .A(dp_rf_out1_ex_i[22]), .B(dp_npc_ex_i[22]), 
        .S(dp_ex_stage_muxA_n6), .Z(dp_ex_stage_muxA_out[22]) );
  MUX2_X1 dp_ex_stage_muxA_U30 ( .A(dp_rf_out1_ex_i[21]), .B(dp_npc_ex_i[21]), 
        .S(dp_ex_stage_muxA_n8), .Z(dp_ex_stage_muxA_out[21]) );
  MUX2_X1 dp_ex_stage_muxA_U29 ( .A(dp_rf_out1_ex_i[20]), .B(dp_npc_ex_i[20]), 
        .S(dp_ex_stage_muxA_n6), .Z(dp_ex_stage_muxA_out[20]) );
  MUX2_X1 dp_ex_stage_muxA_U28 ( .A(dp_rf_out1_ex_i[18]), .B(dp_npc_ex_i[18]), 
        .S(dp_ex_stage_muxA_n5), .Z(dp_ex_stage_muxA_n27) );
  MUX2_X1 dp_ex_stage_muxA_U27 ( .A(dp_rf_out1_ex_i[17]), .B(dp_npc_ex_i[17]), 
        .S(dp_ex_stage_muxA_n8), .Z(dp_ex_stage_muxA_out[17]) );
  MUX2_X1 dp_ex_stage_muxA_U26 ( .A(dp_rf_out1_ex_i[16]), .B(dp_npc_ex_i[16]), 
        .S(dp_ex_stage_muxA_n4), .Z(dp_ex_stage_muxA_out[16]) );
  MUX2_X1 dp_ex_stage_muxA_U25 ( .A(dp_rf_out1_ex_i[15]), .B(dp_npc_ex_i[15]), 
        .S(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_out[15]) );
  MUX2_X1 dp_ex_stage_muxA_U24 ( .A(dp_rf_out1_ex_i[13]), .B(dp_npc_ex_i[13]), 
        .S(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_out[13]) );
  MUX2_X1 dp_ex_stage_muxA_U23 ( .A(dp_rf_out1_ex_i[10]), .B(dp_npc_ex_i[10]), 
        .S(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_out[10]) );
  MUX2_X1 dp_ex_stage_muxA_U22 ( .A(dp_rf_out1_ex_i[9]), .B(dp_npc_ex_i[9]), 
        .S(dp_ex_stage_muxA_n6), .Z(dp_ex_stage_muxA_out[9]) );
  MUX2_X1 dp_ex_stage_muxA_U21 ( .A(dp_rf_out1_ex_i[8]), .B(dp_npc_ex_i[8]), 
        .S(dp_ex_stage_muxA_n8), .Z(dp_ex_stage_muxA_out[8]) );
  MUX2_X1 dp_ex_stage_muxA_U20 ( .A(dp_rf_out1_ex_i[7]), .B(dp_npc_ex_i[7]), 
        .S(dp_ex_stage_muxA_n6), .Z(dp_ex_stage_muxA_out[7]) );
  MUX2_X1 dp_ex_stage_muxA_U19 ( .A(dp_rf_out1_ex_i[6]), .B(dp_npc_ex_i[6]), 
        .S(dp_ex_stage_muxA_n8), .Z(dp_ex_stage_muxA_out[6]) );
  MUX2_X1 dp_ex_stage_muxA_U18 ( .A(dp_rf_out1_ex_i[5]), .B(dp_npc_ex_i[5]), 
        .S(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_out[5]) );
  MUX2_X1 dp_ex_stage_muxA_U17 ( .A(dp_rf_out1_ex_i[4]), .B(dp_npc_ex_i[4]), 
        .S(dp_ex_stage_muxA_n5), .Z(dp_ex_stage_muxA_out[4]) );
  MUX2_X1 dp_ex_stage_muxA_U16 ( .A(dp_rf_out1_ex_i[3]), .B(dp_npc_ex_i[3]), 
        .S(dp_ex_stage_muxA_n8), .Z(dp_ex_stage_muxA_out[3]) );
  MUX2_X1 dp_ex_stage_muxA_U15 ( .A(dp_rf_out1_ex_i[1]), .B(dp_npc_ex_i[1]), 
        .S(dp_ex_stage_muxA_n3), .Z(dp_ex_stage_muxA_out[1]) );
  MUX2_X1 dp_ex_stage_muxA_U14 ( .A(dp_rf_out1_ex_i[0]), .B(dp_npc_ex_i[0]), 
        .S(dp_ex_stage_muxA_n8), .Z(dp_ex_stage_muxA_out[0]) );
  CLKBUF_X3 dp_ex_stage_muxA_U13 ( .A(muxA_sel_i), .Z(dp_ex_stage_muxA_n7) );
  CLKBUF_X1 dp_ex_stage_muxA_U12 ( .A(muxA_sel_i), .Z(dp_ex_stage_muxA_n6) );
  MUX2_X1 dp_ex_stage_muxA_U11 ( .A(dp_rf_out1_ex_i[2]), .B(dp_npc_ex_i[2]), 
        .S(dp_ex_stage_muxA_n8), .Z(dp_ex_stage_muxA_out[2]) );
  BUF_X1 dp_ex_stage_muxA_U10 ( .A(muxA_sel_i), .Z(dp_ex_stage_muxA_n5) );
  CLKBUF_X1 dp_ex_stage_muxA_U9 ( .A(muxA_sel_i), .Z(dp_ex_stage_muxA_n3) );
  MUX2_X1 dp_ex_stage_muxA_U8 ( .A(dp_rf_out1_ex_i[11]), .B(dp_npc_ex_i[11]), 
        .S(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_out[11]) );
  MUX2_X1 dp_ex_stage_muxA_U7 ( .A(dp_rf_out1_ex_i[12]), .B(dp_npc_ex_i[12]), 
        .S(dp_ex_stage_muxA_n3), .Z(dp_ex_stage_muxA_out[12]) );
  BUF_X1 dp_ex_stage_muxA_U6 ( .A(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_n2) );
  CLKBUF_X3 dp_ex_stage_muxA_U5 ( .A(muxA_sel_i), .Z(dp_ex_stage_muxA_n8) );
  BUF_X1 dp_ex_stage_muxA_U4 ( .A(dp_ex_stage_muxA_n7), .Z(dp_ex_stage_muxA_n4) );
  MUX2_X1 dp_ex_stage_muxA_U3 ( .A(dp_rf_out1_ex_i[14]), .B(dp_npc_ex_i[14]), 
        .S(dp_ex_stage_muxA_n5), .Z(dp_ex_stage_muxA_out[14]) );
  BUF_X2 dp_ex_stage_muxA_U2 ( .A(dp_ex_stage_muxA_n27), .Z(
        dp_ex_stage_muxA_out[18]) );
  MUX2_X1 dp_ex_stage_muxA_U1 ( .A(dp_rf_out1_ex_i[19]), .B(dp_npc_ex_i[19]), 
        .S(dp_ex_stage_muxA_n8), .Z(dp_ex_stage_muxA_out[19]) );
  MUX2_X1 dp_ex_stage_muxB_U40 ( .A(dp_data_mem_ex_o[31]), .B(dp_imm_ex_i[31]), 
        .S(dp_ex_stage_muxB_n8), .Z(dp_ex_stage_muxB_out[31]) );
  MUX2_X1 dp_ex_stage_muxB_U39 ( .A(dp_data_mem_ex_o[30]), .B(dp_imm_ex_i[30]), 
        .S(dp_ex_stage_muxB_n8), .Z(dp_ex_stage_muxB_out[30]) );
  MUX2_X1 dp_ex_stage_muxB_U38 ( .A(dp_data_mem_ex_o[29]), .B(dp_imm_ex_i[29]), 
        .S(dp_ex_stage_muxB_n8), .Z(dp_ex_stage_muxB_out[29]) );
  MUX2_X1 dp_ex_stage_muxB_U37 ( .A(dp_data_mem_ex_o[28]), .B(dp_imm_ex_i[28]), 
        .S(dp_ex_stage_muxB_n8), .Z(dp_ex_stage_muxB_out[28]) );
  MUX2_X1 dp_ex_stage_muxB_U36 ( .A(dp_data_mem_ex_o[27]), .B(dp_imm_ex_i[27]), 
        .S(dp_ex_stage_muxB_n8), .Z(dp_ex_stage_muxB_out[27]) );
  MUX2_X1 dp_ex_stage_muxB_U35 ( .A(dp_data_mem_ex_o[26]), .B(dp_imm_ex_i[26]), 
        .S(dp_ex_stage_muxB_n8), .Z(dp_ex_stage_muxB_out[26]) );
  MUX2_X1 dp_ex_stage_muxB_U34 ( .A(dp_data_mem_ex_o[25]), .B(dp_imm_ex_i[25]), 
        .S(dp_ex_stage_muxB_n8), .Z(dp_ex_stage_muxB_out[25]) );
  MUX2_X1 dp_ex_stage_muxB_U33 ( .A(dp_data_mem_ex_o[24]), .B(dp_imm_ex_i[24]), 
        .S(dp_ex_stage_muxB_n8), .Z(dp_ex_stage_muxB_out[24]) );
  MUX2_X1 dp_ex_stage_muxB_U32 ( .A(dp_data_mem_ex_o[23]), .B(dp_imm_ex_i[23]), 
        .S(dp_ex_stage_muxB_n7), .Z(dp_ex_stage_muxB_out[23]) );
  MUX2_X1 dp_ex_stage_muxB_U31 ( .A(dp_data_mem_ex_o[22]), .B(dp_imm_ex_i[22]), 
        .S(dp_ex_stage_muxB_n3), .Z(dp_ex_stage_muxB_out[22]) );
  MUX2_X1 dp_ex_stage_muxB_U30 ( .A(dp_data_mem_ex_o[21]), .B(dp_imm_ex_i[21]), 
        .S(dp_ex_stage_muxB_n3), .Z(dp_ex_stage_muxB_out[21]) );
  MUX2_X1 dp_ex_stage_muxB_U29 ( .A(dp_data_mem_ex_o[20]), .B(dp_imm_ex_i[20]), 
        .S(dp_ex_stage_muxB_n4), .Z(dp_ex_stage_muxB_out[20]) );
  MUX2_X1 dp_ex_stage_muxB_U28 ( .A(dp_data_mem_ex_o[19]), .B(dp_imm_ex_i[19]), 
        .S(dp_ex_stage_muxB_n3), .Z(dp_ex_stage_muxB_out[19]) );
  MUX2_X1 dp_ex_stage_muxB_U27 ( .A(dp_data_mem_ex_o[18]), .B(dp_imm_ex_i[18]), 
        .S(dp_ex_stage_muxB_n7), .Z(dp_ex_stage_muxB_out[18]) );
  MUX2_X1 dp_ex_stage_muxB_U26 ( .A(dp_data_mem_ex_o[17]), .B(dp_imm_ex_i[17]), 
        .S(dp_ex_stage_muxB_n7), .Z(dp_ex_stage_muxB_out[17]) );
  MUX2_X1 dp_ex_stage_muxB_U25 ( .A(dp_data_mem_ex_o[16]), .B(dp_imm_ex_i[16]), 
        .S(dp_ex_stage_muxB_n3), .Z(dp_ex_stage_muxB_out[16]) );
  MUX2_X1 dp_ex_stage_muxB_U24 ( .A(dp_data_mem_ex_o[15]), .B(dp_imm_ex_i[15]), 
        .S(dp_ex_stage_muxB_n2), .Z(dp_ex_stage_muxB_out[15]) );
  MUX2_X1 dp_ex_stage_muxB_U23 ( .A(dp_data_mem_ex_o[14]), .B(dp_imm_ex_i[14]), 
        .S(dp_ex_stage_muxB_n1), .Z(dp_ex_stage_muxB_out[14]) );
  MUX2_X1 dp_ex_stage_muxB_U22 ( .A(dp_data_mem_ex_o[13]), .B(dp_imm_ex_i[13]), 
        .S(dp_ex_stage_muxB_n7), .Z(dp_ex_stage_muxB_out[13]) );
  MUX2_X1 dp_ex_stage_muxB_U21 ( .A(dp_data_mem_ex_o[12]), .B(dp_imm_ex_i[12]), 
        .S(dp_ex_stage_muxB_n3), .Z(dp_ex_stage_muxB_out[12]) );
  MUX2_X1 dp_ex_stage_muxB_U20 ( .A(dp_data_mem_ex_o[11]), .B(dp_imm_ex_i[11]), 
        .S(dp_ex_stage_muxB_n3), .Z(dp_ex_stage_muxB_out[11]) );
  MUX2_X1 dp_ex_stage_muxB_U19 ( .A(dp_data_mem_ex_o[10]), .B(dp_imm_ex_i[10]), 
        .S(dp_ex_stage_muxB_n5), .Z(dp_ex_stage_muxB_out[10]) );
  MUX2_X1 dp_ex_stage_muxB_U18 ( .A(dp_data_mem_ex_o[9]), .B(dp_imm_ex_i[9]), 
        .S(dp_ex_stage_muxB_n3), .Z(dp_ex_stage_muxB_out[9]) );
  MUX2_X1 dp_ex_stage_muxB_U17 ( .A(dp_data_mem_ex_o[8]), .B(dp_imm_ex_i[8]), 
        .S(dp_ex_stage_muxB_n7), .Z(dp_ex_stage_muxB_out[8]) );
  MUX2_X1 dp_ex_stage_muxB_U16 ( .A(dp_data_mem_ex_o[7]), .B(dp_imm_ex_i[7]), 
        .S(dp_ex_stage_muxB_n7), .Z(dp_ex_stage_muxB_out[7]) );
  MUX2_X1 dp_ex_stage_muxB_U15 ( .A(dp_data_mem_ex_o[6]), .B(dp_imm_ex_i[6]), 
        .S(dp_ex_stage_muxB_n5), .Z(dp_ex_stage_muxB_out[6]) );
  MUX2_X1 dp_ex_stage_muxB_U14 ( .A(dp_data_mem_ex_o[5]), .B(dp_imm_ex_i[5]), 
        .S(dp_ex_stage_muxB_n2), .Z(dp_ex_stage_muxB_out[5]) );
  MUX2_X1 dp_ex_stage_muxB_U13 ( .A(dp_data_mem_ex_o[4]), .B(dp_imm_ex_i[4]), 
        .S(dp_ex_stage_muxB_n5), .Z(dp_ex_stage_muxB_out[4]) );
  MUX2_X1 dp_ex_stage_muxB_U12 ( .A(dp_data_mem_ex_o[3]), .B(dp_imm_ex_i[3]), 
        .S(dp_ex_stage_muxB_n7), .Z(dp_ex_stage_muxB_out[3]) );
  MUX2_X1 dp_ex_stage_muxB_U11 ( .A(dp_data_mem_ex_o[2]), .B(dp_imm_ex_i[2]), 
        .S(dp_ex_stage_muxB_n5), .Z(dp_ex_stage_muxB_out[2]) );
  MUX2_X1 dp_ex_stage_muxB_U10 ( .A(dp_data_mem_ex_o[1]), .B(dp_imm_ex_i[1]), 
        .S(muxB_sel_i), .Z(dp_ex_stage_muxB_out[1]) );
  MUX2_X1 dp_ex_stage_muxB_U9 ( .A(dp_data_mem_ex_o[0]), .B(dp_imm_ex_i[0]), 
        .S(muxB_sel_i), .Z(dp_ex_stage_muxB_out[0]) );
  CLKBUF_X1 dp_ex_stage_muxB_U8 ( .A(muxB_sel_i), .Z(dp_ex_stage_muxB_n5) );
  CLKBUF_X1 dp_ex_stage_muxB_U7 ( .A(dp_ex_stage_muxB_n7), .Z(
        dp_ex_stage_muxB_n4) );
  CLKBUF_X3 dp_ex_stage_muxB_U6 ( .A(muxB_sel_i), .Z(dp_ex_stage_muxB_n7) );
  BUF_X1 dp_ex_stage_muxB_U5 ( .A(muxB_sel_i), .Z(dp_ex_stage_muxB_n6) );
  BUF_X2 dp_ex_stage_muxB_U4 ( .A(dp_ex_stage_muxB_n6), .Z(dp_ex_stage_muxB_n3) );
  CLKBUF_X1 dp_ex_stage_muxB_U3 ( .A(dp_ex_stage_muxB_n6), .Z(
        dp_ex_stage_muxB_n2) );
  CLKBUF_X2 dp_ex_stage_muxB_U2 ( .A(dp_ex_stage_muxB_n7), .Z(
        dp_ex_stage_muxB_n8) );
  CLKBUF_X1 dp_ex_stage_muxB_U1 ( .A(dp_ex_stage_muxB_n7), .Z(
        dp_ex_stage_muxB_n1) );
  OAI211_X1 dp_ex_stage_alu_U347 ( .C1(dp_ex_stage_alu_n268), .C2(
        dp_ex_stage_alu_n267), .A(dp_ex_stage_alu_n266), .B(
        dp_ex_stage_alu_n265), .ZN(dp_alu_out_ex_o[0]) );
  AOI21_X1 dp_ex_stage_alu_U346 ( .B1(dp_ex_stage_alu_n263), .B2(
        dp_ex_stage_alu_n189), .A(dp_ex_stage_alu_n262), .ZN(
        dp_ex_stage_alu_n264) );
  INV_X1 dp_ex_stage_alu_U345 ( .A(dp_ex_stage_alu_n21), .ZN(
        dp_ex_stage_alu_n262) );
  MUX2_X1 dp_ex_stage_alu_U344 ( .A(dp_ex_stage_alu_n190), .B(
        dp_ex_stage_alu_n188), .S(dp_ex_stage_alu_n45), .Z(
        dp_ex_stage_alu_n263) );
  MUX2_X1 dp_ex_stage_alu_U343 ( .A(dp_ex_stage_alu_n258), .B(
        dp_ex_stage_alu_n257), .S(dp_ex_stage_alu_n191), .Z(
        dp_ex_stage_alu_n259) );
  AND2_X1 dp_ex_stage_alu_U342 ( .A1(dp_ex_stage_alu_N20), .A2(
        dp_ex_stage_alu_n26), .ZN(dp_ex_stage_alu_n255) );
  NAND2_X1 dp_ex_stage_alu_U341 ( .A1(dp_ex_stage_alu_n254), .A2(
        dp_ex_stage_alu_n26), .ZN(dp_ex_stage_alu_n258) );
  MUX2_X1 dp_ex_stage_alu_U340 ( .A(dp_ex_stage_alu_N17), .B(
        dp_ex_stage_alu_N18), .S(dp_ex_stage_alu_n93), .Z(dp_ex_stage_alu_n254) );
  OAI21_X1 dp_ex_stage_alu_U339 ( .B1(dp_ex_stage_alu_n21), .B2(
        dp_ex_stage_alu_n190), .A(dp_ex_stage_alu_n189), .ZN(
        dp_ex_stage_alu_n261) );
  MUX2_X1 dp_ex_stage_alu_U338 ( .A(dp_ex_stage_alu_n253), .B(
        dp_ex_stage_alu_n252), .S(dp_ex_stage_alu_n2), .Z(dp_ex_stage_alu_n268) );
  NAND2_X1 dp_ex_stage_alu_U337 ( .A1(dp_ex_stage_alu_n251), .A2(
        dp_ex_stage_alu_n51), .ZN(dp_ex_stage_alu_n252) );
  INV_X1 dp_ex_stage_alu_U336 ( .A(alu_op_i[1]), .ZN(dp_ex_stage_alu_n271) );
  MUX2_X1 dp_ex_stage_alu_U335 ( .A(dp_ex_stage_alu_N22), .B(
        dp_ex_stage_alu_N21), .S(alu_op_i[0]), .Z(dp_ex_stage_alu_n251) );
  NAND2_X1 dp_ex_stage_alu_U334 ( .A1(dp_ex_stage_alu_N16), .A2(
        dp_ex_stage_alu_n24), .ZN(dp_ex_stage_alu_n253) );
  NAND3_X1 dp_ex_stage_alu_U333 ( .A1(dp_ex_stage_alu_n206), .A2(
        dp_ex_stage_alu_n40), .A3(dp_ex_stage_alu_n250), .ZN(
        dp_ex_stage_alu_n97) );
  OAI21_X1 dp_ex_stage_alu_U332 ( .B1(dp_ex_stage_alu_n24), .B2(
        dp_ex_stage_alu_n267), .A(alu_op_i[4]), .ZN(dp_ex_stage_alu_n250) );
  NAND3_X1 dp_ex_stage_alu_U331 ( .A1(dp_ex_stage_alu_n205), .A2(
        dp_ex_stage_alu_n191), .A3(dp_ex_stage_alu_n61), .ZN(
        dp_ex_stage_alu_n190) );
  NAND2_X1 dp_ex_stage_alu_U330 ( .A1(dp_ex_stage_alu_n205), .A2(
        dp_ex_stage_alu_n54), .ZN(dp_ex_stage_alu_n188) );
  NAND2_X1 dp_ex_stage_alu_U329 ( .A1(dp_ex_stage_alu_n66), .A2(
        dp_ex_stage_alu_n269), .ZN(dp_ex_stage_alu_n189) );
  INV_X1 dp_ex_stage_alu_U328 ( .A(alu_op_i[4]), .ZN(dp_ex_stage_alu_n269) );
  NAND2_X1 dp_ex_stage_alu_U327 ( .A1(dp_ex_stage_alu_n270), .A2(
        dp_ex_stage_alu_n311), .ZN(dp_ex_stage_alu_n267) );
  INV_X2 dp_ex_stage_alu_U326 ( .A(dp_ex_stage_alu_n241), .ZN(
        dp_ex_stage_alu_n240) );
  INV_X1 dp_ex_stage_alu_U325 ( .A(dp_ex_stage_alu_n223), .ZN(
        dp_ex_stage_alu_n222) );
  CLKBUF_X1 dp_ex_stage_alu_U324 ( .A(dp_ex_stage_alu_n310), .Z(
        dp_ex_stage_alu_n215) );
  AOI22_X1 dp_ex_stage_alu_U323 ( .A1(dp_ex_stage_alu_shifter_out[31]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[31]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n118) );
  AOI22_X1 dp_ex_stage_alu_U322 ( .A1(dp_ex_stage_alu_shifter_out[20]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[20]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n154) );
  AOI22_X1 dp_ex_stage_alu_U321 ( .A1(dp_ex_stage_alu_shifter_out[27]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[27]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n133) );
  AOI22_X1 dp_ex_stage_alu_U320 ( .A1(dp_ex_stage_alu_shifter_out[23]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[23]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n145) );
  NAND4_X1 dp_ex_stage_alu_U319 ( .A1(dp_ex_stage_alu_n272), .A2(
        dp_ex_stage_alu_n271), .A3(dp_ex_stage_alu_n270), .A4(
        dp_ex_stage_alu_n27), .ZN(dp_ex_stage_alu_n90) );
  NOR3_X1 dp_ex_stage_alu_U318 ( .A1(dp_ex_stage_alu_n93), .A2(alu_op_i[4]), 
        .A3(dp_ex_stage_alu_n272), .ZN(dp_ex_stage_alu_n205) );
  INV_X1 dp_ex_stage_alu_U317 ( .A(alu_op_i[3]), .ZN(dp_ex_stage_alu_n311) );
  AOI21_X1 dp_ex_stage_alu_U316 ( .B1(dp_ex_stage_alu_n212), .B2(
        dp_ex_stage_alu_n219), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n155) );
  AOI22_X1 dp_ex_stage_alu_U315 ( .A1(dp_ex_stage_alu_shifter_out[26]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[26]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n136) );
  AOI22_X1 dp_ex_stage_alu_U314 ( .A1(dp_ex_stage_alu_shifter_out[25]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[25]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n139) );
  AOI22_X1 dp_ex_stage_alu_U313 ( .A1(dp_ex_stage_alu_shifter_out[21]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[21]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n151) );
  AOI22_X1 dp_ex_stage_alu_U312 ( .A1(dp_ex_stage_alu_shifter_out[12]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[12]), .B2(
        dp_ex_stage_alu_n218), .ZN(dp_ex_stage_alu_n181) );
  OAI221_X1 dp_ex_stage_alu_U311 ( .B1(dp_ex_stage_alu_n179), .B2(
        dp_ex_stage_alu_n230), .C1(dp_ex_stage_alu_n180), .C2(
        dp_ex_stage_alu_n288), .A(dp_ex_stage_alu_n181), .ZN(
        dp_alu_out_ex_o[12]) );
  AOI22_X1 dp_ex_stage_alu_U310 ( .A1(dp_ex_stage_alu_shifter_out[29]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[29]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n127) );
  AOI22_X1 dp_ex_stage_alu_U309 ( .A1(dp_ex_stage_alu_shifter_out[28]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[28]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n130) );
  AOI22_X1 dp_ex_stage_alu_U308 ( .A1(dp_ex_stage_alu_shifter_out[22]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[22]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n148) );
  AOI22_X1 dp_ex_stage_alu_U307 ( .A1(dp_ex_stage_alu_shifter_out[30]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[30]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n121) );
  AOI22_X1 dp_ex_stage_alu_U306 ( .A1(dp_ex_stage_alu_shifter_out[24]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[24]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n142) );
  INV_X1 dp_ex_stage_alu_U305 ( .A(dp_ex_stage_muxB_out[20]), .ZN(
        dp_ex_stage_alu_n296) );
  INV_X1 dp_ex_stage_alu_U304 ( .A(dp_ex_stage_muxA_out[20]), .ZN(
        dp_ex_stage_alu_n278) );
  AOI21_X1 dp_ex_stage_alu_U303 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n296), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n152) );
  OR2_X1 dp_ex_stage_alu_U302 ( .A1(dp_ex_stage_alu_n153), .A2(
        dp_ex_stage_alu_n296), .ZN(dp_ex_stage_alu_n193) );
  OR2_X1 dp_ex_stage_alu_U301 ( .A1(dp_ex_stage_alu_n152), .A2(
        dp_ex_stage_alu_n278), .ZN(dp_ex_stage_alu_n192) );
  INV_X1 dp_ex_stage_alu_U300 ( .A(dp_ex_stage_alu_n311), .ZN(
        dp_ex_stage_alu_n191) );
  CLKBUF_X1 dp_ex_stage_alu_U299 ( .A(alu_op_i[1]), .Z(dp_ex_stage_alu_n93) );
  INV_X1 dp_ex_stage_alu_U298 ( .A(dp_ex_stage_muxB_out[23]), .ZN(
        dp_ex_stage_alu_n299) );
  INV_X1 dp_ex_stage_alu_U297 ( .A(dp_ex_stage_muxA_out[23]), .ZN(
        dp_ex_stage_alu_n242) );
  AOI21_X1 dp_ex_stage_alu_U296 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n299), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n143) );
  OR2_X1 dp_ex_stage_alu_U295 ( .A1(dp_ex_stage_alu_n144), .A2(
        dp_ex_stage_alu_n299), .ZN(dp_ex_stage_alu_n92) );
  OR2_X1 dp_ex_stage_alu_U294 ( .A1(dp_ex_stage_alu_n143), .A2(
        dp_ex_stage_alu_n242), .ZN(dp_ex_stage_alu_n89) );
  INV_X1 dp_ex_stage_alu_U293 ( .A(dp_ex_stage_muxB_out[27]), .ZN(
        dp_ex_stage_alu_n303) );
  INV_X1 dp_ex_stage_alu_U292 ( .A(dp_ex_stage_muxA_out[27]), .ZN(
        dp_ex_stage_alu_n246) );
  AOI21_X1 dp_ex_stage_alu_U291 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n303), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n131) );
  OR2_X1 dp_ex_stage_alu_U290 ( .A1(dp_ex_stage_alu_n132), .A2(
        dp_ex_stage_alu_n303), .ZN(dp_ex_stage_alu_n88) );
  OR2_X1 dp_ex_stage_alu_U289 ( .A1(dp_ex_stage_alu_n131), .A2(
        dp_ex_stage_alu_n246), .ZN(dp_ex_stage_alu_n87) );
  INV_X1 dp_ex_stage_alu_U288 ( .A(dp_ex_stage_muxB_out[26]), .ZN(
        dp_ex_stage_alu_n302) );
  INV_X1 dp_ex_stage_alu_U287 ( .A(dp_ex_stage_muxA_out[26]), .ZN(
        dp_ex_stage_alu_n245) );
  AOI21_X1 dp_ex_stage_alu_U286 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n302), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n134) );
  OR2_X1 dp_ex_stage_alu_U285 ( .A1(dp_ex_stage_alu_n135), .A2(
        dp_ex_stage_alu_n302), .ZN(dp_ex_stage_alu_n86) );
  OR2_X1 dp_ex_stage_alu_U284 ( .A1(dp_ex_stage_alu_n134), .A2(
        dp_ex_stage_alu_n245), .ZN(dp_ex_stage_alu_n85) );
  INV_X1 dp_ex_stage_alu_U283 ( .A(dp_ex_stage_muxB_out[25]), .ZN(
        dp_ex_stage_alu_n301) );
  INV_X1 dp_ex_stage_alu_U282 ( .A(dp_ex_stage_muxA_out[25]), .ZN(
        dp_ex_stage_alu_n244) );
  AOI21_X1 dp_ex_stage_alu_U281 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n301), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n137) );
  OR2_X1 dp_ex_stage_alu_U280 ( .A1(dp_ex_stage_alu_n138), .A2(
        dp_ex_stage_alu_n301), .ZN(dp_ex_stage_alu_n84) );
  OR2_X1 dp_ex_stage_alu_U279 ( .A1(dp_ex_stage_alu_n137), .A2(
        dp_ex_stage_alu_n244), .ZN(dp_ex_stage_alu_n83) );
  INV_X1 dp_ex_stage_alu_U278 ( .A(dp_ex_stage_muxB_out[22]), .ZN(
        dp_ex_stage_alu_n298) );
  INV_X1 dp_ex_stage_alu_U277 ( .A(dp_ex_stage_muxA_out[22]), .ZN(
        dp_ex_stage_alu_n241) );
  AOI21_X1 dp_ex_stage_alu_U276 ( .B1(dp_ex_stage_alu_n212), .B2(
        dp_ex_stage_alu_n298), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n146) );
  OR2_X1 dp_ex_stage_alu_U275 ( .A1(dp_ex_stage_alu_n147), .A2(
        dp_ex_stage_alu_n298), .ZN(dp_ex_stage_alu_n82) );
  OR2_X1 dp_ex_stage_alu_U274 ( .A1(dp_ex_stage_alu_n146), .A2(
        dp_ex_stage_alu_n39), .ZN(dp_ex_stage_alu_n81) );
  INV_X1 dp_ex_stage_alu_U273 ( .A(dp_ex_stage_muxB_out[21]), .ZN(
        dp_ex_stage_alu_n297) );
  INV_X1 dp_ex_stage_alu_U272 ( .A(dp_ex_stage_muxA_out[21]), .ZN(
        dp_ex_stage_alu_n239) );
  AOI21_X1 dp_ex_stage_alu_U271 ( .B1(dp_ex_stage_alu_n212), .B2(
        dp_ex_stage_alu_n297), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n149) );
  OR2_X1 dp_ex_stage_alu_U270 ( .A1(dp_ex_stage_alu_n150), .A2(
        dp_ex_stage_alu_n297), .ZN(dp_ex_stage_alu_n80) );
  OR2_X1 dp_ex_stage_alu_U269 ( .A1(dp_ex_stage_alu_n149), .A2(
        dp_ex_stage_alu_n239), .ZN(dp_ex_stage_alu_n79) );
  INV_X1 dp_ex_stage_alu_U268 ( .A(dp_ex_stage_alu_n71), .ZN(
        dp_ex_stage_alu_n226) );
  INV_X1 dp_ex_stage_alu_U267 ( .A(dp_ex_stage_alu_n34), .ZN(
        dp_ex_stage_alu_n225) );
  INV_X1 dp_ex_stage_alu_U266 ( .A(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_n221) );
  INV_X1 dp_ex_stage_alu_U265 ( .A(dp_ex_stage_alu_n52), .ZN(
        dp_ex_stage_alu_n274) );
  INV_X1 dp_ex_stage_alu_U264 ( .A(dp_ex_stage_alu_n74), .ZN(
        dp_ex_stage_alu_n228) );
  INV_X1 dp_ex_stage_alu_U263 ( .A(dp_ex_stage_alu_n69), .ZN(
        dp_ex_stage_alu_n224) );
  INV_X1 dp_ex_stage_alu_U262 ( .A(dp_ex_stage_alu_n72), .ZN(
        dp_ex_stage_alu_n227) );
  INV_X1 dp_ex_stage_alu_U261 ( .A(dp_ex_stage_alu_n50), .ZN(
        dp_ex_stage_alu_n220) );
  INV_X1 dp_ex_stage_alu_U260 ( .A(dp_ex_stage_alu_n29), .ZN(
        dp_ex_stage_alu_n234) );
  INV_X1 dp_ex_stage_alu_U259 ( .A(dp_ex_stage_muxA_out[16]), .ZN(
        dp_ex_stage_alu_n235) );
  INV_X1 dp_ex_stage_alu_U258 ( .A(dp_ex_stage_muxB_out[1]), .ZN(
        dp_ex_stage_alu_n219) );
  INV_X1 dp_ex_stage_alu_U257 ( .A(dp_ex_stage_alu_n33), .ZN(
        dp_ex_stage_alu_n229) );
  INV_X1 dp_ex_stage_alu_U256 ( .A(dp_ex_stage_muxA_out[14]), .ZN(
        dp_ex_stage_alu_n233) );
  OAI221_X1 dp_ex_stage_alu_U255 ( .B1(dp_ex_stage_alu_n110), .B2(
        dp_ex_stage_alu_n274), .C1(dp_ex_stage_alu_n111), .C2(
        dp_ex_stage_alu_n223), .A(dp_ex_stage_alu_n112), .ZN(
        dp_alu_out_ex_o[4]) );
  INV_X1 dp_ex_stage_alu_U254 ( .A(dp_ex_stage_muxA_out[18]), .ZN(
        dp_ex_stage_alu_n237) );
  INV_X1 dp_ex_stage_alu_U253 ( .A(dp_ex_stage_alu_n78), .ZN(
        dp_ex_stage_alu_n276) );
  OAI221_X1 dp_ex_stage_alu_U252 ( .B1(dp_ex_stage_alu_n104), .B2(
        dp_ex_stage_alu_n276), .C1(dp_ex_stage_alu_n105), .C2(
        dp_ex_stage_alu_n282), .A(dp_ex_stage_alu_n106), .ZN(
        dp_alu_out_ex_o[6]) );
  OAI221_X1 dp_ex_stage_alu_U251 ( .B1(dp_ex_stage_alu_n107), .B2(
        dp_ex_stage_alu_n275), .C1(dp_ex_stage_alu_n108), .C2(
        dp_ex_stage_alu_n281), .A(dp_ex_stage_alu_n109), .ZN(
        dp_alu_out_ex_o[5]) );
  OAI221_X1 dp_ex_stage_alu_U250 ( .B1(dp_ex_stage_alu_n113), .B2(
        dp_ex_stage_alu_n224), .C1(dp_ex_stage_alu_n114), .C2(
        dp_ex_stage_alu_n221), .A(dp_ex_stage_alu_n115), .ZN(
        dp_alu_out_ex_o[3]) );
  OAI221_X1 dp_ex_stage_alu_U249 ( .B1(dp_ex_stage_alu_n164), .B2(
        dp_ex_stage_alu_n236), .C1(dp_ex_stage_alu_n165), .C2(
        dp_ex_stage_alu_n293), .A(dp_ex_stage_alu_n166), .ZN(
        dp_alu_out_ex_o[17]) );
  AOI21_X1 dp_ex_stage_alu_U248 ( .B1(dp_ex_stage_alu_n212), .B2(
        dp_ex_stage_alu_n300), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n140) );
  NAND2_X1 dp_ex_stage_alu_U247 ( .A1(alu_op_i[4]), .A2(dp_ex_stage_alu_n66), 
        .ZN(dp_ex_stage_alu_shift_arith_i) );
  INV_X1 dp_ex_stage_alu_U246 ( .A(dp_ex_stage_muxB_out[4]), .ZN(
        dp_ex_stage_alu_n223) );
  INV_X1 dp_ex_stage_alu_U245 ( .A(dp_ex_stage_muxA_out[17]), .ZN(
        dp_ex_stage_alu_n236) );
  INV_X1 dp_ex_stage_alu_U244 ( .A(dp_ex_stage_alu_n32), .ZN(
        dp_ex_stage_alu_n230) );
  INV_X1 dp_ex_stage_alu_U243 ( .A(dp_ex_stage_muxA_out[24]), .ZN(
        dp_ex_stage_alu_n243) );
  INV_X1 dp_ex_stage_alu_U242 ( .A(dp_ex_stage_muxA_out[31]), .ZN(
        dp_ex_stage_alu_n249) );
  INV_X1 dp_ex_stage_alu_U241 ( .A(dp_ex_stage_muxA_out[28]), .ZN(
        dp_ex_stage_alu_n248) );
  INV_X1 dp_ex_stage_alu_U240 ( .A(alu_op_i[2]), .ZN(dp_ex_stage_alu_n270) );
  INV_X1 dp_ex_stage_alu_U239 ( .A(dp_ex_stage_muxA_out[13]), .ZN(
        dp_ex_stage_alu_n232) );
  AND4_X1 dp_ex_stage_alu_U238 ( .A1(alu_op_i[2]), .A2(alu_op_i[0]), .A3(
        dp_ex_stage_alu_n311), .A4(dp_ex_stage_alu_n269), .ZN(
        dp_ex_stage_alu_n68) );
  AOI21_X1 dp_ex_stage_alu_U237 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n295), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n158) );
  AOI21_X1 dp_ex_stage_alu_U236 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n283), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n101) );
  OAI221_X1 dp_ex_stage_alu_U234 ( .B1(dp_ex_stage_alu_n101), .B2(
        dp_ex_stage_alu_n225), .C1(dp_ex_stage_alu_n102), .C2(
        dp_ex_stage_alu_n283), .A(dp_ex_stage_alu_n103), .ZN(
        dp_alu_out_ex_o[7]) );
  AOI21_X1 dp_ex_stage_alu_U233 ( .B1(dp_ex_stage_alu_n212), .B2(
        dp_ex_stage_alu_n294), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n161) );
  AOI21_X1 dp_ex_stage_alu_U232 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n289), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n176) );
  OAI221_X1 dp_ex_stage_alu_U231 ( .B1(dp_ex_stage_alu_n176), .B2(
        dp_ex_stage_alu_n232), .C1(dp_ex_stage_alu_n177), .C2(
        dp_ex_stage_alu_n289), .A(dp_ex_stage_alu_n178), .ZN(
        dp_alu_out_ex_o[13]) );
  AOI21_X1 dp_ex_stage_alu_U229 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n290), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n173) );
  OAI221_X1 dp_ex_stage_alu_U228 ( .B1(dp_ex_stage_alu_n173), .B2(
        dp_ex_stage_alu_n233), .C1(dp_ex_stage_alu_n174), .C2(
        dp_ex_stage_alu_n290), .A(dp_ex_stage_alu_n175), .ZN(
        dp_alu_out_ex_o[14]) );
  AOI21_X1 dp_ex_stage_alu_U227 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n291), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n170) );
  OAI221_X1 dp_ex_stage_alu_U226 ( .B1(dp_ex_stage_alu_n170), .B2(
        dp_ex_stage_alu_n234), .C1(dp_ex_stage_alu_n171), .C2(
        dp_ex_stage_alu_n291), .A(dp_ex_stage_alu_n172), .ZN(
        dp_alu_out_ex_o[15]) );
  AOI21_X1 dp_ex_stage_alu_U225 ( .B1(dp_ex_stage_alu_n215), .B2(
        dp_ex_stage_alu_n285), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n94) );
  OAI221_X1 dp_ex_stage_alu_U224 ( .B1(dp_ex_stage_alu_n94), .B2(
        dp_ex_stage_alu_n227), .C1(dp_ex_stage_alu_n95), .C2(
        dp_ex_stage_alu_n285), .A(dp_ex_stage_alu_n96), .ZN(dp_alu_out_ex_o[9]) );
  AOI21_X1 dp_ex_stage_alu_U223 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n284), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n98) );
  OAI221_X1 dp_ex_stage_alu_U222 ( .B1(dp_ex_stage_alu_n98), .B2(
        dp_ex_stage_alu_n226), .C1(dp_ex_stage_alu_n99), .C2(
        dp_ex_stage_alu_n284), .A(dp_ex_stage_alu_n100), .ZN(
        dp_alu_out_ex_o[8]) );
  AOI21_X1 dp_ex_stage_alu_U221 ( .B1(dp_ex_stage_alu_n215), .B2(
        dp_ex_stage_alu_n286), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n185) );
  OAI221_X1 dp_ex_stage_alu_U220 ( .B1(dp_ex_stage_alu_n185), .B2(
        dp_ex_stage_alu_n228), .C1(dp_ex_stage_alu_n186), .C2(
        dp_ex_stage_alu_n286), .A(dp_ex_stage_alu_n187), .ZN(
        dp_alu_out_ex_o[10]) );
  AOI21_X1 dp_ex_stage_alu_U219 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n293), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n164) );
  AOI21_X1 dp_ex_stage_alu_U218 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n287), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n182) );
  OAI221_X1 dp_ex_stage_alu_U217 ( .B1(dp_ex_stage_alu_n182), .B2(
        dp_ex_stage_alu_n229), .C1(dp_ex_stage_alu_n183), .C2(
        dp_ex_stage_alu_n287), .A(dp_ex_stage_alu_n184), .ZN(
        dp_alu_out_ex_o[11]) );
  AOI21_X1 dp_ex_stage_alu_U216 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n288), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n179) );
  AOI21_X1 dp_ex_stage_alu_U215 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n292), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n167) );
  OAI221_X1 dp_ex_stage_alu_U214 ( .B1(dp_ex_stage_alu_n167), .B2(
        dp_ex_stage_alu_n235), .C1(dp_ex_stage_alu_n168), .C2(
        dp_ex_stage_alu_n292), .A(dp_ex_stage_alu_n169), .ZN(
        dp_alu_out_ex_o[16]) );
  AOI21_X1 dp_ex_stage_alu_U213 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n281), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n107) );
  AOI21_X1 dp_ex_stage_alu_U212 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n221), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n113) );
  AOI21_X1 dp_ex_stage_alu_U211 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n220), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n122) );
  OAI221_X1 dp_ex_stage_alu_U210 ( .B1(dp_ex_stage_alu_n122), .B2(
        dp_ex_stage_alu_n43), .C1(dp_ex_stage_alu_n123), .C2(
        dp_ex_stage_alu_n220), .A(dp_ex_stage_alu_n124), .ZN(
        dp_alu_out_ex_o[2]) );
  AOI21_X1 dp_ex_stage_alu_U209 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n223), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n110) );
  AOI21_X1 dp_ex_stage_alu_U208 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n306), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n119) );
  AOI21_X1 dp_ex_stage_alu_U207 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n307), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n116) );
  AOI21_X1 dp_ex_stage_alu_U206 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n304), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n128) );
  AOI21_X1 dp_ex_stage_alu_U205 ( .B1(dp_ex_stage_alu_n213), .B2(
        dp_ex_stage_alu_n305), .A(dp_ex_stage_alu_n202), .ZN(
        dp_ex_stage_alu_n125) );
  AOI221_X1 dp_ex_stage_alu_U204 ( .B1(dp_ex_stage_muxA_out[23]), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n242), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n144) );
  AOI221_X1 dp_ex_stage_alu_U203 ( .B1(dp_ex_stage_muxA_out[26]), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n245), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n135) );
  AOI221_X1 dp_ex_stage_alu_U202 ( .B1(dp_ex_stage_alu_n74), .B2(
        dp_ex_stage_alu_n209), .C1(dp_ex_stage_alu_n212), .C2(
        dp_ex_stage_alu_n228), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n186) );
  INV_X1 dp_ex_stage_alu_U201 ( .A(dp_ex_stage_alu_n70), .ZN(
        dp_ex_stage_alu_n275) );
  INV_X1 dp_ex_stage_alu_U200 ( .A(dp_ex_stage_alu_n76), .ZN(
        dp_ex_stage_alu_n273) );
  INV_X1 dp_ex_stage_alu_U199 ( .A(dp_ex_stage_muxB_out[5]), .ZN(
        dp_ex_stage_alu_n281) );
  INV_X1 dp_ex_stage_alu_U198 ( .A(dp_ex_stage_muxB_out[6]), .ZN(
        dp_ex_stage_alu_n282) );
  INV_X1 dp_ex_stage_alu_U197 ( .A(dp_ex_stage_muxB_out[12]), .ZN(
        dp_ex_stage_alu_n288) );
  INV_X1 dp_ex_stage_alu_U196 ( .A(dp_ex_stage_muxB_out[17]), .ZN(
        dp_ex_stage_alu_n293) );
  INV_X1 dp_ex_stage_alu_U195 ( .A(dp_ex_stage_muxB_out[24]), .ZN(
        dp_ex_stage_alu_n300) );
  INV_X1 dp_ex_stage_alu_U194 ( .A(dp_ex_stage_muxB_out[28]), .ZN(
        dp_ex_stage_alu_n304) );
  INV_X1 dp_ex_stage_alu_U193 ( .A(dp_ex_stage_muxB_out[29]), .ZN(
        dp_ex_stage_alu_n305) );
  INV_X1 dp_ex_stage_alu_U192 ( .A(dp_ex_stage_muxB_out[7]), .ZN(
        dp_ex_stage_alu_n283) );
  INV_X1 dp_ex_stage_alu_U191 ( .A(dp_ex_stage_muxB_out[8]), .ZN(
        dp_ex_stage_alu_n284) );
  INV_X1 dp_ex_stage_alu_U190 ( .A(dp_ex_stage_alu_n35), .ZN(
        dp_ex_stage_alu_n286) );
  INV_X1 dp_ex_stage_alu_U189 ( .A(dp_ex_stage_muxB_out[11]), .ZN(
        dp_ex_stage_alu_n287) );
  INV_X1 dp_ex_stage_alu_U188 ( .A(dp_ex_stage_muxB_out[13]), .ZN(
        dp_ex_stage_alu_n289) );
  INV_X1 dp_ex_stage_alu_U187 ( .A(dp_ex_stage_muxB_out[14]), .ZN(
        dp_ex_stage_alu_n290) );
  INV_X1 dp_ex_stage_alu_U186 ( .A(dp_ex_stage_muxB_out[16]), .ZN(
        dp_ex_stage_alu_n292) );
  INV_X1 dp_ex_stage_alu_U185 ( .A(dp_ex_stage_muxB_out[18]), .ZN(
        dp_ex_stage_alu_n294) );
  INV_X1 dp_ex_stage_alu_U184 ( .A(dp_ex_stage_muxB_out[19]), .ZN(
        dp_ex_stage_alu_n295) );
  INV_X1 dp_ex_stage_alu_U183 ( .A(dp_ex_stage_muxB_out[9]), .ZN(
        dp_ex_stage_alu_n285) );
  INV_X1 dp_ex_stage_alu_U182 ( .A(dp_ex_stage_muxB_out[15]), .ZN(
        dp_ex_stage_alu_n291) );
  AND3_X1 dp_ex_stage_alu_U181 ( .A1(dp_ex_stage_alu_n93), .A2(
        dp_ex_stage_alu_n272), .A3(dp_ex_stage_alu_n54), .ZN(
        dp_ex_stage_alu_n66) );
  INV_X1 dp_ex_stage_alu_U180 ( .A(dp_ex_stage_muxB_out[30]), .ZN(
        dp_ex_stage_alu_n306) );
  INV_X1 dp_ex_stage_alu_U179 ( .A(dp_ex_stage_muxB_out[31]), .ZN(
        dp_ex_stage_alu_n307) );
  AND2_X1 dp_ex_stage_alu_U178 ( .A1(dp_ex_stage_alu_n271), .A2(
        dp_ex_stage_alu_n196), .ZN(dp_ex_stage_alu_n208) );
  BUF_X1 dp_ex_stage_alu_U177 ( .A(dp_ex_stage_alu_n97), .Z(
        dp_ex_stage_alu_n217) );
  AOI22_X1 dp_ex_stage_alu_U176 ( .A1(dp_ex_stage_alu_shifter_out[4]), .A2(
        dp_ex_stage_alu_n196), .B1(dp_ex_stage_alu_adder_out[4]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n112) );
  BUF_X1 dp_ex_stage_alu_U175 ( .A(dp_ex_stage_alu_n68), .Z(
        dp_ex_stage_alu_n195) );
  BUF_X1 dp_ex_stage_alu_U174 ( .A(dp_ex_stage_alu_n97), .Z(
        dp_ex_stage_alu_n218) );
  BUF_X1 dp_ex_stage_alu_U173 ( .A(dp_ex_stage_alu_n97), .Z(
        dp_ex_stage_alu_n216) );
  AOI22_X1 dp_ex_stage_alu_U172 ( .A1(dp_ex_stage_alu_shifter_out[8]), .A2(
        dp_ex_stage_alu_n196), .B1(dp_ex_stage_alu_adder_out[8]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n100) );
  AOI22_X1 dp_ex_stage_alu_U171 ( .A1(dp_ex_stage_alu_shifter_out[16]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[16]), .B2(
        dp_ex_stage_alu_n218), .ZN(dp_ex_stage_alu_n169) );
  INV_X1 dp_ex_stage_alu_U170 ( .A(dp_ex_stage_muxA_out[30]), .ZN(
        dp_ex_stage_alu_n280) );
  BUF_X1 dp_ex_stage_alu_U169 ( .A(dp_ex_stage_alu_n68), .Z(
        dp_ex_stage_alu_n196) );
  INV_X1 dp_ex_stage_alu_U168 ( .A(dp_ex_stage_muxA_out[29]), .ZN(
        dp_ex_stage_alu_n279) );
  INV_X1 dp_ex_stage_alu_U167 ( .A(dp_ex_stage_muxA_out[19]), .ZN(
        dp_ex_stage_alu_n277) );
  BUF_X1 dp_ex_stage_alu_U166 ( .A(dp_ex_stage_alu_n68), .Z(
        dp_ex_stage_alu_n194) );
  AOI221_X1 dp_ex_stage_alu_U165 ( .B1(dp_ex_stage_muxA_out[30]), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n280), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n120) );
  AOI221_X1 dp_ex_stage_alu_U164 ( .B1(dp_ex_stage_muxA_out[29]), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n279), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n126) );
  AOI221_X1 dp_ex_stage_alu_U163 ( .B1(dp_ex_stage_alu_n204), .B2(
        dp_ex_stage_alu_n72), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n227), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n95) );
  AOI221_X1 dp_ex_stage_alu_U162 ( .B1(dp_ex_stage_alu_n33), .B2(
        dp_ex_stage_alu_n209), .C1(dp_ex_stage_alu_n212), .C2(
        dp_ex_stage_alu_n229), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n183) );
  AOI221_X1 dp_ex_stage_alu_U161 ( .B1(dp_ex_stage_muxA_out[19]), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n277), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n159) );
  AOI22_X1 dp_ex_stage_alu_U160 ( .A1(dp_ex_stage_alu_shifter_out[15]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[15]), .B2(
        dp_ex_stage_alu_n218), .ZN(dp_ex_stage_alu_n172) );
  INV_X1 dp_ex_stage_alu_U159 ( .A(dp_ex_stage_alu_n189), .ZN(
        dp_ex_stage_alu_n308) );
  INV_X1 dp_ex_stage_alu_U158 ( .A(dp_ex_stage_alu_n188), .ZN(
        dp_ex_stage_alu_n309) );
  AOI22_X1 dp_ex_stage_alu_U157 ( .A1(dp_ex_stage_alu_shifter_out[11]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[11]), .B2(
        dp_ex_stage_alu_n218), .ZN(dp_ex_stage_alu_n184) );
  INV_X1 dp_ex_stage_alu_U156 ( .A(dp_ex_stage_alu_n190), .ZN(
        dp_ex_stage_alu_n310) );
  AOI21_X1 dp_ex_stage_alu_U155 ( .B1(dp_ex_stage_alu_n214), .B2(
        dp_ex_stage_alu_n282), .A(dp_ex_stage_alu_n203), .ZN(
        dp_ex_stage_alu_n104) );
  AOI22_X1 dp_ex_stage_alu_U154 ( .A1(dp_ex_stage_alu_shifter_out[5]), .A2(
        dp_ex_stage_alu_n196), .B1(dp_ex_stage_alu_adder_out[5]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n109) );
  AOI22_X1 dp_ex_stage_alu_U153 ( .A1(dp_ex_stage_alu_shifter_out[3]), .A2(
        dp_ex_stage_alu_n196), .B1(dp_ex_stage_alu_adder_out[3]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n115) );
  AOI22_X1 dp_ex_stage_alu_U152 ( .A1(dp_ex_stage_alu_shifter_out[6]), .A2(
        dp_ex_stage_alu_n196), .B1(dp_ex_stage_alu_adder_out[6]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n106) );
  AOI22_X1 dp_ex_stage_alu_U151 ( .A1(dp_ex_stage_alu_shifter_out[17]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[17]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n166) );
  AOI22_X1 dp_ex_stage_alu_U150 ( .A1(dp_ex_stage_alu_shifter_out[1]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[1]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n157) );
  AOI22_X1 dp_ex_stage_alu_U149 ( .A1(dp_ex_stage_alu_shifter_out[2]), .A2(
        dp_ex_stage_alu_n195), .B1(dp_ex_stage_alu_adder_out[2]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n124) );
  AOI22_X1 dp_ex_stage_alu_U148 ( .A1(dp_ex_stage_alu_shifter_out[7]), .A2(
        dp_ex_stage_alu_n196), .B1(dp_ex_stage_alu_adder_out[7]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n103) );
  AOI22_X1 dp_ex_stage_alu_U147 ( .A1(dp_ex_stage_alu_shifter_out[9]), .A2(
        dp_ex_stage_alu_n196), .B1(dp_ex_stage_alu_adder_out[9]), .B2(
        dp_ex_stage_alu_n216), .ZN(dp_ex_stage_alu_n96) );
  AOI22_X1 dp_ex_stage_alu_U146 ( .A1(dp_ex_stage_alu_shifter_out[18]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[18]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n163) );
  AOI22_X1 dp_ex_stage_alu_U145 ( .A1(dp_ex_stage_alu_shifter_out[13]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[13]), .B2(
        dp_ex_stage_alu_n218), .ZN(dp_ex_stage_alu_n178) );
  AOI22_X1 dp_ex_stage_alu_U144 ( .A1(dp_ex_stage_alu_shifter_out[14]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[14]), .B2(
        dp_ex_stage_alu_n218), .ZN(dp_ex_stage_alu_n175) );
  AOI22_X1 dp_ex_stage_alu_U143 ( .A1(dp_ex_stage_alu_shifter_out[10]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[10]), .B2(
        dp_ex_stage_alu_n218), .ZN(dp_ex_stage_alu_n187) );
  AOI22_X1 dp_ex_stage_alu_U142 ( .A1(dp_ex_stage_alu_shifter_out[19]), .A2(
        dp_ex_stage_alu_n194), .B1(dp_ex_stage_alu_adder_out[19]), .B2(
        dp_ex_stage_alu_n217), .ZN(dp_ex_stage_alu_n160) );
  BUF_X1 dp_ex_stage_alu_U141 ( .A(dp_ex_stage_alu_n308), .Z(
        dp_ex_stage_alu_n198) );
  BUF_X1 dp_ex_stage_alu_U140 ( .A(dp_ex_stage_alu_n308), .Z(
        dp_ex_stage_alu_n197) );
  BUF_X1 dp_ex_stage_alu_U139 ( .A(dp_ex_stage_alu_n309), .Z(
        dp_ex_stage_alu_n209) );
  BUF_X1 dp_ex_stage_alu_U138 ( .A(dp_ex_stage_alu_n309), .Z(
        dp_ex_stage_alu_n207) );
  BUF_X1 dp_ex_stage_alu_U137 ( .A(dp_ex_stage_alu_n309), .Z(
        dp_ex_stage_alu_n204) );
  BUF_X1 dp_ex_stage_alu_U136 ( .A(dp_ex_stage_alu_n310), .Z(
        dp_ex_stage_alu_n211) );
  BUF_X1 dp_ex_stage_alu_U135 ( .A(dp_ex_stage_alu_n310), .Z(
        dp_ex_stage_alu_n213) );
  BUF_X1 dp_ex_stage_alu_U134 ( .A(dp_ex_stage_alu_n310), .Z(
        dp_ex_stage_alu_n212) );
  BUF_X1 dp_ex_stage_alu_U133 ( .A(dp_ex_stage_alu_n310), .Z(
        dp_ex_stage_alu_n210) );
  BUF_X1 dp_ex_stage_alu_U132 ( .A(dp_ex_stage_alu_n310), .Z(
        dp_ex_stage_alu_n214) );
  BUF_X1 dp_ex_stage_alu_U131 ( .A(dp_ex_stage_alu_n197), .Z(
        dp_ex_stage_alu_n200) );
  BUF_X1 dp_ex_stage_alu_U130 ( .A(dp_ex_stage_alu_n197), .Z(
        dp_ex_stage_alu_n201) );
  BUF_X1 dp_ex_stage_alu_U129 ( .A(dp_ex_stage_alu_n198), .Z(
        dp_ex_stage_alu_n202) );
  BUF_X1 dp_ex_stage_alu_U128 ( .A(dp_ex_stage_alu_n197), .Z(
        dp_ex_stage_alu_n199) );
  BUF_X1 dp_ex_stage_alu_U127 ( .A(dp_ex_stage_alu_n198), .Z(
        dp_ex_stage_alu_n203) );
  INV_X2 dp_ex_stage_alu_U126 ( .A(dp_ex_stage_alu_n232), .ZN(
        dp_ex_stage_alu_n231) );
  OR2_X1 dp_ex_stage_alu_U125 ( .A1(dp_ex_stage_alu_n141), .A2(
        dp_ex_stage_alu_n300), .ZN(dp_ex_stage_alu_n65) );
  OR2_X1 dp_ex_stage_alu_U124 ( .A1(dp_ex_stage_alu_n140), .A2(
        dp_ex_stage_alu_n243), .ZN(dp_ex_stage_alu_n64) );
  OR2_X1 dp_ex_stage_alu_U123 ( .A1(dp_ex_stage_alu_n117), .A2(
        dp_ex_stage_alu_n307), .ZN(dp_ex_stage_alu_n63) );
  OR2_X1 dp_ex_stage_alu_U122 ( .A1(dp_ex_stage_alu_n116), .A2(
        dp_ex_stage_alu_n249), .ZN(dp_ex_stage_alu_n62) );
  INV_X1 dp_ex_stage_alu_U121 ( .A(alu_op_i[2]), .ZN(dp_ex_stage_alu_n61) );
  OR2_X1 dp_ex_stage_alu_U120 ( .A1(dp_ex_stage_alu_n126), .A2(
        dp_ex_stage_alu_n305), .ZN(dp_ex_stage_alu_n60) );
  OR2_X1 dp_ex_stage_alu_U119 ( .A1(dp_ex_stage_alu_n125), .A2(
        dp_ex_stage_alu_n279), .ZN(dp_ex_stage_alu_n59) );
  OR2_X1 dp_ex_stage_alu_U118 ( .A1(dp_ex_stage_alu_n120), .A2(
        dp_ex_stage_alu_n306), .ZN(dp_ex_stage_alu_n58) );
  OR2_X1 dp_ex_stage_alu_U117 ( .A1(dp_ex_stage_alu_n119), .A2(
        dp_ex_stage_alu_n280), .ZN(dp_ex_stage_alu_n57) );
  OR2_X1 dp_ex_stage_alu_U116 ( .A1(dp_ex_stage_alu_n129), .A2(
        dp_ex_stage_alu_n304), .ZN(dp_ex_stage_alu_n56) );
  OR2_X1 dp_ex_stage_alu_U115 ( .A1(dp_ex_stage_alu_n128), .A2(
        dp_ex_stage_alu_n248), .ZN(dp_ex_stage_alu_n55) );
  AOI221_X4 dp_ex_stage_alu_U114 ( .B1(dp_ex_stage_alu_n247), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n248), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n129) );
  NOR2_X1 dp_ex_stage_alu_U113 ( .A1(dp_ex_stage_alu_n259), .A2(
        dp_ex_stage_alu_n17), .ZN(dp_ex_stage_alu_n260) );
  NOR2_X1 dp_ex_stage_alu_U112 ( .A1(dp_ex_stage_alu_n260), .A2(
        dp_ex_stage_alu_n53), .ZN(dp_ex_stage_alu_n266) );
  AND2_X1 dp_ex_stage_alu_U111 ( .A1(dp_ex_stage_alu_n45), .A2(
        dp_ex_stage_alu_n261), .ZN(dp_ex_stage_alu_n53) );
  NAND2_X1 dp_ex_stage_alu_U110 ( .A1(dp_ex_stage_alu_n130), .A2(
        dp_ex_stage_alu_n16), .ZN(dp_alu_out_ex_o[28]) );
  NAND2_X1 dp_ex_stage_alu_U109 ( .A1(dp_ex_stage_alu_n133), .A2(
        dp_ex_stage_alu_n15), .ZN(dp_alu_out_ex_o[27]) );
  NAND2_X1 dp_ex_stage_alu_U108 ( .A1(dp_ex_stage_alu_n139), .A2(
        dp_ex_stage_alu_n14), .ZN(dp_alu_out_ex_o[25]) );
  NAND2_X1 dp_ex_stage_alu_U107 ( .A1(dp_ex_stage_alu_n142), .A2(
        dp_ex_stage_alu_n11), .ZN(dp_alu_out_ex_o[24]) );
  NAND2_X1 dp_ex_stage_alu_U106 ( .A1(dp_ex_stage_alu_n145), .A2(
        dp_ex_stage_alu_n6), .ZN(dp_alu_out_ex_o[23]) );
  NAND2_X1 dp_ex_stage_alu_U105 ( .A1(dp_ex_stage_alu_n151), .A2(
        dp_ex_stage_alu_n10), .ZN(dp_alu_out_ex_o[21]) );
  NAND2_X1 dp_ex_stage_alu_U104 ( .A1(dp_ex_stage_alu_n154), .A2(
        dp_ex_stage_alu_n9), .ZN(dp_alu_out_ex_o[20]) );
  NAND2_X1 dp_ex_stage_alu_U103 ( .A1(dp_ex_stage_alu_n118), .A2(
        dp_ex_stage_alu_n7), .ZN(dp_alu_out_ex_o[31]) );
  NAND2_X1 dp_ex_stage_alu_U102 ( .A1(dp_ex_stage_alu_n121), .A2(
        dp_ex_stage_alu_n5), .ZN(dp_alu_out_ex_o[30]) );
  NAND2_X1 dp_ex_stage_alu_U101 ( .A1(dp_ex_stage_alu_n127), .A2(
        dp_ex_stage_alu_n4), .ZN(dp_alu_out_ex_o[29]) );
  NAND2_X1 dp_ex_stage_alu_U100 ( .A1(dp_ex_stage_alu_n136), .A2(
        dp_ex_stage_alu_n3), .ZN(dp_alu_out_ex_o[26]) );
  NAND2_X1 dp_ex_stage_alu_U99 ( .A1(dp_ex_stage_alu_n148), .A2(
        dp_ex_stage_alu_n8), .ZN(dp_alu_out_ex_o[22]) );
  AOI221_X4 dp_ex_stage_alu_U98 ( .B1(dp_ex_stage_alu_n231), .B2(
        dp_ex_stage_alu_n209), .C1(dp_ex_stage_alu_n212), .C2(
        dp_ex_stage_alu_n232), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n177) );
  OAI21_X2 dp_ex_stage_alu_U97 ( .B1(dp_ex_stage_alu_n90), .B2(
        dp_ex_stage_alu_n311), .A(dp_ex_stage_alu_n91), .ZN(
        dp_ex_stage_alu_N23) );
  AOI221_X4 dp_ex_stage_alu_U96 ( .B1(dp_ex_stage_alu_n71), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n226), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n99) );
  BUF_X2 dp_ex_stage_alu_U95 ( .A(dp_ex_stage_muxA_out[9]), .Z(
        dp_ex_stage_alu_n72) );
  NAND3_X1 dp_ex_stage_alu_U94 ( .A1(dp_ex_stage_alu_n47), .A2(
        dp_ex_stage_alu_n48), .A3(dp_ex_stage_alu_n157), .ZN(
        dp_alu_out_ex_o[1]) );
  OR2_X1 dp_ex_stage_alu_U93 ( .A1(dp_ex_stage_alu_n156), .A2(
        dp_ex_stage_alu_n219), .ZN(dp_ex_stage_alu_n48) );
  OR2_X1 dp_ex_stage_alu_U92 ( .A1(dp_ex_stage_alu_n155), .A2(
        dp_ex_stage_alu_n273), .ZN(dp_ex_stage_alu_n47) );
  BUF_X1 dp_ex_stage_alu_U91 ( .A(dp_ex_stage_alu_n30), .Z(dp_ex_stage_alu_n74) );
  BUF_X4 dp_ex_stage_alu_U90 ( .A(dp_ex_stage_muxB_out[0]), .Z(
        dp_ex_stage_alu_n45) );
  BUF_X2 dp_ex_stage_alu_U89 ( .A(dp_ex_stage_muxA_out[1]), .Z(
        dp_ex_stage_alu_n76) );
  INV_X2 dp_ex_stage_alu_U88 ( .A(dp_ex_stage_alu_n43), .ZN(
        dp_ex_stage_alu_n44) );
  INV_X1 dp_ex_stage_alu_U87 ( .A(dp_ex_stage_muxA_out[2]), .ZN(
        dp_ex_stage_alu_n43) );
  AOI221_X4 dp_ex_stage_alu_U86 ( .B1(dp_ex_stage_muxA_out[18]), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n212), .C2(
        dp_ex_stage_alu_n237), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n162) );
  NAND3_X1 dp_ex_stage_alu_U85 ( .A1(dp_ex_stage_alu_n41), .A2(
        dp_ex_stage_alu_n42), .A3(dp_ex_stage_alu_n163), .ZN(
        dp_alu_out_ex_o[18]) );
  OR2_X1 dp_ex_stage_alu_U84 ( .A1(dp_ex_stage_alu_n162), .A2(
        dp_ex_stage_alu_n294), .ZN(dp_ex_stage_alu_n42) );
  OR2_X1 dp_ex_stage_alu_U83 ( .A1(dp_ex_stage_alu_n161), .A2(
        dp_ex_stage_alu_n237), .ZN(dp_ex_stage_alu_n41) );
  NAND4_X1 dp_ex_stage_alu_U82 ( .A1(dp_ex_stage_alu_n26), .A2(
        dp_ex_stage_alu_n271), .A3(dp_ex_stage_alu_n61), .A4(
        dp_ex_stage_alu_n269), .ZN(dp_ex_stage_alu_n40) );
  CLKBUF_X1 dp_ex_stage_alu_U81 ( .A(dp_ex_stage_alu_n241), .Z(
        dp_ex_stage_alu_n39) );
  INV_X2 dp_ex_stage_alu_U80 ( .A(dp_ex_stage_alu_n235), .ZN(
        dp_ex_stage_alu_n38) );
  BUF_X2 dp_ex_stage_alu_U79 ( .A(dp_ex_stage_muxA_out[8]), .Z(
        dp_ex_stage_alu_n71) );
  NOR3_X1 dp_ex_stage_alu_U78 ( .A1(dp_ex_stage_alu_n36), .A2(
        dp_ex_stage_alu_n37), .A3(dp_ex_stage_alu_n264), .ZN(
        dp_ex_stage_alu_n265) );
  AND2_X1 dp_ex_stage_alu_U77 ( .A1(dp_ex_stage_alu_adder_out[0]), .A2(
        dp_ex_stage_alu_n218), .ZN(dp_ex_stage_alu_n37) );
  AND2_X1 dp_ex_stage_alu_U76 ( .A1(dp_ex_stage_alu_shifter_out[0]), .A2(
        dp_ex_stage_alu_n196), .ZN(dp_ex_stage_alu_n36) );
  AOI221_X4 dp_ex_stage_alu_U75 ( .B1(dp_ex_stage_alu_n238), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n239), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n150) );
  INV_X1 dp_ex_stage_alu_U74 ( .A(dp_ex_stage_alu_n248), .ZN(
        dp_ex_stage_alu_n247) );
  BUF_X1 dp_ex_stage_alu_U73 ( .A(dp_ex_stage_muxB_out[2]), .Z(
        dp_ex_stage_alu_n73) );
  CLKBUF_X1 dp_ex_stage_alu_U72 ( .A(dp_ex_stage_muxB_out[10]), .Z(
        dp_ex_stage_alu_n35) );
  BUF_X2 dp_ex_stage_alu_U71 ( .A(dp_ex_stage_muxA_out[11]), .Z(
        dp_ex_stage_alu_n33) );
  CLKBUF_X1 dp_ex_stage_alu_U70 ( .A(dp_ex_stage_muxA_out[12]), .Z(
        dp_ex_stage_alu_n32) );
  CLKBUF_X1 dp_ex_stage_alu_U69 ( .A(dp_ex_stage_muxA_out[5]), .Z(
        dp_ex_stage_alu_n70) );
  BUF_X4 dp_ex_stage_alu_U68 ( .A(dp_ex_stage_muxB_out[3]), .Z(
        dp_ex_stage_alu_n31) );
  INV_X1 dp_ex_stage_alu_U67 ( .A(dp_ex_stage_alu_n239), .ZN(
        dp_ex_stage_alu_n238) );
  CLKBUF_X1 dp_ex_stage_alu_U66 ( .A(dp_ex_stage_muxA_out[10]), .Z(
        dp_ex_stage_alu_n30) );
  BUF_X2 dp_ex_stage_alu_U65 ( .A(dp_ex_stage_muxA_out[6]), .Z(
        dp_ex_stage_alu_n78) );
  BUF_X2 dp_ex_stage_alu_U64 ( .A(dp_ex_stage_muxA_out[3]), .Z(
        dp_ex_stage_alu_n69) );
  BUF_X2 dp_ex_stage_alu_U63 ( .A(dp_ex_stage_muxA_out[15]), .Z(
        dp_ex_stage_alu_n29) );
  AOI221_X4 dp_ex_stage_alu_U62 ( .B1(dp_ex_stage_muxA_out[17]), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n236), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n165) );
  NOR2_X1 dp_ex_stage_alu_U61 ( .A1(dp_ex_stage_alu_n256), .A2(
        dp_ex_stage_alu_n28), .ZN(dp_ex_stage_alu_n257) );
  AND2_X1 dp_ex_stage_alu_U60 ( .A1(dp_ex_stage_alu_N21), .A2(
        dp_ex_stage_alu_n24), .ZN(dp_ex_stage_alu_n28) );
  CLKBUF_X3 dp_ex_stage_alu_U59 ( .A(dp_ex_stage_muxB_out[1]), .Z(
        dp_ex_stage_alu_n46) );
  NOR2_X1 dp_ex_stage_alu_U58 ( .A1(alu_op_i[2]), .A2(alu_op_i[3]), .ZN(
        dp_ex_stage_alu_n54) );
  INV_X1 dp_ex_stage_alu_U57 ( .A(alu_op_i[4]), .ZN(dp_ex_stage_alu_n27) );
  INV_X1 dp_ex_stage_alu_U56 ( .A(alu_op_i[0]), .ZN(dp_ex_stage_alu_n272) );
  CLKBUF_X1 dp_ex_stage_alu_U55 ( .A(dp_ex_stage_alu_n272), .Z(
        dp_ex_stage_alu_n26) );
  INV_X1 dp_ex_stage_alu_U54 ( .A(dp_ex_stage_alu_n278), .ZN(
        dp_ex_stage_alu_n25) );
  AND2_X1 dp_ex_stage_alu_U53 ( .A1(alu_op_i[0]), .A2(alu_op_i[1]), .ZN(
        dp_ex_stage_alu_n67) );
  CLKBUF_X1 dp_ex_stage_alu_U52 ( .A(dp_ex_stage_alu_n67), .Z(
        dp_ex_stage_alu_n24) );
  BUF_X1 dp_ex_stage_alu_U51 ( .A(dp_ex_stage_alu_n23), .Z(dp_ex_stage_alu_n52) );
  BUF_X1 dp_ex_stage_alu_U50 ( .A(dp_ex_stage_muxA_out[4]), .Z(
        dp_ex_stage_alu_n23) );
  BUF_X2 dp_ex_stage_alu_U49 ( .A(dp_ex_stage_muxB_out[3]), .Z(
        dp_ex_stage_alu_n77) );
  INV_X1 dp_ex_stage_alu_U48 ( .A(dp_ex_stage_alu_n93), .ZN(
        dp_ex_stage_alu_n51) );
  CLKBUF_X1 dp_ex_stage_alu_U47 ( .A(dp_ex_stage_muxB_out[4]), .Z(
        dp_ex_stage_alu_n22) );
  BUF_X2 dp_ex_stage_alu_U46 ( .A(dp_ex_stage_muxA_out[0]), .Z(
        dp_ex_stage_alu_shifter_N202) );
  CLKBUF_X1 dp_ex_stage_alu_U45 ( .A(dp_ex_stage_alu_N23), .Z(
        dp_ex_stage_alu_n20) );
  NAND3_X1 dp_ex_stage_alu_U44 ( .A1(dp_ex_stage_alu_n18), .A2(
        dp_ex_stage_alu_n19), .A3(dp_ex_stage_alu_n160), .ZN(
        dp_alu_out_ex_o[19]) );
  OR2_X1 dp_ex_stage_alu_U43 ( .A1(dp_ex_stage_alu_n159), .A2(
        dp_ex_stage_alu_n295), .ZN(dp_ex_stage_alu_n19) );
  OR2_X1 dp_ex_stage_alu_U42 ( .A1(dp_ex_stage_alu_n158), .A2(
        dp_ex_stage_alu_n277), .ZN(dp_ex_stage_alu_n18) );
  CLKBUF_X1 dp_ex_stage_alu_U41 ( .A(dp_ex_stage_muxB_out[2]), .Z(
        dp_ex_stage_alu_n50) );
  BUF_X1 dp_ex_stage_alu_U40 ( .A(dp_ex_stage_muxA_out[0]), .Z(
        dp_ex_stage_alu_n21) );
  OR2_X1 dp_ex_stage_alu_U39 ( .A1(dp_ex_stage_alu_n2), .A2(
        dp_ex_stage_alu_n61), .ZN(dp_ex_stage_alu_n17) );
  AND2_X1 dp_ex_stage_alu_U38 ( .A1(dp_ex_stage_alu_n56), .A2(
        dp_ex_stage_alu_n55), .ZN(dp_ex_stage_alu_n16) );
  AND2_X1 dp_ex_stage_alu_U37 ( .A1(dp_ex_stage_alu_n88), .A2(
        dp_ex_stage_alu_n87), .ZN(dp_ex_stage_alu_n15) );
  AND2_X1 dp_ex_stage_alu_U36 ( .A1(dp_ex_stage_alu_n84), .A2(
        dp_ex_stage_alu_n83), .ZN(dp_ex_stage_alu_n14) );
  AND2_X1 dp_ex_stage_alu_U35 ( .A1(dp_ex_stage_alu_n65), .A2(
        dp_ex_stage_alu_n64), .ZN(dp_ex_stage_alu_n11) );
  AND2_X1 dp_ex_stage_alu_U34 ( .A1(dp_ex_stage_alu_n80), .A2(
        dp_ex_stage_alu_n79), .ZN(dp_ex_stage_alu_n10) );
  AND2_X1 dp_ex_stage_alu_U33 ( .A1(dp_ex_stage_alu_n193), .A2(
        dp_ex_stage_alu_n192), .ZN(dp_ex_stage_alu_n9) );
  AND2_X1 dp_ex_stage_alu_U32 ( .A1(dp_ex_stage_alu_n82), .A2(
        dp_ex_stage_alu_n81), .ZN(dp_ex_stage_alu_n8) );
  AND2_X1 dp_ex_stage_alu_U31 ( .A1(dp_ex_stage_alu_n63), .A2(
        dp_ex_stage_alu_n62), .ZN(dp_ex_stage_alu_n7) );
  AND2_X1 dp_ex_stage_alu_U30 ( .A1(dp_ex_stage_alu_n92), .A2(
        dp_ex_stage_alu_n89), .ZN(dp_ex_stage_alu_n6) );
  AND2_X1 dp_ex_stage_alu_U29 ( .A1(dp_ex_stage_alu_n58), .A2(
        dp_ex_stage_alu_n57), .ZN(dp_ex_stage_alu_n5) );
  AND2_X1 dp_ex_stage_alu_U28 ( .A1(dp_ex_stage_alu_n60), .A2(
        dp_ex_stage_alu_n59), .ZN(dp_ex_stage_alu_n4) );
  AND2_X1 dp_ex_stage_alu_U27 ( .A1(dp_ex_stage_alu_n86), .A2(
        dp_ex_stage_alu_n85), .ZN(dp_ex_stage_alu_n3) );
  CLKBUF_X2 dp_ex_stage_alu_U26 ( .A(dp_ex_stage_muxB_out[2]), .Z(
        dp_ex_stage_alu_n49) );
  INV_X1 dp_ex_stage_alu_U25 ( .A(dp_ex_stage_alu_n269), .ZN(
        dp_ex_stage_alu_n2) );
  INV_X1 dp_ex_stage_alu_U24 ( .A(dp_ex_stage_alu_n248), .ZN(
        dp_ex_stage_alu_n1) );
  AOI221_X1 dp_ex_stage_alu_U23 ( .B1(dp_ex_stage_alu_n76), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n273), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n156) );
  AOI221_X1 dp_ex_stage_alu_U22 ( .B1(dp_ex_stage_alu_n44), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n43), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n123) );
  AOI221_X1 dp_ex_stage_alu_U21 ( .B1(dp_ex_stage_alu_n69), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n224), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n114) );
  AOI221_X1 dp_ex_stage_alu_U20 ( .B1(dp_ex_stage_alu_n52), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n274), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n111) );
  AOI221_X1 dp_ex_stage_alu_U19 ( .B1(dp_ex_stage_alu_n70), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n275), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n108) );
  AOI221_X1 dp_ex_stage_alu_U18 ( .B1(dp_ex_stage_alu_n78), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n276), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n105) );
  AOI221_X1 dp_ex_stage_alu_U17 ( .B1(dp_ex_stage_alu_n34), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n225), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n102) );
  AOI221_X1 dp_ex_stage_alu_U16 ( .B1(dp_ex_stage_alu_n32), .B2(
        dp_ex_stage_alu_n209), .C1(dp_ex_stage_alu_n212), .C2(
        dp_ex_stage_alu_n230), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n180) );
  AOI221_X1 dp_ex_stage_alu_U15 ( .B1(dp_ex_stage_muxA_out[14]), .B2(
        dp_ex_stage_alu_n209), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n233), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n174) );
  AOI221_X1 dp_ex_stage_alu_U14 ( .B1(dp_ex_stage_alu_n29), .B2(
        dp_ex_stage_alu_n209), .C1(dp_ex_stage_alu_n212), .C2(
        dp_ex_stage_alu_n234), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n171) );
  AOI221_X1 dp_ex_stage_alu_U13 ( .B1(dp_ex_stage_alu_n38), .B2(
        dp_ex_stage_alu_n209), .C1(dp_ex_stage_alu_n212), .C2(
        dp_ex_stage_alu_n235), .A(dp_ex_stage_alu_n201), .ZN(
        dp_ex_stage_alu_n168) );
  AOI221_X1 dp_ex_stage_alu_U12 ( .B1(dp_ex_stage_alu_n25), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n278), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n153) );
  AOI221_X1 dp_ex_stage_alu_U11 ( .B1(dp_ex_stage_alu_n240), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n39), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n147) );
  AOI221_X1 dp_ex_stage_alu_U10 ( .B1(dp_ex_stage_muxA_out[24]), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n243), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n141) );
  AOI221_X1 dp_ex_stage_alu_U9 ( .B1(dp_ex_stage_muxA_out[25]), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n244), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n138) );
  AOI221_X1 dp_ex_stage_alu_U8 ( .B1(dp_ex_stage_muxA_out[27]), .B2(
        dp_ex_stage_alu_n207), .C1(dp_ex_stage_alu_n211), .C2(
        dp_ex_stage_alu_n246), .A(dp_ex_stage_alu_n200), .ZN(
        dp_ex_stage_alu_n132) );
  AOI221_X1 dp_ex_stage_alu_U7 ( .B1(dp_ex_stage_muxA_out[31]), .B2(
        dp_ex_stage_alu_n204), .C1(dp_ex_stage_alu_n210), .C2(
        dp_ex_stage_alu_n249), .A(dp_ex_stage_alu_n199), .ZN(
        dp_ex_stage_alu_n117) );
  BUF_X2 dp_ex_stage_alu_U5 ( .A(dp_ex_stage_muxA_out[7]), .Z(
        dp_ex_stage_alu_n34) );
  MUX2_X1 dp_ex_stage_alu_U4 ( .A(dp_ex_stage_alu_n255), .B(
        dp_ex_stage_alu_N19), .S(dp_ex_stage_alu_n51), .Z(dp_ex_stage_alu_n256) );
  NAND3_X1 dp_ex_stage_alu_U235 ( .A1(dp_ex_stage_alu_n93), .A2(
        dp_ex_stage_alu_n270), .A3(dp_ex_stage_alu_n191), .ZN(
        dp_ex_stage_alu_n206) );
  NAND3_X1 dp_ex_stage_alu_U230 ( .A1(alu_op_i[4]), .A2(dp_ex_stage_alu_n54), 
        .A3(dp_ex_stage_alu_n67), .ZN(dp_ex_stage_alu_n91) );
  OR2_X1 dp_ex_stage_alu_adder_U53 ( .A1(dp_ex_stage_alu_n20), .A2(
        dp_ex_stage_alu_adder_n22), .ZN(dp_ex_stage_alu_adder_carries[0]) );
  XOR2_X1 dp_ex_stage_alu_adder_U52 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_muxB_out[5]), .Z(dp_ex_stage_alu_adder_n20) );
  XOR2_X1 dp_ex_stage_alu_adder_U51 ( .A(dp_ex_stage_alu_adder_n23), .B(
        dp_ex_stage_muxB_out[15]), .Z(dp_ex_stage_alu_adder_n18) );
  XOR2_X1 dp_ex_stage_alu_adder_U50 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_alu_n45), .Z(dp_ex_stage_alu_adder_n17) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U49 ( .A(dp_ex_stage_alu_adder_B_xor_3_), 
        .Z(dp_ex_stage_alu_adder_n16) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U48 ( .A(dp_ex_stage_alu_adder_n20), .Z(
        dp_ex_stage_alu_adder_n14) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U47 ( .A(dp_ex_stage_alu_adder_B_xor_6_), 
        .Z(dp_ex_stage_alu_adder_n10) );
  BUF_X2 dp_ex_stage_alu_adder_U46 ( .A(dp_ex_stage_alu_N23), .Z(
        dp_ex_stage_alu_adder_n15) );
  BUF_X1 dp_ex_stage_alu_adder_U45 ( .A(dp_ex_stage_alu_N23), .Z(
        dp_ex_stage_alu_adder_n21) );
  XOR2_X1 dp_ex_stage_alu_adder_U44 ( .A(dp_ex_stage_alu_adder_n13), .B(
        dp_ex_stage_muxB_out[23]), .Z(dp_ex_stage_alu_adder_B_xor_23_) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U43 ( .A(dp_ex_stage_alu_adder_B_xor_11_), 
        .Z(dp_ex_stage_alu_adder_n8) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U42 ( .A(dp_ex_stage_alu_adder_B_xor_13_), 
        .Z(dp_ex_stage_alu_adder_n7) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U41 ( .A(dp_ex_stage_alu_adder_n15), .Z(
        dp_ex_stage_alu_adder_n11) );
  XOR2_X1 dp_ex_stage_alu_adder_U40 ( .A(dp_ex_stage_alu_adder_n13), .B(
        dp_ex_stage_muxB_out[19]), .Z(dp_ex_stage_alu_adder_B_xor_19_) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U39 ( .A(dp_ex_stage_alu_adder_B_xor_19_), 
        .Z(dp_ex_stage_alu_adder_n6) );
  CLKBUF_X3 dp_ex_stage_alu_adder_U38 ( .A(dp_ex_stage_alu_N23), .Z(
        dp_ex_stage_alu_adder_n23) );
  XOR2_X1 dp_ex_stage_alu_adder_U37 ( .A(dp_ex_stage_alu_adder_n12), .B(
        dp_ex_stage_muxB_out[15]), .Z(dp_ex_stage_alu_adder_n5) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U36 ( .A(dp_ex_stage_alu_adder_B_xor_14_), 
        .Z(dp_ex_stage_alu_adder_n4) );
  XOR2_X1 dp_ex_stage_alu_adder_U35 ( .A(dp_ex_stage_alu_adder_n9), .B(
        dp_ex_stage_muxB_out[9]), .Z(dp_ex_stage_alu_adder_B_xor_9_) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U34 ( .A(dp_ex_stage_alu_adder_B_xor_9_), 
        .Z(dp_ex_stage_alu_adder_n3) );
  BUF_X2 dp_ex_stage_alu_adder_U30 ( .A(dp_ex_stage_alu_adder_n15), .Z(
        dp_ex_stage_alu_adder_n13) );
  CLKBUF_X3 dp_ex_stage_alu_adder_U27 ( .A(dp_ex_stage_alu_N23), .Z(
        dp_ex_stage_alu_adder_n22) );
  XOR2_X1 dp_ex_stage_alu_adder_U23 ( .A(dp_ex_stage_alu_adder_n21), .B(
        dp_ex_stage_muxB_out[7]), .Z(dp_ex_stage_alu_adder_n19) );
  CLKBUF_X1 dp_ex_stage_alu_adder_U18 ( .A(dp_ex_stage_alu_n231), .Z(
        dp_ex_stage_alu_adder_n2) );
  BUF_X1 dp_ex_stage_alu_adder_U6 ( .A(dp_ex_stage_alu_adder_n15), .Z(
        dp_ex_stage_alu_adder_n9) );
  XOR2_X1 dp_ex_stage_alu_adder_U4 ( .A(dp_ex_stage_alu_adder_n13), .B(
        dp_ex_stage_muxB_out[23]), .Z(dp_ex_stage_alu_adder_n1) );
  BUF_X2 dp_ex_stage_alu_adder_U2 ( .A(dp_ex_stage_alu_adder_n15), .Z(
        dp_ex_stage_alu_adder_n12) );
  XOR2_X2 dp_ex_stage_alu_adder_U1 ( .A(dp_ex_stage_alu_adder_n12), .B(
        dp_ex_stage_muxB_out[12]), .Z(dp_ex_stage_alu_adder_B_xor_12_) );
  XOR2_X1 dp_ex_stage_alu_adder_U33 ( .A(dp_ex_stage_alu_adder_n21), .B(
        dp_ex_stage_alu_n45), .Z(dp_ex_stage_alu_adder_B_xor_0_) );
  XOR2_X1 dp_ex_stage_alu_adder_U32 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_alu_n35), .Z(dp_ex_stage_alu_adder_B_xor_10_) );
  XOR2_X1 dp_ex_stage_alu_adder_U31 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_muxB_out[11]), .Z(dp_ex_stage_alu_adder_B_xor_11_) );
  XOR2_X1 dp_ex_stage_alu_adder_U29 ( .A(dp_ex_stage_alu_adder_n23), .B(
        dp_ex_stage_muxB_out[13]), .Z(dp_ex_stage_alu_adder_B_xor_13_) );
  XOR2_X1 dp_ex_stage_alu_adder_U28 ( .A(dp_ex_stage_alu_adder_n12), .B(
        dp_ex_stage_muxB_out[14]), .Z(dp_ex_stage_alu_adder_B_xor_14_) );
  XOR2_X1 dp_ex_stage_alu_adder_U26 ( .A(dp_ex_stage_alu_adder_n11), .B(
        dp_ex_stage_muxB_out[16]), .Z(dp_ex_stage_alu_adder_B_xor_16_) );
  XOR2_X1 dp_ex_stage_alu_adder_U25 ( .A(dp_ex_stage_alu_adder_n23), .B(
        dp_ex_stage_muxB_out[17]), .Z(dp_ex_stage_alu_adder_B_xor_17_) );
  XOR2_X1 dp_ex_stage_alu_adder_U24 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_muxB_out[18]), .Z(dp_ex_stage_alu_adder_B_xor_18_) );
  XOR2_X1 dp_ex_stage_alu_adder_U22 ( .A(dp_ex_stage_alu_adder_n21), .B(
        dp_ex_stage_alu_n46), .Z(dp_ex_stage_alu_adder_B_xor_1_) );
  XOR2_X1 dp_ex_stage_alu_adder_U21 ( .A(dp_ex_stage_alu_adder_n12), .B(
        dp_ex_stage_muxB_out[20]), .Z(dp_ex_stage_alu_adder_B_xor_20_) );
  XOR2_X1 dp_ex_stage_alu_adder_U20 ( .A(dp_ex_stage_alu_adder_n23), .B(
        dp_ex_stage_muxB_out[21]), .Z(dp_ex_stage_alu_adder_B_xor_21_) );
  XOR2_X1 dp_ex_stage_alu_adder_U19 ( .A(dp_ex_stage_alu_adder_n23), .B(
        dp_ex_stage_muxB_out[22]), .Z(dp_ex_stage_alu_adder_B_xor_22_) );
  XOR2_X1 dp_ex_stage_alu_adder_U17 ( .A(dp_ex_stage_alu_adder_n11), .B(
        dp_ex_stage_muxB_out[24]), .Z(dp_ex_stage_alu_adder_B_xor_24_) );
  XOR2_X1 dp_ex_stage_alu_adder_U16 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_muxB_out[25]), .Z(dp_ex_stage_alu_adder_B_xor_25_) );
  XOR2_X1 dp_ex_stage_alu_adder_U15 ( .A(dp_ex_stage_alu_adder_n23), .B(
        dp_ex_stage_muxB_out[26]), .Z(dp_ex_stage_alu_adder_B_xor_26_) );
  XOR2_X1 dp_ex_stage_alu_adder_U14 ( .A(dp_ex_stage_alu_adder_n23), .B(
        dp_ex_stage_muxB_out[27]), .Z(dp_ex_stage_alu_adder_B_xor_27_) );
  XOR2_X1 dp_ex_stage_alu_adder_U13 ( .A(dp_ex_stage_alu_adder_n23), .B(
        dp_ex_stage_muxB_out[28]), .Z(dp_ex_stage_alu_adder_B_xor_28_) );
  XOR2_X1 dp_ex_stage_alu_adder_U12 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_muxB_out[29]), .Z(dp_ex_stage_alu_adder_B_xor_29_) );
  XOR2_X1 dp_ex_stage_alu_adder_U11 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_alu_n50), .Z(dp_ex_stage_alu_adder_B_xor_2_) );
  XOR2_X1 dp_ex_stage_alu_adder_U10 ( .A(dp_ex_stage_alu_adder_n12), .B(
        dp_ex_stage_muxB_out[30]), .Z(dp_ex_stage_alu_adder_B_xor_30_) );
  XOR2_X1 dp_ex_stage_alu_adder_U9 ( .A(dp_ex_stage_alu_adder_n13), .B(
        dp_ex_stage_muxB_out[31]), .Z(dp_ex_stage_alu_adder_B_xor_31_) );
  XOR2_X1 dp_ex_stage_alu_adder_U8 ( .A(dp_ex_stage_alu_adder_n9), .B(
        dp_ex_stage_alu_n77), .Z(dp_ex_stage_alu_adder_B_xor_3_) );
  XOR2_X1 dp_ex_stage_alu_adder_U7 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_alu_n222), .Z(dp_ex_stage_alu_adder_B_xor_4_) );
  XOR2_X1 dp_ex_stage_alu_adder_U5 ( .A(dp_ex_stage_muxB_out[6]), .B(
        dp_ex_stage_alu_adder_n13), .Z(dp_ex_stage_alu_adder_B_xor_6_) );
  XOR2_X1 dp_ex_stage_alu_adder_U3 ( .A(dp_ex_stage_alu_adder_n22), .B(
        dp_ex_stage_muxB_out[8]), .Z(dp_ex_stage_alu_adder_B_xor_8_) );
  CLKBUF_X1 dp_ex_stage_alu_adder_SparseTree_U6 ( .A(
        dp_ex_stage_alu_adder_SparseTree_n1), .Z(
        dp_ex_stage_alu_adder_carries[2]) );
  CLKBUF_X1 dp_ex_stage_alu_adder_SparseTree_U5 ( .A(
        dp_ex_stage_alu_adder_SparseTree_gen_12__9_), .Z(
        dp_ex_stage_alu_adder_SparseTree_n4) );
  CLKBUF_X1 dp_ex_stage_alu_adder_SparseTree_U4 ( .A(
        dp_ex_stage_alu_adder_SparseTree_gen_24__17_), .Z(
        dp_ex_stage_alu_adder_SparseTree_n3) );
  CLKBUF_X1 dp_ex_stage_alu_adder_SparseTree_U3 ( .A(
        dp_ex_stage_alu_adder_SparseTree_n9), .Z(
        dp_ex_stage_alu_adder_carries[1]) );
  CLKBUF_X2 dp_ex_stage_alu_adder_SparseTree_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_n7), .Z(
        dp_ex_stage_alu_adder_carries[4]) );
  CLKBUF_X1 dp_ex_stage_alu_adder_SparseTree_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_n8), .Z(
        dp_ex_stage_alu_adder_SparseTree_n1) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_1_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_0_), .A2(dp_ex_stage_alu_shifter_N202), 
        .ZN(dp_ex_stage_alu_adder_SparseTree_gen_1__1_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_1_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_0_), .B(dp_ex_stage_alu_shifter_N202), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_1__1_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_2_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_1_), .A2(dp_ex_stage_alu_n76), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_2__2_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_2_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_1_), .B(dp_ex_stage_alu_n76), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_2__2_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_3_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_2_), .A2(dp_ex_stage_alu_n44), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_3__3_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_3_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_2_), .B(dp_ex_stage_alu_n44), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_3__3_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_4_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_3_), .A2(dp_ex_stage_alu_n69), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_4__4_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_4_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_3_), .B(dp_ex_stage_alu_n69), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_4__4_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_5_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_4_), .A2(dp_ex_stage_alu_n52), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_5__5_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_5_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_4_), .B(dp_ex_stage_alu_n52), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_5__5_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_6_U1 ( .A1(
        dp_ex_stage_alu_adder_n20), .A2(dp_ex_stage_muxA_out[5]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_6__6_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_6_U2 ( .A(
        dp_ex_stage_alu_adder_n20), .B(dp_ex_stage_muxA_out[5]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_6__6_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_7_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_6_), .A2(dp_ex_stage_alu_n78), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_7__7_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_7_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_6_), .B(dp_ex_stage_alu_n78), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_7__7_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_8_U1 ( .A1(
        dp_ex_stage_alu_adder_n19), .A2(dp_ex_stage_alu_n34), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_8__8_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_8_U2 ( .A(
        dp_ex_stage_alu_adder_n19), .B(dp_ex_stage_alu_n34), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_8__8_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_9_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_8_), .A2(dp_ex_stage_alu_n71), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_9__9_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_9_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_8_), .B(dp_ex_stage_alu_n71), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_9__9_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_10_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_9_), .A2(dp_ex_stage_alu_n72), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_10__10_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_10_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_9_), .B(dp_ex_stage_alu_n72), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_10__10_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_11_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_10_), .A2(dp_ex_stage_alu_n74), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_11__11_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_11_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_10_), .B(dp_ex_stage_alu_n74), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_11__11_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_12_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_11_), .A2(dp_ex_stage_muxA_out[11]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_12__12_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_12_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_11_), .B(dp_ex_stage_muxA_out[11]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_12__12_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_13_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_12_), .A2(dp_ex_stage_alu_n32), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_13__13_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_13_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_12_), .B(dp_ex_stage_alu_n32), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_13__13_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_14_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_13_), .A2(dp_ex_stage_alu_n231), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_14__14_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_14_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_13_), .B(dp_ex_stage_alu_n231), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_14__14_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_15_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_14_), .A2(dp_ex_stage_muxA_out[14]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_15__15_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_15_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_14_), .B(dp_ex_stage_muxA_out[14]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_15__15_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_16_U1 ( .A1(
        dp_ex_stage_alu_adder_n18), .A2(dp_ex_stage_alu_n29), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_16__16_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_16_U2 ( .A(
        dp_ex_stage_alu_adder_n18), .B(dp_ex_stage_alu_n29), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_16__16_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_17_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_16_), .A2(dp_ex_stage_alu_n38), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_17__17_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_17_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_16_), .B(dp_ex_stage_alu_n38), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_17__17_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_n1), .A2(
        dp_ex_stage_muxA_out[17]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_18__18_) );
  CLKBUF_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_U1 ( .A(
        dp_ex_stage_alu_adder_B_xor_17_), .Z(
        dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_n1) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_17_), .B(dp_ex_stage_muxA_out[17]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_18__18_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_19_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_18_), .A2(dp_ex_stage_muxA_out[18]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_19__19_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_19_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_18_), .B(dp_ex_stage_muxA_out[18]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_19__19_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_20_U1 ( .A1(
        dp_ex_stage_muxA_out[19]), .A2(dp_ex_stage_alu_adder_B_xor_19_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_20__20_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_20_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_19_), .B(dp_ex_stage_muxA_out[19]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_20__20_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_21_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_20_), .A2(dp_ex_stage_alu_n25), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_21__21_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_21_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_20_), .B(dp_ex_stage_alu_n25), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_21__21_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_n1), .A2(
        dp_ex_stage_alu_n238), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_22__22_) );
  CLKBUF_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_U1 ( .A(
        dp_ex_stage_alu_adder_B_xor_21_), .Z(
        dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_n1) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_21_), .B(dp_ex_stage_alu_n238), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_22__22_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_23_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_22_), .A2(dp_ex_stage_alu_n240), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_23__23_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_23_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_22_), .B(dp_ex_stage_alu_n240), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_23__23_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_24_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_23_), .A2(dp_ex_stage_muxA_out[23]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_24__24_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_24_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_23_), .B(dp_ex_stage_muxA_out[23]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_24__24_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_25_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_24_), .A2(dp_ex_stage_muxA_out[24]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_25__25_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_25_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_24_), .B(dp_ex_stage_muxA_out[24]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_25__25_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_26_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_25_), .A2(dp_ex_stage_muxA_out[25]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_26__26_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_26_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_25_), .B(dp_ex_stage_muxA_out[25]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_26__26_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_27_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_26_), .A2(dp_ex_stage_muxA_out[26]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_27__27_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_27_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_26_), .B(dp_ex_stage_muxA_out[26]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_27__27_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_28_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_27_), .A2(dp_ex_stage_muxA_out[27]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_28__28_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_28_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_27_), .B(dp_ex_stage_muxA_out[27]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_28__28_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_29_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_28_), .A2(dp_ex_stage_alu_n247), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_29__29_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_29_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_28_), .B(dp_ex_stage_alu_n247), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_29__29_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_30_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_29_), .A2(dp_ex_stage_muxA_out[29]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_30__30_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_30_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_29_), .B(dp_ex_stage_muxA_out[29]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_30__30_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_31_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_30_), .A2(dp_ex_stage_muxA_out[30]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_31__31_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_31_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_30_), .B(dp_ex_stage_muxA_out[30]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_31__31_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_32_U1 ( .A1(
        dp_ex_stage_alu_adder_B_xor_31_), .A2(dp_ex_stage_muxA_out[31]), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_32__32_) );
  XOR2_X1 dp_ex_stage_alu_adder_SparseTree_PG_net_i_32_U2 ( .A(
        dp_ex_stage_alu_adder_B_xor_31_), .B(dp_ex_stage_muxA_out[31]), .Z(
        dp_ex_stage_alu_adder_SparseTree_prop_32__32_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G10_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_1__1_), .B2(
        dp_ex_stage_alu_adder_carries[0]), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_1__1_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G10_n2) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G10_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G10_n2), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_1__0_) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G20_1_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G20_1_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_2__0_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G20_1_U1 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_1__0_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_2__2_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_2__2_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G20_1_n3) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_4__4_), .B2(
        dp_ex_stage_alu_adder_SparseTree_gen_3__3_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_4__4_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_n2) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_U2 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_3__3_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_4__4_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_4__3_) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_n2), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_4__3_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_5__5_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_6__6_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_6__5_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_5__5_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_6__6_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_6__6_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_6__5_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_8__8_), .B2(
        dp_ex_stage_alu_adder_SparseTree_gen_7__7_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_8__8_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_n3) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_U2 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_7__7_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_8__8_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_8__7_) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_8__7_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_10__10_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_9__9_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_10__9_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_10__10_), .B2(
        dp_ex_stage_alu_adder_SparseTree_gen_9__9_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_10__10_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_10__9_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_11__11_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_12__12_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_12__11_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_11__11_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_12__12_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_12__12_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_12__11_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_13__13_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_14__14_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_14__13_) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_14__13_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_U1 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_13__13_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_14__14_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_14__14_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_n3) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_16__16_), .B2(
        dp_ex_stage_alu_adder_SparseTree_gen_15__15_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_16__16_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_n3) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_U2 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_15__15_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_16__16_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_16__15_) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_16__15_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_18__18_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_17__17_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_18__17_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_17__17_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_18__18_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_18__18_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_18__17_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_19__19_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_20__20_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_20__19_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_20__20_), .B2(
        dp_ex_stage_alu_adder_SparseTree_gen_19__19_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_20__20_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_20__19_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_22__22_), .B2(
        dp_ex_stage_alu_adder_SparseTree_gen_21__21_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_22__22_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_22__21_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_U1 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_22__22_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_21__21_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_22__21_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_24__24_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_23__23_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_24__23_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_24__24_), .B2(
        dp_ex_stage_alu_adder_SparseTree_gen_23__23_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_24__24_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_24__23_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_25__25_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_26__26_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_26__25_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_25__25_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_26__26_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_26__26_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_26__25_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_27__27_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_28__28_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_28__27_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_27__27_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_28__28_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_28__28_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_28__27_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_29__29_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_30__30_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_30__30_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_30__29_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_U1 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_29__29_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_30__30_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_30__29_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_31__31_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_32__32_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_32__32_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_32__31_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_U1 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_31__31_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_32__32_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_32__31_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_2__0_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_4__3_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_4__3_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_n9) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_U3 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_8__5_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_6__5_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_8__7_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_8__7_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_n3) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_U1 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_6__5_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_8__7_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_8__5_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_10__9_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_12__11_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_12__9_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_10__9_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_12__11_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_12__11_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_12__9_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_14__13_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_16__15_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_16__13_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_14__13_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_16__15_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_16__15_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_16__13_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_18__17_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_20__19_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_20__17_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_18__17_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_20__19_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_20__19_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_20__17_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_22__21_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_24__23_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_24__21_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_22__21_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_24__23_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_24__23_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_24__21_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_26__25_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_28__27_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_28__25_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_26__25_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_28__27_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_28__27_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_28__25_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_30__29_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_32__31_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_32__31_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_32__29_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_U1 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_30__29_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_32__31_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_32__29_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_n9), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_8__5_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_8__5_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_n8) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_U3 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_16__9_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_12__9_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_16__13_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_16__13_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_n3) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_U1 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_12__9_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_16__13_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_16__9_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_U3 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_20__17_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_24__21_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_24__17_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_20__17_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_24__21_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_24__21_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_24__17_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_28__25_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_32__29_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_32__29_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_32__25_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_U1 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_28__25_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_32__29_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_32__25_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_n8), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_16__9_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_16__9_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_n7) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_12__9_), .B2(
        dp_ex_stage_alu_adder_SparseTree_n1), .A(
        dp_ex_stage_alu_adder_SparseTree_n4), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_n3), .ZN(
        dp_ex_stage_alu_adder_carries[3]) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_n3), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_32__25_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_32__25_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_n3) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_U2 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_24__17_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_32__25_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_32__17_) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_32__17_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_U3 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_gen_24__17_), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_28__25_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_28__25_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_gen_28__17_) );
  AND2_X1 dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_U1 ( .A1(
        dp_ex_stage_alu_adder_SparseTree_prop_24__17_), .A2(
        dp_ex_stage_alu_adder_SparseTree_prop_28__25_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_prop_28__17_) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_prop_32__17_), .B2(
        dp_ex_stage_alu_adder_carries[4]), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_32__17_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_n3), .ZN(
        dp_ex_stage_alu_adder_Cout) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_n7), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_28__17_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_28__17_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_n3), .ZN(
        dp_ex_stage_alu_adder_carries[7]) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_U2 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_n3), .ZN(
        dp_ex_stage_alu_adder_carries[6]) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_U1 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_n7), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_24__17_), .A(
        dp_ex_stage_alu_adder_SparseTree_n3), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_n3) );
  AOI21_X1 dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_U2 ( .B1(
        dp_ex_stage_alu_adder_SparseTree_n7), .B2(
        dp_ex_stage_alu_adder_SparseTree_prop_20__17_), .A(
        dp_ex_stage_alu_adder_SparseTree_gen_20__17_), .ZN(
        dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_n3) );
  INV_X1 dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_U1 ( .A(
        dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_n3), .ZN(
        dp_ex_stage_alu_adder_carries[5]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_alu_n69), .B(dp_ex_stage_alu_adder_n16), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_alu_n44), .B(dp_ex_stage_alu_adder_B_xor_2_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_alu_n76), .B(dp_ex_stage_alu_adder_B_xor_1_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_shifter_N202), .B(dp_ex_stage_alu_adder_n17), .CI(
        1'b0), .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0[0]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_alu_n69), .B(dp_ex_stage_alu_adder_n16), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_alu_n44), .B(dp_ex_stage_alu_adder_B_xor_2_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_alu_n76), .B(dp_ex_stage_alu_adder_B_xor_1_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_shifter_N202), .B(dp_ex_stage_alu_adder_n17), .CI(
        1'b1), .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1[0]) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U9 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0[0]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1[0]), .B2(
        dp_ex_stage_alu_adder_carries[0]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n9) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U8 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0[3]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5), .B1(
        dp_ex_stage_alu_adder_carries[0]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n6) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U7 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n6), .ZN(
        dp_ex_stage_alu_adder_out[3]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U6 ( .A(
        dp_ex_stage_alu_adder_carries[0]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U5 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0[1]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1[1]), .B2(
        dp_ex_stage_alu_adder_carries[0]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n8) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U4 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n8), .ZN(
        dp_ex_stage_alu_adder_out[1]) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U3 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0[2]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1[2]), .B2(
        dp_ex_stage_alu_adder_carries[0]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n7) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n7), .ZN(
        dp_ex_stage_alu_adder_out[2]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U1 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n9), .ZN(
        dp_ex_stage_alu_adder_out[0]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_alu_n34), .B(dp_ex_stage_alu_adder_n19), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_alu_n78), .B(dp_ex_stage_alu_adder_n10), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_muxA_out[5]), .B(dp_ex_stage_alu_adder_n14), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n52), .B(dp_ex_stage_alu_adder_B_xor_4_), .CI(1'b0), 
        .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0[0]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_alu_n34), .B(dp_ex_stage_alu_adder_n19), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_alu_n78), .B(dp_ex_stage_alu_adder_n10), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_muxA_out[5]), .B(dp_ex_stage_alu_adder_n14), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n52), .B(dp_ex_stage_alu_adder_B_xor_4_), .CI(1'b1), 
        .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1[0]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U9 ( .A(
        dp_ex_stage_alu_adder_carries[1]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U8 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0[0]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1[0]), .B2(
        dp_ex_stage_alu_adder_carries[1]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n10) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U7 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0[1]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1[1]), .B2(
        dp_ex_stage_alu_adder_carries[1]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n11) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U6 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0[2]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1[2]), .B2(
        dp_ex_stage_alu_adder_carries[1]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n12) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U5 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0[3]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5), .B1(
        dp_ex_stage_alu_adder_carries[1]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n13) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U4 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n10), .ZN(
        dp_ex_stage_alu_adder_out[4]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U3 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n11), .ZN(
        dp_ex_stage_alu_adder_out[5]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n12), .ZN(
        dp_ex_stage_alu_adder_out[6]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U1 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n13), .ZN(
        dp_ex_stage_alu_adder_out[7]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[11]), .B(dp_ex_stage_alu_adder_n8), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_alu_n74), .B(dp_ex_stage_alu_adder_B_xor_10_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_alu_n72), .B(dp_ex_stage_alu_adder_n3), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n71), .B(dp_ex_stage_alu_adder_B_xor_8_), .CI(1'b0), 
        .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0[0]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[11]), .B(dp_ex_stage_alu_adder_n8), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_alu_n74), .B(dp_ex_stage_alu_adder_B_xor_10_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_alu_n72), .B(dp_ex_stage_alu_adder_n3), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n71), .B(dp_ex_stage_alu_adder_B_xor_8_), .CI(1'b1), 
        .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1[0]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U9 ( .A(
        dp_ex_stage_alu_adder_carries[2]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U8 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0[1]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1[1]), .B2(
        dp_ex_stage_alu_adder_carries[2]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n11) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U7 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0[0]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1[0]), .B2(
        dp_ex_stage_alu_adder_carries[2]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n10) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U6 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0[2]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1[2]), .B2(
        dp_ex_stage_alu_adder_carries[2]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n12) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U5 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0[3]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5), .B1(
        dp_ex_stage_alu_adder_carries[2]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n13) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U4 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n10), .ZN(
        dp_ex_stage_alu_adder_out[8]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U3 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n13), .ZN(
        dp_ex_stage_alu_adder_out[11]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n11), .ZN(
        dp_ex_stage_alu_adder_out[9]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U1 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n12), .ZN(
        dp_ex_stage_alu_adder_out[10]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_alu_n29), .B(dp_ex_stage_alu_adder_n5), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_muxA_out[14]), .B(dp_ex_stage_alu_adder_n4), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_alu_adder_n2), .B(dp_ex_stage_alu_adder_n7), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n32), .B(dp_ex_stage_alu_adder_B_xor_12_), .CI(1'b0), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry[1]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0[0]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_alu_n29), .B(dp_ex_stage_alu_adder_n5), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_muxA_out[14]), .B(dp_ex_stage_alu_adder_n4), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_alu_adder_n2), .B(dp_ex_stage_alu_adder_n7), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n32), .B(dp_ex_stage_alu_adder_B_xor_12_), .CI(1'b1), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry[1]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1[0]) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U9 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0[3]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5), .B1(
        dp_ex_stage_alu_adder_carries[3]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n13) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U8 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0[0]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1[0]), .B2(
        dp_ex_stage_alu_adder_carries[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n10) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U7 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n10), .ZN(
        dp_ex_stage_alu_adder_out[12]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U6 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n13), .ZN(
        dp_ex_stage_alu_adder_out[15]) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U5 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0[1]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1[1]), .B2(
        dp_ex_stage_alu_adder_carries[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n11) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U4 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0[2]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1[2]), .B2(
        dp_ex_stage_alu_adder_carries[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n12) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U3 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n11), .ZN(
        dp_ex_stage_alu_adder_out[13]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n12), .ZN(
        dp_ex_stage_alu_adder_out[14]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U1 ( .A(
        dp_ex_stage_alu_adder_carries[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[19]), .B(dp_ex_stage_alu_adder_n6), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_muxA_out[18]), .B(dp_ex_stage_alu_adder_B_xor_18_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_muxA_out[17]), .B(dp_ex_stage_alu_adder_B_xor_17_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n38), .B(dp_ex_stage_alu_adder_B_xor_16_), .CI(1'b0), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry[1]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0[0]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[19]), .B(dp_ex_stage_alu_adder_n6), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_muxA_out[18]), .B(dp_ex_stage_alu_adder_B_xor_18_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_muxA_out[17]), .B(dp_ex_stage_alu_adder_B_xor_17_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n38), .B(dp_ex_stage_alu_adder_B_xor_16_), .CI(1'b1), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry[1]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1[0]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U9 ( .A(
        dp_ex_stage_alu_adder_carries[4]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U8 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0[0]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5), .B1(
        dp_ex_stage_alu_adder_carries[4]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1[0]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n10) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U7 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0[1]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1[1]), .B2(
        dp_ex_stage_alu_adder_carries[4]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n11) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U6 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0[2]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5), .B1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1[2]), .B2(
        dp_ex_stage_alu_adder_carries[4]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n12) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U5 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0[3]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5), .B1(
        dp_ex_stage_alu_adder_carries[4]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n13) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U4 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n10), .ZN(
        dp_ex_stage_alu_adder_out[16]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U3 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n11), .ZN(
        dp_ex_stage_alu_adder_out[17]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n12), .ZN(
        dp_ex_stage_alu_adder_out[18]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U1 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n13), .ZN(
        dp_ex_stage_alu_adder_out[19]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[23]), .B(dp_ex_stage_alu_adder_n1), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_alu_n240), .B(dp_ex_stage_alu_adder_B_xor_22_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_alu_n238), .B(dp_ex_stage_alu_adder_B_xor_21_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n25), .B(dp_ex_stage_alu_adder_B_xor_20_), .CI(1'b0), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry[1]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0[0]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[23]), .B(dp_ex_stage_alu_adder_n1), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_alu_n240), .B(dp_ex_stage_alu_adder_B_xor_22_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_alu_n238), .B(dp_ex_stage_alu_adder_B_xor_21_), .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n25), .B(dp_ex_stage_alu_adder_B_xor_20_), .CI(1'b1), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry[1]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1[0]) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U10 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n1), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0[0]), .B1(
        dp_ex_stage_alu_adder_carries[5]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1[0]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n11) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U9 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n11), .ZN(
        dp_ex_stage_alu_adder_out[20]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U8 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n14), .ZN(
        dp_ex_stage_alu_adder_out[23]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U7 ( .A(
        dp_ex_stage_alu_adder_carries[5]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n10) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U6 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0[3]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n10), .B1(
        dp_ex_stage_alu_adder_carries[5]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n14) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U5 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0[2]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n1), .B1(
        dp_ex_stage_alu_adder_carries[5]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1[2]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n13) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U4 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n10), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0[1]), .B1(
        dp_ex_stage_alu_adder_carries[5]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1[1]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n12) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U3 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n13), .ZN(
        dp_ex_stage_alu_adder_out[22]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n12), .ZN(
        dp_ex_stage_alu_adder_out[21]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U1 ( .A(
        dp_ex_stage_alu_adder_carries[5]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n1) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[27]), .B(dp_ex_stage_alu_adder_B_xor_27_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_muxA_out[26]), .B(dp_ex_stage_alu_adder_B_xor_26_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_muxA_out[25]), .B(dp_ex_stage_alu_adder_B_xor_25_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_muxA_out[24]), .B(dp_ex_stage_alu_adder_B_xor_24_), 
        .CI(1'b0), .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0[0]) );
  NAND3_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U6 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n2), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n3), .A3(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n4), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_3_) );
  NAND2_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U5 ( .A1(
        dp_ex_stage_alu_adder_B_xor_26_), .A2(dp_ex_stage_muxA_out[26]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n4) );
  NAND2_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U4 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_), .A2(dp_ex_stage_muxA_out[26]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n3) );
  NAND2_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U3 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_), .A2(dp_ex_stage_alu_adder_B_xor_26_), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n2) );
  XOR2_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_), .B(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n1), .Z(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1[2]) );
  XOR2_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U1 ( .A(
        dp_ex_stage_alu_adder_B_xor_26_), .B(dp_ex_stage_muxA_out[26]), .Z(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n1) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[27]), .B(dp_ex_stage_alu_adder_B_xor_27_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_3_), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_muxA_out[25]), .B(dp_ex_stage_alu_adder_B_xor_25_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_1_), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_muxA_out[24]), .B(dp_ex_stage_alu_adder_B_xor_24_), 
        .CI(1'b1), .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_1_), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1[0]) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U10 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n1), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0[3]), .B1(
        dp_ex_stage_alu_adder_carries[6]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n14) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U9 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0[2]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n1), .B1(
        dp_ex_stage_alu_adder_carries[6]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1[2]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n13) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U8 ( .A(
        dp_ex_stage_alu_adder_carries[6]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n10) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U7 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0[1]), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n10), .B1(
        dp_ex_stage_alu_adder_carries[6]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1[1]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n12) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U6 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n10), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0[0]), .B1(
        dp_ex_stage_alu_adder_carries[6]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1[0]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n11) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U5 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n13), .ZN(
        dp_ex_stage_alu_adder_out[26]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U4 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n11), .ZN(
        dp_ex_stage_alu_adder_out[24]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U3 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n14), .ZN(
        dp_ex_stage_alu_adder_out[27]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n12), .ZN(
        dp_ex_stage_alu_adder_out[25]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U1 ( .A(
        dp_ex_stage_alu_adder_carries[6]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n1) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[31]), .B(dp_ex_stage_alu_adder_B_xor_31_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_muxA_out[30]), .B(dp_ex_stage_alu_adder_B_xor_30_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_muxA_out[29]), .B(dp_ex_stage_alu_adder_B_xor_29_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n247), .B(dp_ex_stage_alu_adder_B_xor_28_), .CI(
        1'b0), .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0[0]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_U1_3 ( 
        .A(dp_ex_stage_muxA_out[31]), .B(dp_ex_stage_alu_adder_B_xor_31_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry[3]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_Co), .S(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1[3]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_U1_2 ( 
        .A(dp_ex_stage_muxA_out[30]), .B(dp_ex_stage_alu_adder_B_xor_30_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry[2]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry[3]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1[2]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_U1_1 ( 
        .A(dp_ex_stage_muxA_out[29]), .B(dp_ex_stage_alu_adder_B_xor_29_), 
        .CI(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry[1]), .CO(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry[2]), 
        .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1[1]) );
  FA_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_U1_0 ( 
        .A(dp_ex_stage_alu_n247), .B(dp_ex_stage_alu_adder_B_xor_28_), .CI(
        1'b1), .CO(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry[1]), .S(dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1[0]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U10 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n14), .ZN(
        dp_ex_stage_alu_adder_out[31]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U9 ( .A(
        dp_ex_stage_alu_adder_carries[7]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n10) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U8 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n1), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0[3]), .B1(
        dp_ex_stage_alu_adder_carries[7]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1[3]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n14) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U7 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n10), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0[0]), .B1(
        dp_ex_stage_alu_adder_carries[7]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1[0]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n11) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U6 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n10), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0[1]), .B1(
        dp_ex_stage_alu_adder_carries[7]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1[1]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n12) );
  AOI22_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U5 ( .A1(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n1), .A2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0[2]), .B1(
        dp_ex_stage_alu_adder_carries[7]), .B2(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1[2]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n13) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U4 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n12), .ZN(
        dp_ex_stage_alu_adder_out[29]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U3 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n11), .ZN(
        dp_ex_stage_alu_adder_out[28]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U2 ( .A(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n13), .ZN(
        dp_ex_stage_alu_adder_out[30]) );
  INV_X1 dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U1 ( .A(
        dp_ex_stage_alu_adder_carries[7]), .ZN(
        dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n1) );
  AOI222_X1 dp_ex_stage_alu_shifter_U150 ( .A1(dp_ex_stage_alu_shifter_N207), 
        .A2(dp_ex_stage_alu_shifter_n115), .B1(dp_ex_stage_alu_shifter_N110), 
        .B2(dp_ex_stage_alu_shifter_n112), .C1(dp_ex_stage_alu_shifter_N142), 
        .C2(dp_ex_stage_alu_shifter_n109), .ZN(dp_ex_stage_alu_shifter_n36) );
  NAND2_X1 dp_ex_stage_alu_shifter_U149 ( .A1(dp_ex_stage_alu_shifter_n33), 
        .A2(dp_ex_stage_alu_shifter_n34), .ZN(dp_ex_stage_alu_shifter_out[6])
         );
  NAND2_X1 dp_ex_stage_alu_shifter_U148 ( .A1(dp_ex_stage_alu_shifter_n37), 
        .A2(dp_ex_stage_alu_shifter_n38), .ZN(dp_ex_stage_alu_shifter_out[4])
         );
  NAND2_X1 dp_ex_stage_alu_shifter_U147 ( .A1(dp_ex_stage_alu_shifter_n35), 
        .A2(dp_ex_stage_alu_shifter_n36), .ZN(dp_ex_stage_alu_shifter_out[5])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U146 ( .A1(dp_ex_stage_alu_shifter_N213), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N116), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N148), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n86) );
  AOI222_X1 dp_ex_stage_alu_shifter_U145 ( .A1(dp_ex_stage_alu_shifter_N208), 
        .A2(dp_ex_stage_alu_shifter_n115), .B1(dp_ex_stage_alu_shifter_N111), 
        .B2(dp_ex_stage_alu_shifter_n112), .C1(dp_ex_stage_alu_shifter_N143), 
        .C2(dp_ex_stage_alu_shifter_n109), .ZN(dp_ex_stage_alu_shifter_n34) );
  AOI222_X1 dp_ex_stage_alu_shifter_U144 ( .A1(dp_ex_stage_alu_shifter_N206), 
        .A2(dp_ex_stage_alu_shifter_n115), .B1(dp_ex_stage_alu_shifter_N109), 
        .B2(dp_ex_stage_alu_shifter_n112), .C1(dp_ex_stage_alu_shifter_N141), 
        .C2(dp_ex_stage_alu_shifter_n109), .ZN(dp_ex_stage_alu_shifter_n38) );
  AOI222_X1 dp_ex_stage_alu_shifter_U143 ( .A1(dp_ex_stage_alu_shifter_N205), 
        .A2(dp_ex_stage_alu_shifter_n115), .B1(dp_ex_stage_alu_shifter_N108), 
        .B2(dp_ex_stage_alu_shifter_n112), .C1(dp_ex_stage_alu_shifter_N140), 
        .C2(dp_ex_stage_alu_shifter_n109), .ZN(dp_ex_stage_alu_shifter_n40) );
  NAND2_X1 dp_ex_stage_alu_shifter_U142 ( .A1(dp_ex_stage_alu_shifter_n39), 
        .A2(dp_ex_stage_alu_shifter_n40), .ZN(dp_ex_stage_alu_shifter_out[3])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U141 ( .A1(dp_ex_stage_alu_shifter_N219), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N122), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N154), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n74) );
  NAND2_X1 dp_ex_stage_alu_shifter_U140 ( .A1(dp_ex_stage_alu_shifter_n73), 
        .A2(dp_ex_stage_alu_shifter_n74), .ZN(dp_ex_stage_alu_shifter_out[17])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U139 ( .A1(dp_ex_stage_alu_shifter_N203), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N106), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N138), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n68) );
  NAND2_X1 dp_ex_stage_alu_shifter_U138 ( .A1(dp_ex_stage_alu_shifter_n67), 
        .A2(dp_ex_stage_alu_shifter_n68), .ZN(dp_ex_stage_alu_shifter_out[1])
         );
  NAND2_X1 dp_ex_stage_alu_shifter_U137 ( .A1(dp_ex_stage_alu_shifter_n90), 
        .A2(dp_ex_stage_alu_shifter_n89), .ZN(dp_ex_stage_alu_shifter_out[0])
         );
  NAND2_X1 dp_ex_stage_alu_shifter_U136 ( .A1(dp_ex_stage_alu_shifter_n45), 
        .A2(dp_ex_stage_alu_shifter_n46), .ZN(dp_ex_stage_alu_shifter_out[2])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U135 ( .A1(dp_ex_stage_alu_shifter_N218), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N121), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N153), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n76) );
  NAND2_X1 dp_ex_stage_alu_shifter_U134 ( .A1(dp_ex_stage_alu_shifter_n75), 
        .A2(dp_ex_stage_alu_shifter_n76), .ZN(dp_ex_stage_alu_shifter_out[16])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U133 ( .A1(dp_ex_stage_alu_shifter_N221), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N124), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N156), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n70) );
  NAND2_X1 dp_ex_stage_alu_shifter_U132 ( .A1(dp_ex_stage_alu_shifter_n69), 
        .A2(dp_ex_stage_alu_shifter_n70), .ZN(dp_ex_stage_alu_shifter_out[19])
         );
  NAND2_X1 dp_ex_stage_alu_shifter_U131 ( .A1(dp_ex_stage_alu_shifter_n83), 
        .A2(dp_ex_stage_alu_shifter_n84), .ZN(dp_ex_stage_alu_shifter_out[12])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U130 ( .A1(dp_ex_stage_alu_shifter_N212), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N115), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N147), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n88) );
  NAND2_X1 dp_ex_stage_alu_shifter_U129 ( .A1(dp_ex_stage_alu_shifter_n87), 
        .A2(dp_ex_stage_alu_shifter_n88), .ZN(dp_ex_stage_alu_shifter_out[10])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U128 ( .A1(dp_ex_stage_alu_shifter_N210), 
        .A2(dp_ex_stage_alu_shifter_n115), .B1(dp_ex_stage_alu_shifter_N113), 
        .B2(dp_ex_stage_alu_shifter_n112), .C1(dp_ex_stage_alu_shifter_N145), 
        .C2(dp_ex_stage_alu_shifter_n109), .ZN(dp_ex_stage_alu_shifter_n30) );
  NAND2_X1 dp_ex_stage_alu_shifter_U127 ( .A1(dp_ex_stage_alu_shifter_n29), 
        .A2(dp_ex_stage_alu_shifter_n30), .ZN(dp_ex_stage_alu_shifter_out[8])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U126 ( .A1(dp_ex_stage_alu_shifter_N211), 
        .A2(dp_ex_stage_alu_shifter_n115), .B1(dp_ex_stage_alu_shifter_N114), 
        .B2(dp_ex_stage_alu_shifter_n112), .C1(dp_ex_stage_alu_shifter_N146), 
        .C2(dp_ex_stage_alu_shifter_n109), .ZN(dp_ex_stage_alu_shifter_n22) );
  NAND2_X1 dp_ex_stage_alu_shifter_U125 ( .A1(dp_ex_stage_alu_shifter_n21), 
        .A2(dp_ex_stage_alu_shifter_n22), .ZN(dp_ex_stage_alu_shifter_out[9])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U124 ( .A1(dp_ex_stage_alu_shifter_N220), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N123), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N155), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n72) );
  NAND2_X1 dp_ex_stage_alu_shifter_U123 ( .A1(dp_ex_stage_alu_shifter_n71), 
        .A2(dp_ex_stage_alu_shifter_n72), .ZN(dp_ex_stage_alu_shifter_out[18])
         );
  NOR2_X1 dp_ex_stage_alu_shifter_U122 ( .A1(dp_ex_stage_alu_n208), .A2(1'b1), 
        .ZN(dp_ex_stage_alu_shifter_n28) );
  NOR2_X1 dp_ex_stage_alu_shifter_U121 ( .A1(dp_ex_stage_alu_shifter_n118), 
        .A2(1'b1), .ZN(dp_ex_stage_alu_shifter_n26) );
  AND2_X1 dp_ex_stage_alu_shifter_U120 ( .A1(dp_ex_stage_alu_shift_arith_i), 
        .A2(1'b1), .ZN(dp_ex_stage_alu_shifter_n91) );
  INV_X1 dp_ex_stage_alu_shifter_U119 ( .A(1'b1), .ZN(
        dp_ex_stage_alu_shifter_n117) );
  NOR2_X1 dp_ex_stage_alu_shifter_U118 ( .A1(dp_ex_stage_alu_shifter_n117), 
        .A2(dp_ex_stage_alu_shift_arith_i), .ZN(dp_ex_stage_alu_shifter_n92)
         );
  BUF_X1 dp_ex_stage_alu_shifter_U117 ( .A(dp_ex_stage_alu_shifter_n26), .Z(
        dp_ex_stage_alu_shifter_n106) );
  BUF_X1 dp_ex_stage_alu_shifter_U116 ( .A(dp_ex_stage_alu_shifter_n28), .Z(
        dp_ex_stage_alu_shifter_n100) );
  BUF_X1 dp_ex_stage_alu_shifter_U115 ( .A(dp_ex_stage_alu_shifter_n26), .Z(
        dp_ex_stage_alu_shifter_n104) );
  BUF_X1 dp_ex_stage_alu_shifter_U114 ( .A(dp_ex_stage_alu_shifter_n26), .Z(
        dp_ex_stage_alu_shifter_n105) );
  BUF_X1 dp_ex_stage_alu_shifter_U113 ( .A(dp_ex_stage_alu_shifter_n28), .Z(
        dp_ex_stage_alu_shifter_n98) );
  BUF_X1 dp_ex_stage_alu_shifter_U112 ( .A(dp_ex_stage_alu_shifter_n28), .Z(
        dp_ex_stage_alu_shifter_n99) );
  AND2_X1 dp_ex_stage_alu_shifter_U111 ( .A1(dp_ex_stage_alu_shifter_n91), 
        .A2(dp_ex_stage_alu_shifter_n118), .ZN(dp_ex_stage_alu_shifter_n25) );
  AND2_X1 dp_ex_stage_alu_shifter_U110 ( .A1(dp_ex_stage_alu_shifter_n92), 
        .A2(dp_ex_stage_alu_shifter_n118), .ZN(dp_ex_stage_alu_shifter_n24) );
  AND2_X1 dp_ex_stage_alu_shifter_U109 ( .A1(dp_ex_stage_alu_n208), .A2(
        dp_ex_stage_alu_shifter_n91), .ZN(dp_ex_stage_alu_shifter_n27) );
  AND2_X1 dp_ex_stage_alu_shifter_U108 ( .A1(dp_ex_stage_alu_n208), .A2(
        dp_ex_stage_alu_shifter_n92), .ZN(dp_ex_stage_alu_shifter_n23) );
  AOI222_X1 dp_ex_stage_alu_shifter_U107 ( .A1(dp_ex_stage_alu_shifter_N229), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N132), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N164), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n52) );
  AOI222_X1 dp_ex_stage_alu_shifter_U106 ( .A1(dp_ex_stage_alu_shifter_N54), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N249), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N22), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n77) );
  NAND2_X1 dp_ex_stage_alu_shifter_U105 ( .A1(dp_ex_stage_alu_shifter_n77), 
        .A2(dp_ex_stage_alu_shifter_n78), .ZN(dp_ex_stage_alu_shifter_out[15])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U104 ( .A1(dp_ex_stage_alu_shifter_N59), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N254), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N27), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n65) );
  NAND2_X1 dp_ex_stage_alu_shifter_U103 ( .A1(dp_ex_stage_alu_shifter_n65), 
        .A2(dp_ex_stage_alu_shifter_n66), .ZN(dp_ex_stage_alu_shifter_out[20])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U102 ( .A1(dp_ex_stage_alu_shifter_N62), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N257), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N30), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n59) );
  NAND2_X1 dp_ex_stage_alu_shifter_U101 ( .A1(dp_ex_stage_alu_shifter_n59), 
        .A2(dp_ex_stage_alu_shifter_n60), .ZN(dp_ex_stage_alu_shifter_out[23])
         );
  INV_X1 dp_ex_stage_alu_shifter_U100 ( .A(dp_ex_stage_alu_n208), .ZN(
        dp_ex_stage_alu_shifter_n118) );
  NAND2_X1 dp_ex_stage_alu_shifter_U99 ( .A1(dp_ex_stage_alu_shifter_n85), 
        .A2(dp_ex_stage_alu_shifter_n86), .ZN(dp_ex_stage_alu_shifter_out[11])
         );
  BUF_X1 dp_ex_stage_alu_shifter_U98 ( .A(dp_ex_stage_alu_shifter_n25), .Z(
        dp_ex_stage_alu_shifter_n109) );
  BUF_X1 dp_ex_stage_alu_shifter_U97 ( .A(dp_ex_stage_alu_shifter_n24), .Z(
        dp_ex_stage_alu_shifter_n112) );
  BUF_X1 dp_ex_stage_alu_shifter_U96 ( .A(dp_ex_stage_alu_shifter_n23), .Z(
        dp_ex_stage_alu_shifter_n115) );
  BUF_X1 dp_ex_stage_alu_shifter_U95 ( .A(dp_ex_stage_alu_shifter_n23), .Z(
        dp_ex_stage_alu_shifter_n113) );
  CLKBUF_X3 dp_ex_stage_alu_shifter_U94 ( .A(dp_ex_stage_muxB_out[4]), .Z(
        dp_ex_stage_alu_shifter_n116) );
  AOI222_X1 dp_ex_stage_alu_shifter_U93 ( .A1(dp_ex_stage_alu_shifter_N69), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N264), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N37), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n43) );
  NAND2_X1 dp_ex_stage_alu_shifter_U92 ( .A1(dp_ex_stage_alu_shifter_n43), 
        .A2(dp_ex_stage_alu_shifter_n44), .ZN(dp_ex_stage_alu_shifter_out[30])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U91 ( .A1(dp_ex_stage_alu_shifter_N70), 
        .A2(dp_ex_stage_alu_shifter_n106), .B1(dp_ex_stage_alu_shifter_N265), 
        .B2(dp_ex_stage_alu_shifter_n103), .C1(dp_ex_stage_alu_shifter_N38), 
        .C2(dp_ex_stage_alu_shifter_n100), .ZN(dp_ex_stage_alu_shifter_n41) );
  NAND2_X1 dp_ex_stage_alu_shifter_U90 ( .A1(dp_ex_stage_alu_shifter_n41), 
        .A2(dp_ex_stage_alu_shifter_n42), .ZN(dp_ex_stage_alu_shifter_out[31])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U89 ( .A1(dp_ex_stage_alu_shifter_N67), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N262), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N35), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n49) );
  NAND2_X1 dp_ex_stage_alu_shifter_U88 ( .A1(dp_ex_stage_alu_shifter_n49), 
        .A2(dp_ex_stage_alu_shifter_n50), .ZN(dp_ex_stage_alu_shifter_out[28])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U87 ( .A1(dp_ex_stage_alu_shifter_N68), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N263), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N36), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n47) );
  NAND2_X1 dp_ex_stage_alu_shifter_U86 ( .A1(dp_ex_stage_alu_shifter_n47), 
        .A2(dp_ex_stage_alu_shifter_n48), .ZN(dp_ex_stage_alu_shifter_out[29])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U85 ( .A1(dp_ex_stage_alu_shifter_N63), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N258), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N31), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n57) );
  NAND2_X1 dp_ex_stage_alu_shifter_U84 ( .A1(dp_ex_stage_alu_shifter_n57), 
        .A2(dp_ex_stage_alu_shifter_n58), .ZN(dp_ex_stage_alu_shifter_out[24])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U83 ( .A1(dp_ex_stage_alu_shifter_N61), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N256), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N29), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n61) );
  NAND2_X1 dp_ex_stage_alu_shifter_U82 ( .A1(dp_ex_stage_alu_shifter_n61), 
        .A2(dp_ex_stage_alu_shifter_n62), .ZN(dp_ex_stage_alu_shifter_out[22])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U81 ( .A1(dp_ex_stage_alu_shifter_N65), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N260), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N33), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n53) );
  NAND2_X1 dp_ex_stage_alu_shifter_U80 ( .A1(dp_ex_stage_alu_shifter_n53), 
        .A2(dp_ex_stage_alu_shifter_n54), .ZN(dp_ex_stage_alu_shifter_out[26])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U79 ( .A1(dp_ex_stage_alu_shifter_N64), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N259), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N32), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n55) );
  NAND2_X1 dp_ex_stage_alu_shifter_U78 ( .A1(dp_ex_stage_alu_shifter_n55), 
        .A2(dp_ex_stage_alu_shifter_n56), .ZN(dp_ex_stage_alu_shifter_out[25])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U77 ( .A1(dp_ex_stage_alu_shifter_N60), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N255), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N28), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n63) );
  NAND2_X1 dp_ex_stage_alu_shifter_U76 ( .A1(dp_ex_stage_alu_shifter_n63), 
        .A2(dp_ex_stage_alu_shifter_n64), .ZN(dp_ex_stage_alu_shifter_out[21])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U75 ( .A1(dp_ex_stage_alu_shifter_N66), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N261), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N34), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n51) );
  NAND2_X1 dp_ex_stage_alu_shifter_U74 ( .A1(dp_ex_stage_alu_shifter_n51), 
        .A2(dp_ex_stage_alu_shifter_n52), .ZN(dp_ex_stage_alu_shifter_out[27])
         );
  NAND2_X1 dp_ex_stage_alu_shifter_U73 ( .A1(dp_ex_stage_alu_shifter_n31), 
        .A2(dp_ex_stage_alu_shifter_n32), .ZN(dp_ex_stage_alu_shifter_out[7])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U72 ( .A1(dp_ex_stage_alu_shifter_N52), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N247), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N20), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n81) );
  NAND2_X1 dp_ex_stage_alu_shifter_U71 ( .A1(dp_ex_stage_alu_shifter_n81), 
        .A2(dp_ex_stage_alu_shifter_n82), .ZN(dp_ex_stage_alu_shifter_out[13])
         );
  AOI222_X1 dp_ex_stage_alu_shifter_U70 ( .A1(dp_ex_stage_alu_shifter_N53), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N248), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N21), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n79) );
  NAND2_X1 dp_ex_stage_alu_shifter_U69 ( .A1(dp_ex_stage_alu_shifter_n79), 
        .A2(dp_ex_stage_alu_shifter_n80), .ZN(dp_ex_stage_alu_shifter_out[14])
         );
  BUF_X1 dp_ex_stage_alu_shifter_U68 ( .A(dp_ex_stage_alu_shifter_n27), .Z(
        dp_ex_stage_alu_shifter_n103) );
  BUF_X1 dp_ex_stage_alu_shifter_U67 ( .A(dp_ex_stage_alu_shifter_n23), .Z(
        dp_ex_stage_alu_shifter_n114) );
  BUF_X1 dp_ex_stage_alu_shifter_U66 ( .A(dp_ex_stage_alu_shifter_n24), .Z(
        dp_ex_stage_alu_shifter_n111) );
  BUF_X1 dp_ex_stage_alu_shifter_U65 ( .A(dp_ex_stage_alu_shifter_n27), .Z(
        dp_ex_stage_alu_shifter_n101) );
  BUF_X1 dp_ex_stage_alu_shifter_U64 ( .A(dp_ex_stage_alu_shifter_n27), .Z(
        dp_ex_stage_alu_shifter_n102) );
  AOI222_X1 dp_ex_stage_alu_shifter_U63 ( .A1(dp_ex_stage_alu_shifter_N51), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N246), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N19), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n83) );
  AOI222_X1 dp_ex_stage_alu_shifter_U62 ( .A1(dp_ex_stage_alu_shifter_N49), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N244), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N17), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n87) );
  AOI222_X1 dp_ex_stage_alu_shifter_U61 ( .A1(dp_ex_stage_alu_shifter_N56), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N251), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N24), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n73) );
  AOI222_X1 dp_ex_stage_alu_shifter_U60 ( .A1(dp_ex_stage_alu_shifter_N57), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N252), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N25), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n71) );
  AOI222_X1 dp_ex_stage_alu_shifter_U59 ( .A1(dp_ex_stage_alu_shifter_N58), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N253), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N26), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n69) );
  AOI222_X1 dp_ex_stage_alu_shifter_U58 ( .A1(dp_ex_stage_alu_shifter_N55), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N250), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N23), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n75) );
  AOI222_X1 dp_ex_stage_alu_shifter_U57 ( .A1(dp_ex_stage_alu_shifter_N39), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N234), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N7), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n89) );
  AOI222_X1 dp_ex_stage_alu_shifter_U56 ( .A1(dp_ex_stage_alu_shifter_N40), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N235), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N8), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n67) );
  AOI222_X1 dp_ex_stage_alu_shifter_U55 ( .A1(dp_ex_stage_alu_shifter_N41), 
        .A2(dp_ex_stage_alu_shifter_n105), .B1(dp_ex_stage_alu_shifter_N236), 
        .B2(dp_ex_stage_alu_shifter_n102), .C1(dp_ex_stage_alu_shifter_N9), 
        .C2(dp_ex_stage_alu_shifter_n99), .ZN(dp_ex_stage_alu_shifter_n45) );
  AOI222_X1 dp_ex_stage_alu_shifter_U54 ( .A1(dp_ex_stage_alu_shifter_N45), 
        .A2(dp_ex_stage_alu_shifter_n106), .B1(dp_ex_stage_alu_shifter_N240), 
        .B2(dp_ex_stage_alu_shifter_n103), .C1(dp_ex_stage_alu_shifter_N13), 
        .C2(dp_ex_stage_alu_shifter_n100), .ZN(dp_ex_stage_alu_shifter_n33) );
  AOI222_X1 dp_ex_stage_alu_shifter_U53 ( .A1(dp_ex_stage_alu_shifter_N48), 
        .A2(dp_ex_stage_alu_shifter_n106), .B1(dp_ex_stage_alu_shifter_N243), 
        .B2(dp_ex_stage_alu_shifter_n103), .C1(dp_ex_stage_alu_shifter_N16), 
        .C2(dp_ex_stage_alu_shifter_n100), .ZN(dp_ex_stage_alu_shifter_n21) );
  AOI222_X1 dp_ex_stage_alu_shifter_U52 ( .A1(dp_ex_stage_alu_shifter_N47), 
        .A2(dp_ex_stage_alu_shifter_n106), .B1(dp_ex_stage_alu_shifter_N242), 
        .B2(dp_ex_stage_alu_shifter_n103), .C1(dp_ex_stage_alu_shifter_N15), 
        .C2(dp_ex_stage_alu_shifter_n100), .ZN(dp_ex_stage_alu_shifter_n29) );
  AOI222_X1 dp_ex_stage_alu_shifter_U51 ( .A1(dp_ex_stage_alu_shifter_N42), 
        .A2(dp_ex_stage_alu_shifter_n106), .B1(dp_ex_stage_alu_shifter_N237), 
        .B2(dp_ex_stage_alu_shifter_n103), .C1(dp_ex_stage_alu_shifter_N10), 
        .C2(dp_ex_stage_alu_shifter_n100), .ZN(dp_ex_stage_alu_shifter_n39) );
  AOI222_X1 dp_ex_stage_alu_shifter_U50 ( .A1(dp_ex_stage_alu_shifter_N43), 
        .A2(dp_ex_stage_alu_shifter_n106), .B1(dp_ex_stage_alu_shifter_N238), 
        .B2(dp_ex_stage_alu_shifter_n103), .C1(dp_ex_stage_alu_shifter_N11), 
        .C2(dp_ex_stage_alu_shifter_n100), .ZN(dp_ex_stage_alu_shifter_n37) );
  AOI222_X1 dp_ex_stage_alu_shifter_U49 ( .A1(dp_ex_stage_alu_shifter_N44), 
        .A2(dp_ex_stage_alu_shifter_n106), .B1(dp_ex_stage_alu_shifter_N239), 
        .B2(dp_ex_stage_alu_shifter_n103), .C1(dp_ex_stage_alu_shifter_N12), 
        .C2(dp_ex_stage_alu_shifter_n100), .ZN(dp_ex_stage_alu_shifter_n35) );
  AOI222_X1 dp_ex_stage_alu_shifter_U48 ( .A1(dp_ex_stage_alu_shifter_N50), 
        .A2(dp_ex_stage_alu_shifter_n104), .B1(dp_ex_stage_alu_shifter_N245), 
        .B2(dp_ex_stage_alu_shifter_n101), .C1(dp_ex_stage_alu_shifter_N18), 
        .C2(dp_ex_stage_alu_shifter_n98), .ZN(dp_ex_stage_alu_shifter_n85) );
  AOI222_X1 dp_ex_stage_alu_shifter_U47 ( .A1(dp_ex_stage_alu_shifter_N46), 
        .A2(dp_ex_stage_alu_shifter_n106), .B1(dp_ex_stage_alu_shifter_N241), 
        .B2(dp_ex_stage_alu_shifter_n103), .C1(dp_ex_stage_alu_shifter_N14), 
        .C2(dp_ex_stage_alu_shifter_n100), .ZN(dp_ex_stage_alu_shifter_n31) );
  AOI222_X1 dp_ex_stage_alu_shifter_U46 ( .A1(dp_ex_stage_alu_shifter_N217), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N120), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N152), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n78) );
  AOI222_X1 dp_ex_stage_alu_shifter_U45 ( .A1(dp_ex_stage_alu_shifter_N215), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N118), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N150), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n82) );
  AOI222_X1 dp_ex_stage_alu_shifter_U44 ( .A1(dp_ex_stage_alu_shifter_N216), 
        .A2(dp_ex_stage_alu_shifter_n113), .B1(dp_ex_stage_alu_shifter_N119), 
        .B2(dp_ex_stage_alu_shifter_n110), .C1(dp_ex_stage_alu_shifter_N151), 
        .C2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n80) );
  AOI222_X1 dp_ex_stage_alu_shifter_U43 ( .A1(dp_ex_stage_alu_shifter_N230), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N133), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N165), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n50) );
  AOI222_X1 dp_ex_stage_alu_shifter_U42 ( .A1(dp_ex_stage_alu_shifter_N232), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N135), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N167), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n44) );
  AOI222_X1 dp_ex_stage_alu_shifter_U41 ( .A1(dp_ex_stage_alu_shifter_N231), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N134), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N166), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n48) );
  AOI222_X1 dp_ex_stage_alu_shifter_U40 ( .A1(dp_ex_stage_alu_shifter_N233), 
        .A2(dp_ex_stage_alu_shifter_n115), .B1(dp_ex_stage_alu_shifter_N136), 
        .B2(dp_ex_stage_alu_shifter_n112), .C1(dp_ex_stage_alu_shifter_N168), 
        .C2(dp_ex_stage_alu_shifter_n109), .ZN(dp_ex_stage_alu_shifter_n42) );
  AOI222_X1 dp_ex_stage_alu_shifter_U39 ( .A1(dp_ex_stage_alu_shifter_N209), 
        .A2(dp_ex_stage_alu_shifter_n115), .B1(dp_ex_stage_alu_shifter_N112), 
        .B2(dp_ex_stage_alu_shifter_n112), .C1(dp_ex_stage_alu_shifter_N144), 
        .C2(dp_ex_stage_alu_shifter_n109), .ZN(dp_ex_stage_alu_shifter_n32) );
  AOI222_X1 dp_ex_stage_alu_shifter_U38 ( .A1(dp_ex_stage_alu_shifter_N227), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N130), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N162), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n56) );
  AOI222_X1 dp_ex_stage_alu_shifter_U37 ( .A1(dp_ex_stage_alu_shifter_N228), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N131), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N163), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n54) );
  AOI222_X1 dp_ex_stage_alu_shifter_U36 ( .A1(dp_ex_stage_alu_shifter_N224), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N127), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N159), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n62) );
  AOI222_X1 dp_ex_stage_alu_shifter_U35 ( .A1(dp_ex_stage_alu_shifter_N223), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N126), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N158), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n64) );
  AOI222_X1 dp_ex_stage_alu_shifter_U34 ( .A1(dp_ex_stage_alu_shifter_N225), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N128), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N160), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n60) );
  AOI222_X1 dp_ex_stage_alu_shifter_U33 ( .A1(dp_ex_stage_alu_shifter_N226), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N129), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N161), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n58) );
  AOI222_X1 dp_ex_stage_alu_shifter_U32 ( .A1(dp_ex_stage_alu_shifter_N222), 
        .A2(dp_ex_stage_alu_shifter_n114), .B1(dp_ex_stage_alu_shifter_N125), 
        .B2(dp_ex_stage_alu_shifter_n111), .C1(dp_ex_stage_alu_shifter_N157), 
        .C2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n66) );
  AND3_X1 dp_ex_stage_alu_shifter_U31 ( .A1(dp_ex_stage_alu_shifter_n95), .A2(
        dp_ex_stage_alu_shifter_n96), .A3(dp_ex_stage_alu_shifter_n97), .ZN(
        dp_ex_stage_alu_shifter_n84) );
  NAND2_X1 dp_ex_stage_alu_shifter_U30 ( .A1(dp_ex_stage_alu_shifter_N149), 
        .A2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n97) );
  NAND2_X1 dp_ex_stage_alu_shifter_U29 ( .A1(dp_ex_stage_alu_shifter_N117), 
        .A2(dp_ex_stage_alu_shifter_n110), .ZN(dp_ex_stage_alu_shifter_n96) );
  NAND2_X1 dp_ex_stage_alu_shifter_U28 ( .A1(dp_ex_stage_alu_shifter_N214), 
        .A2(dp_ex_stage_alu_shifter_n113), .ZN(dp_ex_stage_alu_shifter_n95) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_U27 ( .A(dp_ex_stage_muxA_out[24]), .Z(
        dp_ex_stage_alu_shifter_n94) );
  NOR3_X1 dp_ex_stage_alu_shifter_U26 ( .A1(dp_ex_stage_alu_shifter_n93), .A2(
        dp_ex_stage_alu_shifter_n20), .A3(dp_ex_stage_alu_shifter_n19), .ZN(
        dp_ex_stage_alu_shifter_n90) );
  AND2_X1 dp_ex_stage_alu_shifter_U25 ( .A1(dp_ex_stage_alu_shifter_N137), 
        .A2(dp_ex_stage_alu_shifter_n107), .ZN(dp_ex_stage_alu_shifter_n93) );
  AND2_X1 dp_ex_stage_alu_shifter_U24 ( .A1(dp_ex_stage_alu_shifter_N105), 
        .A2(dp_ex_stage_alu_shifter_n110), .ZN(dp_ex_stage_alu_shifter_n20) );
  AND2_X1 dp_ex_stage_alu_shifter_U23 ( .A1(dp_ex_stage_alu_shifter_N202), 
        .A2(dp_ex_stage_alu_shifter_n113), .ZN(dp_ex_stage_alu_shifter_n19) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_U22 ( .A(dp_ex_stage_muxA_out[27]), .Z(
        dp_ex_stage_alu_shifter_n12) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_U21 ( .A(dp_ex_stage_muxA_out[26]), .Z(
        dp_ex_stage_alu_shifter_n11) );
  AND3_X1 dp_ex_stage_alu_shifter_U20 ( .A1(dp_ex_stage_alu_shifter_n8), .A2(
        dp_ex_stage_alu_shifter_n9), .A3(dp_ex_stage_alu_shifter_n10), .ZN(
        dp_ex_stage_alu_shifter_n46) );
  NAND2_X1 dp_ex_stage_alu_shifter_U19 ( .A1(dp_ex_stage_alu_shifter_N139), 
        .A2(dp_ex_stage_alu_shifter_n108), .ZN(dp_ex_stage_alu_shifter_n10) );
  NAND2_X1 dp_ex_stage_alu_shifter_U18 ( .A1(dp_ex_stage_alu_shifter_N107), 
        .A2(dp_ex_stage_alu_shifter_n111), .ZN(dp_ex_stage_alu_shifter_n9) );
  NAND2_X1 dp_ex_stage_alu_shifter_U17 ( .A1(dp_ex_stage_alu_shifter_N204), 
        .A2(dp_ex_stage_alu_shifter_n114), .ZN(dp_ex_stage_alu_shifter_n8) );
  INV_X1 dp_ex_stage_alu_shifter_U16 ( .A(dp_ex_stage_alu_shifter_n6), .ZN(
        dp_ex_stage_alu_shifter_n7) );
  INV_X1 dp_ex_stage_alu_shifter_U15 ( .A(dp_ex_stage_muxA_out[25]), .ZN(
        dp_ex_stage_alu_shifter_n6) );
  INV_X2 dp_ex_stage_alu_shifter_U14 ( .A(dp_ex_stage_alu_shifter_n4), .ZN(
        dp_ex_stage_alu_shifter_n5) );
  INV_X1 dp_ex_stage_alu_shifter_U13 ( .A(dp_ex_stage_alu_n46), .ZN(
        dp_ex_stage_alu_shifter_n4) );
  INV_X1 dp_ex_stage_alu_shifter_U10 ( .A(dp_ex_stage_alu_shifter_n2), .ZN(
        dp_ex_stage_alu_shifter_n3) );
  INV_X1 dp_ex_stage_alu_shifter_U9 ( .A(dp_ex_stage_alu_n45), .ZN(
        dp_ex_stage_alu_shifter_n2) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_U8 ( .A(dp_ex_stage_muxA_out[31]), .Z(
        dp_ex_stage_alu_shifter_n1) );
  BUF_X1 dp_ex_stage_alu_shifter_U7 ( .A(dp_ex_stage_alu_shifter_n25), .Z(
        dp_ex_stage_alu_shifter_n107) );
  BUF_X1 dp_ex_stage_alu_shifter_U6 ( .A(dp_ex_stage_alu_shifter_n24), .Z(
        dp_ex_stage_alu_shifter_n110) );
  BUF_X1 dp_ex_stage_alu_shifter_U5 ( .A(dp_ex_stage_alu_shifter_n25), .Z(
        dp_ex_stage_alu_shifter_n108) );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U59 ( .A1(
        dp_ex_stage_alu_shifter_N202), .A2(dp_ex_stage_alu_shifter_sll_48_n4), 
        .ZN(dp_ex_stage_alu_shifter_sll_48_ML_int_1__0_) );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U58 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__0_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n8), .ZN(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__0_) );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U57 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__1_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n8), .ZN(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__1_) );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U56 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__0_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n12), .ZN(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__0_) );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U55 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__1_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n12), .ZN(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__1_) );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U54 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__2_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n12), .ZN(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__2_) );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U53 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__3_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n12), .ZN(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__3_) );
  NAND2_X1 dp_ex_stage_alu_shifter_sll_48_U52 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__0_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n34) );
  NAND2_X1 dp_ex_stage_alu_shifter_sll_48_U51 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__1_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n33) );
  NAND2_X1 dp_ex_stage_alu_shifter_sll_48_U50 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__2_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n32) );
  NAND2_X1 dp_ex_stage_alu_shifter_sll_48_U49 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__3_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n31) );
  NAND2_X1 dp_ex_stage_alu_shifter_sll_48_U48 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__4_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n30) );
  NAND2_X1 dp_ex_stage_alu_shifter_sll_48_U47 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__5_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n29) );
  NAND2_X1 dp_ex_stage_alu_shifter_sll_48_U46 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__6_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n28) );
  NAND2_X1 dp_ex_stage_alu_shifter_sll_48_U45 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__7_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n27) );
  NOR2_X1 dp_ex_stage_alu_shifter_sll_48_U44 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_n17), .A2(
        dp_ex_stage_alu_shifter_sll_48_n34), .ZN(dp_ex_stage_alu_shifter_N234)
         );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U43 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__10_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(dp_ex_stage_alu_shifter_N244)
         );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U42 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__11_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(dp_ex_stage_alu_shifter_N245)
         );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U41 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__12_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(dp_ex_stage_alu_shifter_N246)
         );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U40 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__13_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(dp_ex_stage_alu_shifter_N247)
         );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U39 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__14_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(dp_ex_stage_alu_shifter_N248)
         );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U38 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__15_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(dp_ex_stage_alu_shifter_N249)
         );
  NOR2_X1 dp_ex_stage_alu_shifter_sll_48_U37 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_n17), .A2(
        dp_ex_stage_alu_shifter_sll_48_n33), .ZN(dp_ex_stage_alu_shifter_N235)
         );
  NOR2_X1 dp_ex_stage_alu_shifter_sll_48_U36 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_n17), .A2(
        dp_ex_stage_alu_shifter_sll_48_n32), .ZN(dp_ex_stage_alu_shifter_N236)
         );
  NOR2_X1 dp_ex_stage_alu_shifter_sll_48_U35 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_n17), .A2(
        dp_ex_stage_alu_shifter_sll_48_n31), .ZN(dp_ex_stage_alu_shifter_N237)
         );
  NOR2_X1 dp_ex_stage_alu_shifter_sll_48_U34 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_n17), .A2(
        dp_ex_stage_alu_shifter_sll_48_n30), .ZN(dp_ex_stage_alu_shifter_N238)
         );
  NOR2_X1 dp_ex_stage_alu_shifter_sll_48_U33 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_n17), .A2(
        dp_ex_stage_alu_shifter_sll_48_n29), .ZN(dp_ex_stage_alu_shifter_N239)
         );
  NOR2_X1 dp_ex_stage_alu_shifter_sll_48_U32 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_n17), .A2(
        dp_ex_stage_alu_shifter_sll_48_n28), .ZN(dp_ex_stage_alu_shifter_N240)
         );
  NOR2_X1 dp_ex_stage_alu_shifter_sll_48_U31 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_n17), .A2(
        dp_ex_stage_alu_shifter_sll_48_n27), .ZN(dp_ex_stage_alu_shifter_N241)
         );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U30 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__8_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(dp_ex_stage_alu_shifter_N242)
         );
  AND2_X1 dp_ex_stage_alu_shifter_sll_48_U29 ( .A1(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__9_), .A2(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(dp_ex_stage_alu_shifter_N243)
         );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U28 ( .A(dp_ex_stage_alu_shifter_n116), 
        .ZN(dp_ex_stage_alu_shifter_sll_48_n18) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U27 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n14) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U26 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n15), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n13) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U25 ( .A(dp_ex_stage_alu_n49), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n12) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U24 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n12), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n11) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U23 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n8), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n7) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U22 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n4), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n3) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U21 ( .A(dp_ex_stage_alu_shifter_n5), 
        .ZN(dp_ex_stage_alu_shifter_sll_48_n8) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U20 ( .A(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n15) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U19 ( .A(dp_ex_stage_alu_n45), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n4) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U18 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n4), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n2) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U17 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n4), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n1) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U16 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n33), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n23) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U15 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n32), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n21) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U14 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n31), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n25) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U13 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n34), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n19) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U12 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n28), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n22) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U11 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n27), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n26) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U10 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n29), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n24) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U9 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n30), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n20) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U8 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n8), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n6) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U7 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n8), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n5) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U6 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n12), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n10) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U5 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n12), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n9) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U4 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n17) );
  INV_X1 dp_ex_stage_alu_shifter_sll_48_U3 ( .A(
        dp_ex_stage_alu_shifter_sll_48_n18), .ZN(
        dp_ex_stage_alu_shifter_sll_48_n16) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_1 ( .A(dp_ex_stage_alu_n76), .B(
        dp_ex_stage_alu_shifter_N202), .S(dp_ex_stage_alu_shifter_sll_48_n1), 
        .Z(dp_ex_stage_alu_shifter_sll_48_ML_int_1__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_2 ( .A(dp_ex_stage_alu_n44), .B(
        dp_ex_stage_alu_n76), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_3 ( .A(dp_ex_stage_alu_n69), .B(
        dp_ex_stage_alu_n44), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_4 ( .A(dp_ex_stage_alu_n52), .B(
        dp_ex_stage_alu_n69), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_5 ( .A(dp_ex_stage_alu_n70), .B(
        dp_ex_stage_alu_n52), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_6 ( .A(dp_ex_stage_alu_n78), .B(
        dp_ex_stage_alu_n70), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_7 ( .A(dp_ex_stage_alu_n34), .B(
        dp_ex_stage_alu_n78), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_8 ( .A(dp_ex_stage_alu_n71), .B(
        dp_ex_stage_alu_n34), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_9 ( .A(dp_ex_stage_alu_n72), .B(
        dp_ex_stage_alu_n71), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_10 ( .A(dp_ex_stage_alu_n74), 
        .B(dp_ex_stage_alu_n72), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_11 ( .A(dp_ex_stage_alu_n33), 
        .B(dp_ex_stage_alu_n74), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_12 ( .A(dp_ex_stage_muxA_out[12]), .B(dp_ex_stage_alu_n33), .S(dp_ex_stage_alu_shifter_sll_48_n1), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_13 ( .A(dp_ex_stage_alu_n231), 
        .B(dp_ex_stage_muxA_out[12]), .S(dp_ex_stage_alu_shifter_sll_48_n2), 
        .Z(dp_ex_stage_alu_shifter_sll_48_ML_int_1__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_14 ( .A(dp_ex_stage_muxA_out[14]), .B(dp_ex_stage_alu_n231), .S(dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_15 ( .A(dp_ex_stage_alu_n29), 
        .B(dp_ex_stage_muxA_out[14]), .S(dp_ex_stage_alu_shifter_sll_48_n2), 
        .Z(dp_ex_stage_alu_shifter_sll_48_ML_int_1__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_16 ( .A(dp_ex_stage_alu_n38), 
        .B(dp_ex_stage_alu_n29), .S(dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_17 ( .A(dp_ex_stage_muxA_out[17]), .B(dp_ex_stage_alu_n38), .S(dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_18 ( .A(dp_ex_stage_muxA_out[18]), .B(dp_ex_stage_muxA_out[17]), .S(dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_19 ( .A(dp_ex_stage_muxA_out[19]), .B(dp_ex_stage_muxA_out[18]), .S(dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_20 ( .A(dp_ex_stage_muxA_out[20]), .B(dp_ex_stage_muxA_out[19]), .S(dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_21 ( .A(dp_ex_stage_muxA_out[21]), .B(dp_ex_stage_muxA_out[20]), .S(dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_22 ( .A(dp_ex_stage_alu_n240), 
        .B(dp_ex_stage_muxA_out[21]), .S(dp_ex_stage_alu_shifter_sll_48_n2), 
        .Z(dp_ex_stage_alu_shifter_sll_48_ML_int_1__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_23 ( .A(dp_ex_stage_muxA_out[23]), .B(dp_ex_stage_alu_n240), .S(dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_24 ( .A(
        dp_ex_stage_alu_shifter_n94), .B(dp_ex_stage_muxA_out[23]), .S(
        dp_ex_stage_alu_shifter_sll_48_n2), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_25 ( .A(
        dp_ex_stage_alu_shifter_n7), .B(dp_ex_stage_alu_shifter_n94), .S(
        dp_ex_stage_alu_shifter_sll_48_n3), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_26 ( .A(
        dp_ex_stage_alu_shifter_n11), .B(dp_ex_stage_alu_shifter_n7), .S(
        dp_ex_stage_alu_shifter_sll_48_n3), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_27 ( .A(
        dp_ex_stage_alu_shifter_n12), .B(dp_ex_stage_alu_shifter_n11), .S(
        dp_ex_stage_alu_shifter_sll_48_n3), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_28 ( .A(dp_ex_stage_alu_n1), .B(
        dp_ex_stage_alu_shifter_n12), .S(dp_ex_stage_alu_shifter_sll_48_n3), 
        .Z(dp_ex_stage_alu_shifter_sll_48_ML_int_1__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_29 ( .A(dp_ex_stage_muxA_out[29]), .B(dp_ex_stage_alu_n1), .S(dp_ex_stage_alu_shifter_sll_48_n3), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_30 ( .A(dp_ex_stage_muxA_out[30]), .B(dp_ex_stage_muxA_out[29]), .S(dp_ex_stage_alu_shifter_sll_48_n3), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_0_31 ( .A(dp_ex_stage_muxA_out[31]), .B(dp_ex_stage_muxA_out[30]), .S(dp_ex_stage_alu_shifter_sll_48_n3), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_2 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__2_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__0_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_3 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__3_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__1_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_4 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__4_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__2_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_5 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__5_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__3_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_6 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__6_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__4_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_7 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__7_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__5_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_8 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__8_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__6_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_9 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__9_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__7_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_10 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__10_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__8_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_11 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__11_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__9_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_12 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__12_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__10_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_13 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__13_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__11_), .S(
        dp_ex_stage_alu_shifter_sll_48_n5), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_14 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__14_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__12_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_15 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__15_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__13_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_16 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__16_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__14_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_17 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__17_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__15_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_18 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__18_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__16_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_19 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__19_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__17_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_20 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__20_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__18_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_21 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__21_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__19_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_22 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__22_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__20_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_23 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__23_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__21_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_24 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__24_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__22_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_25 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__25_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__23_), .S(
        dp_ex_stage_alu_shifter_sll_48_n6), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_26 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__26_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__24_), .S(
        dp_ex_stage_alu_shifter_sll_48_n7), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_27 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__27_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__25_), .S(
        dp_ex_stage_alu_shifter_sll_48_n7), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_28 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__28_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__26_), .S(
        dp_ex_stage_alu_shifter_sll_48_n7), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_29 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__29_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__27_), .S(
        dp_ex_stage_alu_shifter_sll_48_n7), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_30 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__30_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__28_), .S(
        dp_ex_stage_alu_shifter_sll_48_n7), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_1_31 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__31_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_1__29_), .S(
        dp_ex_stage_alu_shifter_sll_48_n7), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_4 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__4_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__0_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_5 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__5_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__1_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_6 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__6_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__2_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_7 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__7_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__3_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_8 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__8_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__4_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_9 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__9_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__5_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_10 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__10_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__6_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_11 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__11_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__7_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_12 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__12_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__8_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_13 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__13_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__9_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_14 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__14_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__10_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_15 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__15_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__11_), .S(
        dp_ex_stage_alu_shifter_sll_48_n9), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_16 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__16_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__12_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_17 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__17_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__13_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_18 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__18_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__14_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_19 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__19_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__15_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_20 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__20_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__16_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_21 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__21_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__17_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_22 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__22_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__18_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_23 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__23_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__19_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_24 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__24_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__20_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_25 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__25_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__21_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_26 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__26_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__22_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_27 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__27_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__23_), .S(
        dp_ex_stage_alu_shifter_sll_48_n10), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_28 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__28_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__24_), .S(
        dp_ex_stage_alu_shifter_sll_48_n11), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_29 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__29_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__25_), .S(
        dp_ex_stage_alu_shifter_sll_48_n11), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_30 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__30_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__26_), .S(
        dp_ex_stage_alu_shifter_sll_48_n11), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_2_31 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__31_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_2__27_), .S(
        dp_ex_stage_alu_shifter_sll_48_n11), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_8 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__8_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__0_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_9 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__9_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__1_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_10 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__10_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__2_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_11 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__11_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__3_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_12 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__12_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__4_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_13 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__13_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__5_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_14 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__14_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__6_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_15 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__15_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__7_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_16 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__16_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__8_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_17 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__17_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__9_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_18 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__18_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__10_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_19 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__19_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__11_), .S(
        dp_ex_stage_alu_shifter_sll_48_n13), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_20 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__20_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__12_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_21 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__21_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__13_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_22 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__22_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__14_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_23 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__23_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__15_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_24 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__24_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__16_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_25 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__25_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__17_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_26 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__26_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__18_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_27 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__27_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__19_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_28 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__28_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__20_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_29 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__29_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__21_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_30 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__30_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__22_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_3_31 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__31_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_3__23_), .S(
        dp_ex_stage_alu_shifter_sll_48_n14), .Z(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_16 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__16_), .B(
        dp_ex_stage_alu_shifter_sll_48_n19), .S(
        dp_ex_stage_alu_shifter_sll_48_n17), .Z(dp_ex_stage_alu_shifter_N250)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_17 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__17_), .B(
        dp_ex_stage_alu_shifter_sll_48_n23), .S(
        dp_ex_stage_alu_shifter_sll_48_n17), .Z(dp_ex_stage_alu_shifter_N251)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_18 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__18_), .B(
        dp_ex_stage_alu_shifter_sll_48_n21), .S(
        dp_ex_stage_alu_shifter_sll_48_n17), .Z(dp_ex_stage_alu_shifter_N252)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_19 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__19_), .B(
        dp_ex_stage_alu_shifter_sll_48_n25), .S(
        dp_ex_stage_alu_shifter_sll_48_n17), .Z(dp_ex_stage_alu_shifter_N253)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_20 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__20_), .B(
        dp_ex_stage_alu_shifter_sll_48_n20), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N254)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_21 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__21_), .B(
        dp_ex_stage_alu_shifter_sll_48_n24), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N255)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_22 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__22_), .B(
        dp_ex_stage_alu_shifter_sll_48_n22), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N256)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_23 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__23_), .B(
        dp_ex_stage_alu_shifter_sll_48_n26), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N257)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_24 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__24_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__8_), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N258)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_25 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__25_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__9_), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N259)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_26 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__26_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__10_), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N260)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_27 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__27_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__11_), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N261)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_28 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__28_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__12_), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N262)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_29 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__29_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__13_), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N263)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_30 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__30_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__14_), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N264)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sll_48_M1_4_31 ( .A(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__31_), .B(
        dp_ex_stage_alu_shifter_sll_48_ML_int_4__15_), .S(
        dp_ex_stage_alu_shifter_sll_48_n16), .Z(dp_ex_stage_alu_shifter_N265)
         );
  NAND2_X1 dp_ex_stage_alu_shifter_sla_46_U225 ( .A1(
        dp_ex_stage_alu_shifter_n5), .A2(dp_ex_stage_alu_shifter_sla_46_n13), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n95) );
  NAND2_X1 dp_ex_stage_alu_shifter_sla_46_U224 ( .A1(dp_ex_stage_alu_n45), 
        .A2(dp_ex_stage_alu_shifter_n5), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n96) );
  NOR2_X1 dp_ex_stage_alu_shifter_sla_46_U223 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n13), .A2(dp_ex_stage_alu_shifter_n5), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n98) );
  NOR2_X1 dp_ex_stage_alu_shifter_sla_46_U222 ( .A1(dp_ex_stage_alu_n45), .A2(
        dp_ex_stage_alu_shifter_n5), .ZN(dp_ex_stage_alu_shifter_sla_46_n99)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U221 ( .A1(dp_ex_stage_alu_n70), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n7), .B1(dp_ex_stage_alu_n78), .B2(
        dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n193) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U220 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n57), .C1(
        dp_ex_stage_alu_shifter_sla_46_n20), .C2(
        dp_ex_stage_alu_shifter_sla_46_n4), .A(
        dp_ex_stage_alu_shifter_sla_46_n193), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n155) );
  NOR2_X1 dp_ex_stage_alu_shifter_sla_46_U219 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n14), .A2(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n133) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U218 ( .A1(dp_ex_stage_alu_n72), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n9), .B1(
        dp_ex_stage_alu_shifter_sla_46_n24), .B2(
        dp_ex_stage_alu_shifter_sla_46_n12), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n192) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U217 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n3), .B2(
        dp_ex_stage_alu_shifter_sla_46_n22), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n21), .A(
        dp_ex_stage_alu_shifter_sla_46_n192), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n154) );
  AND2_X1 dp_ex_stage_alu_shifter_sla_46_U216 ( .A1(dp_ex_stage_alu_n31), .A2(
        dp_ex_stage_alu_shifter_sla_46_n14), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n137) );
  NAND2_X1 dp_ex_stage_alu_shifter_sla_46_U215 ( .A1(dp_ex_stage_alu_n31), 
        .A2(dp_ex_stage_alu_shifter_N202), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n158) );
  NOR2_X1 dp_ex_stage_alu_shifter_sla_46_U214 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n14), .A2(
        dp_ex_stage_alu_shifter_sla_46_n158), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n139) );
  AOI21_X1 dp_ex_stage_alu_shifter_sla_46_U213 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n137), .B2(
        dp_ex_stage_alu_shifter_sla_46_n48), .A(
        dp_ex_stage_alu_shifter_sla_46_n139), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n190) );
  NAND2_X1 dp_ex_stage_alu_shifter_sla_46_U212 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n17), .A2(dp_ex_stage_alu_shifter_N202), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n80) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U211 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n17), .B2(
        dp_ex_stage_alu_shifter_sla_46_n125), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N212)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U210 ( .A1(dp_ex_stage_alu_n78), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n9), .B1(dp_ex_stage_alu_n34), .B2(
        dp_ex_stage_alu_shifter_sla_46_n12), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n189) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U209 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n3), .B2(
        dp_ex_stage_alu_shifter_sla_46_n58), .C1(
        dp_ex_stage_alu_shifter_sla_46_n6), .C2(
        dp_ex_stage_alu_shifter_sla_46_n57), .A(
        dp_ex_stage_alu_shifter_sla_46_n189), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n151) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U208 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n24), .A2(
        dp_ex_stage_alu_shifter_sla_46_n9), .B1(dp_ex_stage_alu_n33), .B2(
        dp_ex_stage_alu_shifter_sla_46_n12), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n188) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U207 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n3), .B2(
        dp_ex_stage_alu_shifter_sla_46_n23), .C1(
        dp_ex_stage_alu_shifter_sla_46_n6), .C2(
        dp_ex_stage_alu_shifter_sla_46_n22), .A(
        dp_ex_stage_alu_shifter_sla_46_n188), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n149) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U206 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n9), .A2(dp_ex_stage_alu_n44), .B1(
        dp_ex_stage_alu_n69), .B2(dp_ex_stage_alu_shifter_sla_46_n12), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n187) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U205 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n56), .B2(
        dp_ex_stage_alu_shifter_sla_46_n3), .C1(
        dp_ex_stage_alu_shifter_sla_46_n55), .C2(
        dp_ex_stage_alu_shifter_sla_46_n4), .A(
        dp_ex_stage_alu_shifter_sla_46_n187), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n150) );
  AOI21_X1 dp_ex_stage_alu_shifter_sla_46_U204 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n137), .B2(
        dp_ex_stage_alu_shifter_sla_46_n150), .A(
        dp_ex_stage_alu_shifter_sla_46_n139), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n186) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U203 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n17), .B2(
        dp_ex_stage_alu_shifter_sla_46_n120), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N213)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U202 ( .A1(dp_ex_stage_alu_n34), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n8), .B1(dp_ex_stage_alu_n71), .B2(
        dp_ex_stage_alu_shifter_sla_46_n12), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n185) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U201 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n3), .B2(
        dp_ex_stage_alu_shifter_sla_46_n60), .C1(
        dp_ex_stage_alu_shifter_sla_46_n6), .C2(
        dp_ex_stage_alu_shifter_sla_46_n58), .A(
        dp_ex_stage_alu_shifter_sla_46_n185), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n145) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U200 ( .A1(dp_ex_stage_alu_n33), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n8), .B1(dp_ex_stage_muxA_out[12]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n184) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U199 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n25), .C1(
        dp_ex_stage_alu_shifter_sla_46_n6), .C2(
        dp_ex_stage_alu_shifter_sla_46_n23), .A(
        dp_ex_stage_alu_shifter_sla_46_n184), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n143) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U198 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n9), .A2(dp_ex_stage_alu_n69), .B1(
        dp_ex_stage_alu_n52), .B2(dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n183) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U197 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n19), .C1(
        dp_ex_stage_alu_shifter_sla_46_n56), .C2(
        dp_ex_stage_alu_shifter_sla_46_n4), .A(
        dp_ex_stage_alu_shifter_sla_46_n183), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n144) );
  AOI21_X1 dp_ex_stage_alu_shifter_sla_46_U196 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n137), .B2(
        dp_ex_stage_alu_shifter_sla_46_n144), .A(
        dp_ex_stage_alu_shifter_sla_46_n139), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n182) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U195 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n17), .B2(
        dp_ex_stage_alu_shifter_sla_46_n113), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N214)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_sla_46_U194 ( .A(
        dp_ex_stage_alu_shifter_N202), .B(dp_ex_stage_alu_n76), .S(
        dp_ex_stage_alu_shifter_sla_46_n10), .Z(
        dp_ex_stage_alu_shifter_sla_46_n138) );
  AND2_X1 dp_ex_stage_alu_shifter_sla_46_U193 ( .A1(dp_ex_stage_alu_n49), .A2(
        dp_ex_stage_alu_n31), .ZN(dp_ex_stage_alu_shifter_sla_46_n174) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U192 ( .A1(dp_ex_stage_alu_n52), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n8), .B1(dp_ex_stage_alu_n70), .B2(
        dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n181) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U191 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n20), .C1(
        dp_ex_stage_alu_shifter_sla_46_n6), .C2(
        dp_ex_stage_alu_shifter_sla_46_n19), .A(
        dp_ex_stage_alu_shifter_sla_46_n181), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n132) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U190 ( .A1(dp_ex_stage_alu_n71), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n8), .B1(dp_ex_stage_alu_n72), .B2(
        dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n180) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U189 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n21), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n60), .A(
        dp_ex_stage_alu_shifter_sla_46_n180), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n134) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U188 ( .A1(dp_ex_stage_muxA_out[12]), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n8), .B1(
        dp_ex_stage_alu_shifter_sla_46_n28), .B2(
        dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n179) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U187 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n26), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n25), .A(
        dp_ex_stage_alu_shifter_sla_46_n179), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n131) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U186 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n133), .A2(
        dp_ex_stage_alu_shifter_sla_46_n134), .B1(
        dp_ex_stage_alu_shifter_sla_46_n131), .B2(
        dp_ex_stage_alu_shifter_sla_46_n135), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n178) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U185 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n138), .B2(
        dp_ex_stage_alu_shifter_sla_46_n174), .C1(
        dp_ex_stage_alu_shifter_sla_46_n132), .C2(
        dp_ex_stage_alu_shifter_sla_46_n137), .A(
        dp_ex_stage_alu_shifter_sla_46_n59), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n107) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U184 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n16), .B2(
        dp_ex_stage_alu_shifter_sla_46_n107), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N215)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U183 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n28), .A2(
        dp_ex_stage_alu_shifter_sla_46_n8), .B1(
        dp_ex_stage_alu_shifter_sla_46_n30), .B2(
        dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n177) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U182 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n27), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n26), .A(
        dp_ex_stage_alu_shifter_sla_46_n177), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n127) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U181 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n174), .A2(
        dp_ex_stage_alu_shifter_sla_46_n48), .B1(
        dp_ex_stage_alu_shifter_sla_46_n137), .B2(
        dp_ex_stage_alu_shifter_sla_46_n155), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n176) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U180 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n154), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n127), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n47), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n100) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U179 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n16), .B2(
        dp_ex_stage_alu_shifter_sla_46_n100), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N216)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U178 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n30), .A2(
        dp_ex_stage_alu_shifter_sla_46_n8), .B1(dp_ex_stage_alu_n29), .B2(
        dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n175) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U177 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n29), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n27), .A(
        dp_ex_stage_alu_shifter_sla_46_n175), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n122) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U176 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n174), .A2(
        dp_ex_stage_alu_shifter_sla_46_n150), .B1(
        dp_ex_stage_alu_shifter_sla_46_n137), .B2(
        dp_ex_stage_alu_shifter_sla_46_n151), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n173) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U175 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n149), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n122), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n54), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n88) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U174 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n16), .B2(
        dp_ex_stage_alu_shifter_sla_46_n88), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N217)
         );
  NAND2_X1 dp_ex_stage_alu_shifter_sla_46_U173 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n133), .A2(
        dp_ex_stage_alu_shifter_sla_46_n18), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n87) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U172 ( .A1(dp_ex_stage_alu_n29), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n8), .B1(
        dp_ex_stage_alu_shifter_sla_46_n33), .B2(
        dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n172) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U171 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n31), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n29), .A(
        dp_ex_stage_alu_shifter_sla_46_n172), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n115) );
  AND2_X1 dp_ex_stage_alu_shifter_sla_46_U170 ( .A1(dp_ex_stage_alu_n31), .A2(
        dp_ex_stage_alu_shifter_sla_46_n18), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n171) );
  AND2_X1 dp_ex_stage_alu_shifter_sla_46_U169 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n171), .A2(dp_ex_stage_alu_n49), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n90) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U168 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n90), .B2(
        dp_ex_stage_alu_shifter_sla_46_n144), .C1(
        dp_ex_stage_alu_shifter_sla_46_n93), .C2(
        dp_ex_stage_alu_shifter_sla_46_n145), .A(
        dp_ex_stage_alu_shifter_sla_46_n53), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n170) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U167 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n61), .B2(
        dp_ex_stage_alu_shifter_sla_46_n87), .C1(
        dp_ex_stage_alu_shifter_sla_46_n62), .C2(
        dp_ex_stage_alu_shifter_sla_46_n119), .A(
        dp_ex_stage_alu_shifter_sla_46_n170), .ZN(dp_ex_stage_alu_shifter_N218) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U166 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n33), .A2(
        dp_ex_stage_alu_shifter_sla_46_n8), .B1(
        dp_ex_stage_alu_shifter_sla_46_n35), .B2(
        dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n169) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U165 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n32), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n31), .A(
        dp_ex_stage_alu_shifter_sla_46_n169), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n109) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U164 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n55), .B2(
        dp_ex_stage_alu_shifter_sla_46_n14), .A(
        dp_ex_stage_alu_shifter_sla_46_n158), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n161) );
  AOI21_X1 dp_ex_stage_alu_shifter_sla_46_U163 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n138), .B2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n161), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n163) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U162 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n131), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n134), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n132), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n168) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U161 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n63), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n163), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n168), .ZN(dp_ex_stage_alu_shifter_N219) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U160 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n35), .A2(
        dp_ex_stage_alu_shifter_sla_46_n8), .B1(dp_ex_stage_muxA_out[18]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n167) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U159 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n34), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n32), .A(
        dp_ex_stage_alu_shifter_sla_46_n167), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n102) );
  AOI21_X1 dp_ex_stage_alu_shifter_sla_46_U158 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n48), .B2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n161), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n106) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U157 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n127), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n154), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n155), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n166) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U156 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n64), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n106), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n166), .ZN(dp_ex_stage_alu_shifter_N220) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U155 ( .A1(dp_ex_stage_muxA_out[18]), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n8), .B1(dp_ex_stage_muxA_out[19]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n165) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U154 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n36), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n34), .A(
        dp_ex_stage_alu_shifter_sla_46_n165), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n91) );
  AOI21_X1 dp_ex_stage_alu_shifter_sla_46_U153 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n150), .B2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n161), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n86) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U152 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n122), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n149), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n151), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n164) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U151 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n65), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n86), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n164), .ZN(dp_ex_stage_alu_shifter_N221) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U150 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n16), .B2(
        dp_ex_stage_alu_shifter_sla_46_n163), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N203)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U149 ( .A1(dp_ex_stage_muxA_out[19]), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n7), .B1(dp_ex_stage_muxA_out[20]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n162) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U148 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n37), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n36), .A(
        dp_ex_stage_alu_shifter_sla_46_n162), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n117) );
  AOI21_X1 dp_ex_stage_alu_shifter_sla_46_U147 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n144), .B2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n161), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n85) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U146 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n115), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n143), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n145), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n160) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U145 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n66), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n85), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n160), .ZN(dp_ex_stage_alu_shifter_N222) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U144 ( .A1(dp_ex_stage_muxA_out[20]), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n7), .B1(dp_ex_stage_muxA_out[21]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n159) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U143 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n69), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n37), .A(
        dp_ex_stage_alu_shifter_sla_46_n159), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n111) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U142 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n109), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n131), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n134), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n157) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U141 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n67), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n84), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n157), .ZN(dp_ex_stage_alu_shifter_N223) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U140 ( .A1(dp_ex_stage_muxA_out[21]), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n7), .B1(dp_ex_stage_alu_n240), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n156) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U139 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n71), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n69), .A(
        dp_ex_stage_alu_shifter_sla_46_n156), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n104) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U138 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n102), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n127), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n154), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n153) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U137 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n68), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n83), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n153), .ZN(dp_ex_stage_alu_shifter_N224) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U136 ( .A1(dp_ex_stage_alu_n240), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n7), .B1(dp_ex_stage_muxA_out[23]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n152) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U135 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n38), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n71), .A(
        dp_ex_stage_alu_shifter_sla_46_n152), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n94) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U134 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n91), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n122), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n149), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n148) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U133 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n70), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n82), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n148), .ZN(dp_ex_stage_alu_shifter_N225) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U132 ( .A1(dp_ex_stage_muxA_out[23]), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n7), .B1(
        dp_ex_stage_alu_shifter_n94), .B2(dp_ex_stage_alu_shifter_sla_46_n10), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n147) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U131 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n39), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n38), .A(
        dp_ex_stage_alu_shifter_sla_46_n147), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n146) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U130 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n117), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n115), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n143), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n142) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U129 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n72), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n81), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n142), .ZN(dp_ex_stage_alu_shifter_N226) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U128 ( .A1(
        dp_ex_stage_alu_shifter_n94), .A2(dp_ex_stage_alu_shifter_sla_46_n7), 
        .B1(dp_ex_stage_alu_shifter_n7), .B2(
        dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n141) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U127 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n40), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n39), .A(
        dp_ex_stage_alu_shifter_sla_46_n141), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n140) );
  AOI21_X1 dp_ex_stage_alu_shifter_sla_46_U126 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n137), .B2(
        dp_ex_stage_alu_shifter_sla_46_n138), .A(
        dp_ex_stage_alu_shifter_sla_46_n139), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n136) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U125 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n132), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n134), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n51), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n79) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U124 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n111), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n109), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n131), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n130) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U123 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n73), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n79), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n130), .ZN(dp_ex_stage_alu_shifter_N227) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U122 ( .A1(
        dp_ex_stage_alu_shifter_n7), .A2(dp_ex_stage_alu_shifter_sla_46_n7), 
        .B1(dp_ex_stage_alu_shifter_n11), .B2(
        dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n129) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U121 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n41), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n40), .A(
        dp_ex_stage_alu_shifter_sla_46_n129), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n128) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U120 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n104), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n102), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n127), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n126) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U119 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n74), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n125), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n126), .ZN(dp_ex_stage_alu_shifter_N228) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U118 ( .A1(
        dp_ex_stage_alu_shifter_n11), .A2(dp_ex_stage_alu_shifter_sla_46_n7), 
        .B1(dp_ex_stage_alu_shifter_n12), .B2(
        dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n124) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U117 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n42), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n41), .A(
        dp_ex_stage_alu_shifter_sla_46_n124), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n123) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U116 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n78), .A2(
        dp_ex_stage_alu_shifter_sla_46_n94), .B1(
        dp_ex_stage_alu_shifter_sla_46_n93), .B2(
        dp_ex_stage_alu_shifter_sla_46_n91), .C1(
        dp_ex_stage_alu_shifter_sla_46_n90), .C2(
        dp_ex_stage_alu_shifter_sla_46_n122), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n121) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U115 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n75), .B2(
        dp_ex_stage_alu_shifter_sla_46_n119), .C1(
        dp_ex_stage_alu_shifter_sla_46_n120), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n121), .ZN(dp_ex_stage_alu_shifter_N229) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U114 ( .A1(
        dp_ex_stage_alu_shifter_n12), .A2(dp_ex_stage_alu_shifter_sla_46_n7), 
        .B1(dp_ex_stage_alu_n1), .B2(dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n118) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U113 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n43), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n42), .A(
        dp_ex_stage_alu_shifter_sla_46_n118), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n116) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U112 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n90), .A2(
        dp_ex_stage_alu_shifter_sla_46_n115), .B1(
        dp_ex_stage_alu_shifter_sla_46_n77), .B2(
        dp_ex_stage_alu_shifter_sla_46_n116), .C1(
        dp_ex_stage_alu_shifter_sla_46_n93), .C2(
        dp_ex_stage_alu_shifter_sla_46_n117), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n114) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U111 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n72), .B2(
        dp_ex_stage_alu_shifter_sla_46_n87), .C1(
        dp_ex_stage_alu_shifter_sla_46_n113), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n114), .ZN(dp_ex_stage_alu_shifter_N230) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U110 ( .A1(dp_ex_stage_alu_n1), .A2(
        dp_ex_stage_alu_shifter_sla_46_n7), .B1(dp_ex_stage_muxA_out[29]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n112) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U109 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n44), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n43), .A(
        dp_ex_stage_alu_shifter_sla_46_n112), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n110) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U108 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n90), .A2(
        dp_ex_stage_alu_shifter_sla_46_n109), .B1(
        dp_ex_stage_alu_shifter_sla_46_n77), .B2(
        dp_ex_stage_alu_shifter_sla_46_n110), .C1(
        dp_ex_stage_alu_shifter_sla_46_n93), .C2(
        dp_ex_stage_alu_shifter_sla_46_n111), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n108) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U107 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n73), .B2(
        dp_ex_stage_alu_shifter_sla_46_n87), .C1(
        dp_ex_stage_alu_shifter_sla_46_n107), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n108), .ZN(dp_ex_stage_alu_shifter_N231) );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U106 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n16), .B2(
        dp_ex_stage_alu_shifter_sla_46_n106), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N204)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U105 ( .A1(dp_ex_stage_muxA_out[29]), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n7), .B1(dp_ex_stage_muxA_out[30]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n10), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n105) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U104 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n1), .B2(
        dp_ex_stage_alu_shifter_sla_46_n45), .C1(
        dp_ex_stage_alu_shifter_sla_46_n4), .C2(
        dp_ex_stage_alu_shifter_sla_46_n44), .A(
        dp_ex_stage_alu_shifter_sla_46_n105), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n103) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U103 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n90), .A2(
        dp_ex_stage_alu_shifter_sla_46_n102), .B1(
        dp_ex_stage_alu_shifter_sla_46_n77), .B2(
        dp_ex_stage_alu_shifter_sla_46_n103), .C1(
        dp_ex_stage_alu_shifter_sla_46_n93), .C2(
        dp_ex_stage_alu_shifter_sla_46_n104), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n101) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U102 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n74), .B2(
        dp_ex_stage_alu_shifter_sla_46_n87), .C1(
        dp_ex_stage_alu_shifter_sla_46_n100), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n101), .ZN(dp_ex_stage_alu_shifter_N232) );
  AOI22_X1 dp_ex_stage_alu_shifter_sla_46_U101 ( .A1(dp_ex_stage_muxA_out[30]), 
        .A2(dp_ex_stage_alu_shifter_sla_46_n8), .B1(dp_ex_stage_muxA_out[31]), 
        .B2(dp_ex_stage_alu_shifter_sla_46_n11), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n97) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U100 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n2), .B2(
        dp_ex_stage_alu_shifter_sla_46_n76), .C1(
        dp_ex_stage_alu_shifter_sla_46_n5), .C2(
        dp_ex_stage_alu_shifter_sla_46_n45), .A(
        dp_ex_stage_alu_shifter_sla_46_n97), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n92) );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U99 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n90), .A2(
        dp_ex_stage_alu_shifter_sla_46_n91), .B1(
        dp_ex_stage_alu_shifter_sla_46_n77), .B2(
        dp_ex_stage_alu_shifter_sla_46_n92), .C1(
        dp_ex_stage_alu_shifter_sla_46_n93), .C2(
        dp_ex_stage_alu_shifter_sla_46_n94), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n89) );
  OAI221_X1 dp_ex_stage_alu_shifter_sla_46_U98 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n75), .B2(
        dp_ex_stage_alu_shifter_sla_46_n87), .C1(
        dp_ex_stage_alu_shifter_sla_46_n88), .C2(
        dp_ex_stage_alu_shifter_sla_46_n18), .A(
        dp_ex_stage_alu_shifter_sla_46_n89), .ZN(dp_ex_stage_alu_shifter_N233)
         );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U97 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n16), .B2(
        dp_ex_stage_alu_shifter_sla_46_n86), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N205)
         );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U96 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n16), .B2(
        dp_ex_stage_alu_shifter_sla_46_n85), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N206)
         );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U95 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n15), .B2(
        dp_ex_stage_alu_shifter_sla_46_n84), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N207)
         );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U94 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n15), .B2(
        dp_ex_stage_alu_shifter_sla_46_n83), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N208)
         );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U93 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n15), .B2(
        dp_ex_stage_alu_shifter_sla_46_n82), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N209)
         );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U92 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n15), .B2(
        dp_ex_stage_alu_shifter_sla_46_n81), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N210)
         );
  OAI21_X1 dp_ex_stage_alu_shifter_sla_46_U91 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n15), .B2(
        dp_ex_stage_alu_shifter_sla_46_n79), .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(dp_ex_stage_alu_shifter_N211)
         );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U90 ( .A(dp_ex_stage_alu_n1), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n45) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U89 ( .A(dp_ex_stage_alu_shifter_n12), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n44) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U88 ( .A(dp_ex_stage_alu_shifter_n11), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n43) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U87 ( .A(dp_ex_stage_alu_shifter_n7), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n42) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U86 ( .A(dp_ex_stage_alu_shifter_n94), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n41) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U85 ( .A(dp_ex_stage_muxA_out[23]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n40) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U84 ( .A(dp_ex_stage_alu_n240), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n39) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U83 ( .A(dp_ex_stage_muxA_out[21]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n38) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U82 ( .A(dp_ex_stage_muxA_out[18]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n37) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U81 ( .A(dp_ex_stage_muxA_out[17]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n36) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U80 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n36), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n35) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U79 ( .A(dp_ex_stage_alu_n38), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n34) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U78 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n34), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n33) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U77 ( .A(dp_ex_stage_alu_n29), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n32) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U76 ( .A(dp_ex_stage_muxA_out[14]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n31) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U75 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n31), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n30) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U74 ( .A(dp_ex_stage_alu_n231), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n29) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U73 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n29), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n28) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U72 ( .A(dp_ex_stage_muxA_out[12]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n27) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U71 ( .A(dp_ex_stage_alu_n33), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n26) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U70 ( .A(dp_ex_stage_alu_n74), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n25) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U69 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n25), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n24) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U68 ( .A(dp_ex_stage_alu_n72), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n23) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U67 ( .A(dp_ex_stage_alu_n71), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n22) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U66 ( .A(dp_ex_stage_alu_n34), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n21) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U65 ( .A(dp_ex_stage_alu_n69), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n20) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U64 ( .A(dp_ex_stage_alu_n44), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n19) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U63 ( .A(dp_ex_stage_alu_n49), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n14) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U62 ( .A(dp_ex_stage_alu_n45), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n13) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U61 ( .A(dp_ex_stage_alu_n52), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n57) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U60 ( .A(dp_ex_stage_alu_n78), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n60) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U59 ( .A(dp_ex_stage_alu_shifter_N202), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n55) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U58 ( .A(dp_ex_stage_alu_n70), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n58) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U57 ( .A(dp_ex_stage_alu_n76), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n56) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U56 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n191), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n48) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U55 ( .A(dp_ex_stage_muxA_out[20]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n71) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U54 ( .A(dp_ex_stage_muxA_out[19]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n69) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U53 ( .A(dp_ex_stage_muxA_out[29]), 
        .ZN(dp_ex_stage_alu_shifter_sla_46_n76) );
  BUF_X1 dp_ex_stage_alu_shifter_sla_46_U52 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n96), .Z(
        dp_ex_stage_alu_shifter_sla_46_n6) );
  BUF_X1 dp_ex_stage_alu_shifter_sla_46_U51 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n99), .Z(
        dp_ex_stage_alu_shifter_sla_46_n12) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U50 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n117), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n66) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U49 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n111), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n67) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U48 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n178), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n59) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U47 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n158), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n52) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U46 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n91), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n65) );
  BUF_X1 dp_ex_stage_alu_shifter_sla_46_U45 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n96), .Z(
        dp_ex_stage_alu_shifter_sla_46_n5) );
  BUF_X2 dp_ex_stage_alu_shifter_sla_46_U44 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n96), .Z(
        dp_ex_stage_alu_shifter_sla_46_n4) );
  AND2_X1 dp_ex_stage_alu_shifter_sla_46_U43 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n171), .A2(
        dp_ex_stage_alu_shifter_sla_46_n14), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n93) );
  BUF_X2 dp_ex_stage_alu_shifter_sla_46_U42 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n99), .Z(
        dp_ex_stage_alu_shifter_sla_46_n11) );
  BUF_X2 dp_ex_stage_alu_shifter_sla_46_U41 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n99), .Z(
        dp_ex_stage_alu_shifter_sla_46_n10) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U40 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n80), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n53) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U39 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n136), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n51) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U38 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n182), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n50) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U37 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n190), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n46) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U36 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n186), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n49) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U35 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n173), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n54) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U34 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n176), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n47) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U33 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n146), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n72) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U32 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n140), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n73) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U31 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n128), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n74) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U30 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n123), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n75) );
  BUF_X1 dp_ex_stage_alu_shifter_sla_46_U29 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n95), .Z(
        dp_ex_stage_alu_shifter_sla_46_n3) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U28 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n104), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n68) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U27 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n94), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n70) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U26 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n143), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n61) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U25 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n115), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n62) );
  BUF_X1 dp_ex_stage_alu_shifter_sla_46_U24 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n98), .Z(
        dp_ex_stage_alu_shifter_sla_46_n9) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U23 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n109), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n63) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U22 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n102), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n64) );
  BUF_X1 dp_ex_stage_alu_shifter_sla_46_U21 ( .A(dp_ex_stage_alu_shifter_n116), 
        .Z(dp_ex_stage_alu_shifter_sla_46_n15) );
  BUF_X2 dp_ex_stage_alu_shifter_sla_46_U20 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n95), .Z(
        dp_ex_stage_alu_shifter_sla_46_n1) );
  BUF_X2 dp_ex_stage_alu_shifter_sla_46_U19 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n95), .Z(
        dp_ex_stage_alu_shifter_sla_46_n2) );
  BUF_X1 dp_ex_stage_alu_shifter_sla_46_U18 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n98), .Z(
        dp_ex_stage_alu_shifter_sla_46_n8) );
  BUF_X1 dp_ex_stage_alu_shifter_sla_46_U17 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n98), .Z(
        dp_ex_stage_alu_shifter_sla_46_n7) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U16 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n119), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n77) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U15 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n87), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n78) );
  INV_X1 dp_ex_stage_alu_shifter_sla_46_U14 ( .A(
        dp_ex_stage_alu_shifter_sla_46_n15), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n18) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_sla_46_U13 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_sla_46_n17)
         );
  CLKBUF_X1 dp_ex_stage_alu_shifter_sla_46_U12 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_sla_46_n16)
         );
  AOI222_X1 dp_ex_stage_alu_shifter_sla_46_U11 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n10), .A2(dp_ex_stage_alu_n44), .B1(
        dp_ex_stage_alu_n76), .B2(dp_ex_stage_alu_shifter_sla_46_n9), .C1(
        dp_ex_stage_alu_shifter_N202), .C2(dp_ex_stage_alu_shifter_n5), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n191) );
  NOR2_X2 dp_ex_stage_alu_shifter_sla_46_U10 ( .A1(dp_ex_stage_alu_n49), .A2(
        dp_ex_stage_alu_n31), .ZN(dp_ex_stage_alu_shifter_sla_46_n135) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U9 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n150), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n151), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n52), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n82) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U8 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n151), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n149), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n49), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n120) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U7 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n155), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n154), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n46), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n125) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U6 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n145), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n143), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n50), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n113) );
  NAND2_X2 dp_ex_stage_alu_shifter_sla_46_U5 ( .A1(
        dp_ex_stage_alu_shifter_sla_46_n135), .A2(
        dp_ex_stage_alu_shifter_sla_46_n18), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n119) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U4 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n138), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n132), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n52), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n84) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U3 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n48), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n155), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n52), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n83) );
  AOI221_X1 dp_ex_stage_alu_shifter_sla_46_U2 ( .B1(
        dp_ex_stage_alu_shifter_sla_46_n144), .B2(
        dp_ex_stage_alu_shifter_sla_46_n133), .C1(
        dp_ex_stage_alu_shifter_sla_46_n145), .C2(
        dp_ex_stage_alu_shifter_sla_46_n135), .A(
        dp_ex_stage_alu_shifter_sla_46_n52), .ZN(
        dp_ex_stage_alu_shifter_sla_46_n81) );
  NAND2_X1 dp_ex_stage_alu_shifter_srl_41_U222 ( .A1(dp_ex_stage_alu_n46), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n3), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n120) );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U221 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n55), .A2(
        dp_ex_stage_alu_shifter_srl_41_n78), .B1(
        dp_ex_stage_alu_shifter_srl_41_n54), .B2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n189) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U220 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n24), .A2(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n137) );
  NAND2_X1 dp_ex_stage_alu_shifter_srl_41_U219 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n137), .A2(
        dp_ex_stage_alu_shifter_srl_41_n29), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n114) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U218 ( .A1(dp_ex_stage_muxA_out[23]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n79), .B1(dp_ex_stage_alu_n240), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n77), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n188) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U217 ( .A1(dp_ex_stage_muxA_out[17]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_alu_n38), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n187) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U216 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n68), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n45), .A(
        dp_ex_stage_alu_shifter_srl_41_n187), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n96) );
  NAND2_X1 dp_ex_stage_alu_shifter_srl_41_U215 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n24), .A2(
        dp_ex_stage_alu_shifter_srl_41_n25), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n164) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U214 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n24), .A2(
        dp_ex_stage_alu_shifter_srl_41_n25), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n152) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U213 ( .A1(dp_ex_stage_muxA_out[29]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_alu_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n186) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U212 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n25), .A2(dp_ex_stage_alu_n49), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n140) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U211 ( .A1(dp_ex_stage_muxA_out[25]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_muxA_out[24]), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n185) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U210 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n119), .B2(
        dp_ex_stage_alu_shifter_srl_41_n51), .C1(
        dp_ex_stage_alu_shifter_srl_41_n21), .C2(
        dp_ex_stage_alu_shifter_srl_41_n50), .A(
        dp_ex_stage_alu_shifter_srl_41_n185), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n138) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U209 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n152), .A2(
        dp_ex_stage_alu_shifter_srl_41_n134), .B1(
        dp_ex_stage_alu_shifter_srl_41_n140), .B2(
        dp_ex_stage_alu_shifter_srl_41_n138), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n184) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U208 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n97), .B2(
        dp_ex_stage_alu_shifter_srl_41_n137), .C1(
        dp_ex_stage_alu_shifter_srl_41_n96), .C2(
        dp_ex_stage_alu_shifter_srl_41_n82), .A(
        dp_ex_stage_alu_shifter_srl_41_n70), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n154) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U207 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n25), .A2(
        dp_ex_stage_alu_shifter_srl_41_n28), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n181) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U206 ( .A1(dp_ex_stage_alu_n231), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(
        dp_ex_stage_alu_shifter_srl_41_n37), .B2(
        dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n183) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U205 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n42), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n40), .A(
        dp_ex_stage_alu_shifter_srl_41_n183), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n95) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U204 ( .A1(dp_ex_stage_alu_n76), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(
        dp_ex_stage_alu_shifter_N202), .B2(dp_ex_stage_alu_shifter_srl_41_n18), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n182) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U203 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n31), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n30), .A(
        dp_ex_stage_alu_shifter_srl_41_n182), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n179) );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U202 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n34), .A2(
        dp_ex_stage_alu_shifter_srl_41_n78), .B1(
        dp_ex_stage_alu_shifter_srl_41_n33), .B2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n180) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U201 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n111), .B2(
        dp_ex_stage_alu_shifter_srl_41_n114), .C1(
        dp_ex_stage_alu_shifter_srl_41_n154), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n178), .ZN(dp_ex_stage_alu_shifter_N137) );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U200 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n36), .A2(
        dp_ex_stage_alu_shifter_srl_41_n78), .B1(
        dp_ex_stage_alu_shifter_srl_41_n35), .B2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n177) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U199 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n79), .B2(dp_ex_stage_alu_n231), .C1(
        dp_ex_stage_alu_shifter_srl_41_n77), .C2(
        dp_ex_stage_alu_shifter_srl_41_n37), .A(
        dp_ex_stage_alu_shifter_srl_41_n177), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n130) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U198 ( .A1(dp_ex_stage_muxA_out[27]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_muxA_out[26]), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n176) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U197 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n119), .B2(
        dp_ex_stage_alu_shifter_srl_41_n74), .C1(
        dp_ex_stage_alu_shifter_srl_41_n21), .C2(
        dp_ex_stage_alu_shifter_srl_41_n52), .A(
        dp_ex_stage_alu_shifter_srl_41_n176), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n142) );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U196 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n76), .A2(
        dp_ex_stage_alu_shifter_srl_41_n75), .B1(
        dp_ex_stage_alu_shifter_srl_41_n78), .B2(
        dp_ex_stage_alu_shifter_srl_41_n53), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n126) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U195 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n142), .A2(
        dp_ex_stage_alu_shifter_srl_41_n82), .B1(
        dp_ex_stage_alu_shifter_srl_41_n126), .B2(
        dp_ex_stage_alu_shifter_srl_41_n137), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n135) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U194 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n41), .A2(
        dp_ex_stage_alu_shifter_srl_41_n20), .B1(
        dp_ex_stage_alu_shifter_srl_41_n39), .B2(
        dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n175) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U193 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n44), .C1(
        dp_ex_stage_alu_shifter_srl_41_n21), .C2(
        dp_ex_stage_alu_shifter_srl_41_n43), .A(
        dp_ex_stage_alu_shifter_srl_41_n175), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n106) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U192 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n20), .A2(dp_ex_stage_muxA_out[19]), 
        .B1(dp_ex_stage_alu_shifter_srl_41_n18), .B2(dp_ex_stage_muxA_out[18]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n174) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U191 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n119), .B2(
        dp_ex_stage_alu_shifter_srl_41_n46), .C1(
        dp_ex_stage_alu_shifter_srl_41_n69), .C2(
        dp_ex_stage_alu_shifter_srl_41_n22), .A(
        dp_ex_stage_alu_shifter_srl_41_n174), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n107) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U190 ( .A1(dp_ex_stage_muxA_out[23]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_alu_n240), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n173) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U189 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n119), .B2(
        dp_ex_stage_alu_shifter_srl_41_n49), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n48), .A(
        dp_ex_stage_alu_shifter_srl_41_n173), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n143) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U188 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n80), .A2(
        dp_ex_stage_alu_shifter_srl_41_n106), .B1(
        dp_ex_stage_alu_shifter_srl_41_n88), .B2(
        dp_ex_stage_alu_shifter_srl_41_n107), .C1(
        dp_ex_stage_alu_shifter_srl_41_n90), .C2(
        dp_ex_stage_alu_shifter_srl_41_n143), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n172) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U187 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n130), .B2(
        dp_ex_stage_alu_shifter_srl_41_n84), .C1(
        dp_ex_stage_alu_shifter_srl_41_n135), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n172), .ZN(dp_ex_stage_alu_shifter_N147) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U186 ( .A1(dp_ex_stage_alu_n38), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(
        dp_ex_stage_alu_shifter_srl_41_n41), .B2(
        dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n171) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U185 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n45), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n44), .A(
        dp_ex_stage_alu_shifter_srl_41_n171), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n101) );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U184 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n38), .A2(
        dp_ex_stage_alu_shifter_srl_41_n78), .B1(
        dp_ex_stage_alu_shifter_srl_41_n36), .B2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n170) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U183 ( .A1(dp_ex_stage_muxA_out[24]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_muxA_out[23]), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n169) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U182 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n119), .B2(
        dp_ex_stage_alu_shifter_srl_41_n50), .C1(
        dp_ex_stage_alu_shifter_srl_41_n21), .C2(
        dp_ex_stage_alu_shifter_srl_41_n49), .A(
        dp_ex_stage_alu_shifter_srl_41_n169), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n141) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U181 ( .A1(dp_ex_stage_alu_n240), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n79), .B1(dp_ex_stage_muxA_out[21]), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n77), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n168) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U180 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n69), .B2(
        dp_ex_stage_alu_shifter_srl_41_n78), .C1(
        dp_ex_stage_alu_shifter_srl_41_n68), .C2(
        dp_ex_stage_alu_shifter_srl_41_n76), .A(
        dp_ex_stage_alu_shifter_srl_41_n168), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n102) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U179 ( .A1(dp_ex_stage_alu_n1), .A2(
        dp_ex_stage_alu_shifter_srl_41_n19), .B1(dp_ex_stage_muxA_out[27]), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n167) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U178 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n53), .A2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n125) );
  MUX2_X1 dp_ex_stage_alu_shifter_srl_41_U177 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n139), .B(
        dp_ex_stage_alu_shifter_srl_41_n125), .S(dp_ex_stage_alu_n49), .Z(
        dp_ex_stage_alu_shifter_srl_41_n150) );
  NOR3_X1 dp_ex_stage_alu_shifter_srl_41_U176 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n29), .A2(dp_ex_stage_alu_n31), .A3(
        dp_ex_stage_alu_shifter_srl_41_n73), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n166) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U175 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n90), .B2(
        dp_ex_stage_alu_shifter_srl_41_n141), .C1(
        dp_ex_stage_alu_shifter_srl_41_n88), .C2(
        dp_ex_stage_alu_shifter_srl_41_n102), .A(
        dp_ex_stage_alu_shifter_srl_41_n166), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n165) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U174 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n64), .B2(
        dp_ex_stage_alu_shifter_srl_41_n114), .C1(
        dp_ex_stage_alu_shifter_srl_41_n118), .C2(
        dp_ex_stage_alu_shifter_srl_41_n84), .A(
        dp_ex_stage_alu_shifter_srl_41_n165), .ZN(dp_ex_stage_alu_shifter_N148) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U173 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n29), .A2(
        dp_ex_stage_alu_shifter_srl_41_n164), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n156) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U172 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n96), .B2(
        dp_ex_stage_alu_shifter_srl_41_n80), .C1(
        dp_ex_stage_alu_shifter_srl_41_n95), .C2(
        dp_ex_stage_alu_shifter_srl_41_n81), .A(
        dp_ex_stage_alu_shifter_srl_41_n2), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n163) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U171 ( .A1(dp_ex_stage_muxA_out[18]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_muxA_out[17]), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n162) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U170 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n119), .B2(
        dp_ex_stage_alu_shifter_srl_41_n69), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n68), .A(
        dp_ex_stage_alu_shifter_srl_41_n162), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n89) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U169 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n39), .A2(
        dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_alu_n231), .B2(
        dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n161) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U168 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n43), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n42), .A(
        dp_ex_stage_alu_shifter_srl_41_n161), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n87) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U167 ( .A1(dp_ex_stage_muxA_out[26]), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_muxA_out[25]), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n160) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U166 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n119), .B2(
        dp_ex_stage_alu_shifter_srl_41_n52), .C1(
        dp_ex_stage_alu_shifter_srl_41_n21), .C2(
        dp_ex_stage_alu_shifter_srl_41_n51), .A(
        dp_ex_stage_alu_shifter_srl_41_n160), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n136) );
  OAI222_X1 dp_ex_stage_alu_shifter_srl_41_U165 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n78), .A2(
        dp_ex_stage_alu_shifter_srl_41_n75), .B1(
        dp_ex_stage_alu_shifter_srl_41_n21), .B2(
        dp_ex_stage_alu_shifter_srl_41_n53), .C1(
        dp_ex_stage_alu_shifter_srl_41_n76), .C2(
        dp_ex_stage_alu_shifter_srl_41_n74), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n133) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U164 ( .A1(dp_ex_stage_alu_n240), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_muxA_out[21]), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n159) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U163 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n119), .B2(
        dp_ex_stage_alu_shifter_srl_41_n48), .C1(
        dp_ex_stage_alu_shifter_srl_41_n21), .C2(
        dp_ex_stage_alu_shifter_srl_41_n47), .A(
        dp_ex_stage_alu_shifter_srl_41_n159), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n91) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U162 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n90), .A2(
        dp_ex_stage_alu_shifter_srl_41_n136), .B1(
        dp_ex_stage_alu_shifter_srl_41_n156), .B2(
        dp_ex_stage_alu_shifter_srl_41_n133), .C1(
        dp_ex_stage_alu_shifter_srl_41_n88), .C2(
        dp_ex_stage_alu_shifter_srl_41_n91), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n158) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U161 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n65), .B2(
        dp_ex_stage_alu_shifter_srl_41_n114), .C1(
        dp_ex_stage_alu_shifter_srl_41_n62), .C2(
        dp_ex_stage_alu_shifter_srl_41_n84), .A(
        dp_ex_stage_alu_shifter_srl_41_n158), .ZN(dp_ex_stage_alu_shifter_N150) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U160 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n90), .A2(
        dp_ex_stage_alu_shifter_srl_41_n142), .B1(
        dp_ex_stage_alu_shifter_srl_41_n156), .B2(
        dp_ex_stage_alu_shifter_srl_41_n126), .C1(
        dp_ex_stage_alu_shifter_srl_41_n88), .C2(
        dp_ex_stage_alu_shifter_srl_41_n143), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n157) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U159 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n66), .B2(
        dp_ex_stage_alu_shifter_srl_41_n114), .C1(
        dp_ex_stage_alu_shifter_srl_41_n63), .C2(
        dp_ex_stage_alu_shifter_srl_41_n84), .A(
        dp_ex_stage_alu_shifter_srl_41_n157), .ZN(dp_ex_stage_alu_shifter_N151) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U158 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n90), .A2(
        dp_ex_stage_alu_shifter_srl_41_n139), .B1(
        dp_ex_stage_alu_shifter_srl_41_n156), .B2(
        dp_ex_stage_alu_shifter_srl_41_n125), .C1(
        dp_ex_stage_alu_shifter_srl_41_n88), .C2(
        dp_ex_stage_alu_shifter_srl_41_n141), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n155) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U157 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n67), .B2(
        dp_ex_stage_alu_shifter_srl_41_n114), .C1(
        dp_ex_stage_alu_shifter_srl_41_n64), .C2(
        dp_ex_stage_alu_shifter_srl_41_n84), .A(
        dp_ex_stage_alu_shifter_srl_41_n155), .ZN(dp_ex_stage_alu_shifter_N152) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U156 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n28), .A2(
        dp_ex_stage_alu_shifter_srl_41_n154), .ZN(dp_ex_stage_alu_shifter_N153) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U155 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n152), .A2(
        dp_ex_stage_alu_shifter_srl_41_n133), .B1(
        dp_ex_stage_alu_shifter_srl_41_n140), .B2(
        dp_ex_stage_alu_shifter_srl_41_n136), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n153) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U154 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n91), .B2(
        dp_ex_stage_alu_shifter_srl_41_n137), .C1(
        dp_ex_stage_alu_shifter_srl_41_n89), .C2(
        dp_ex_stage_alu_shifter_srl_41_n82), .A(
        dp_ex_stage_alu_shifter_srl_41_n71), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n144) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U153 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n27), .A2(
        dp_ex_stage_alu_shifter_srl_41_n144), .ZN(dp_ex_stage_alu_shifter_N154) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U152 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n152), .A2(
        dp_ex_stage_alu_shifter_srl_41_n126), .B1(
        dp_ex_stage_alu_shifter_srl_41_n140), .B2(
        dp_ex_stage_alu_shifter_srl_41_n142), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n151) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U151 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n143), .B2(
        dp_ex_stage_alu_shifter_srl_41_n137), .C1(
        dp_ex_stage_alu_shifter_srl_41_n107), .C2(
        dp_ex_stage_alu_shifter_srl_41_n82), .A(
        dp_ex_stage_alu_shifter_srl_41_n72), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n127) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U150 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n27), .A2(
        dp_ex_stage_alu_shifter_srl_41_n127), .ZN(dp_ex_stage_alu_shifter_N155) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U149 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n102), .A2(
        dp_ex_stage_alu_shifter_srl_41_n82), .B1(
        dp_ex_stage_alu_shifter_srl_41_n141), .B2(
        dp_ex_stage_alu_shifter_srl_41_n137), .C1(
        dp_ex_stage_alu_shifter_srl_41_n150), .C2(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n115) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U148 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n27), .A2(
        dp_ex_stage_alu_shifter_srl_41_n115), .ZN(dp_ex_stage_alu_shifter_N156) );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U147 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n56), .A2(
        dp_ex_stage_alu_shifter_srl_41_n78), .B1(
        dp_ex_stage_alu_shifter_srl_41_n55), .B2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n149) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U146 ( .A1(dp_ex_stage_alu_n44), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_alu_n76), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n148) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U145 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n54), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n31), .A(
        dp_ex_stage_alu_shifter_srl_41_n148), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n146) );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U144 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n35), .A2(
        dp_ex_stage_alu_shifter_srl_41_n78), .B1(
        dp_ex_stage_alu_shifter_srl_41_n34), .B2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n147) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U143 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n79), .B2(
        dp_ex_stage_alu_shifter_srl_41_n37), .C1(
        dp_ex_stage_alu_shifter_srl_41_n77), .C2(dp_ex_stage_alu_n33), .A(
        dp_ex_stage_alu_shifter_srl_41_n147), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n83) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U142 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n90), .A2(
        dp_ex_stage_alu_shifter_srl_41_n87), .B1(
        dp_ex_stage_alu_shifter_srl_41_n81), .B2(
        dp_ex_stage_alu_shifter_srl_41_n146), .C1(
        dp_ex_stage_alu_shifter_srl_41_n88), .C2(
        dp_ex_stage_alu_shifter_srl_41_n58), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n145) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U141 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n108), .B2(
        dp_ex_stage_alu_shifter_srl_41_n114), .C1(
        dp_ex_stage_alu_shifter_srl_41_n144), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n145), .ZN(dp_ex_stage_alu_shifter_N138) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U140 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n27), .A2(
        dp_ex_stage_alu_shifter_srl_41_n112), .ZN(dp_ex_stage_alu_shifter_N157) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U139 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n136), .A2(
        dp_ex_stage_alu_shifter_srl_41_n137), .B1(
        dp_ex_stage_alu_shifter_srl_41_n133), .B2(
        dp_ex_stage_alu_shifter_srl_41_n140), .C1(
        dp_ex_stage_alu_shifter_srl_41_n91), .C2(
        dp_ex_stage_alu_shifter_srl_41_n82), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n109) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U138 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n27), .A2(
        dp_ex_stage_alu_shifter_srl_41_n109), .ZN(dp_ex_stage_alu_shifter_N158) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U137 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n142), .A2(
        dp_ex_stage_alu_shifter_srl_41_n137), .B1(
        dp_ex_stage_alu_shifter_srl_41_n126), .B2(
        dp_ex_stage_alu_shifter_srl_41_n140), .C1(
        dp_ex_stage_alu_shifter_srl_41_n143), .C2(
        dp_ex_stage_alu_shifter_srl_41_n82), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n104) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U136 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n26), .A2(
        dp_ex_stage_alu_shifter_srl_41_n104), .ZN(dp_ex_stage_alu_shifter_N159) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U135 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n26), .A2(
        dp_ex_stage_alu_shifter_srl_41_n99), .ZN(dp_ex_stage_alu_shifter_N160)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U134 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n138), .A2(
        dp_ex_stage_alu_shifter_srl_41_n82), .B1(
        dp_ex_stage_alu_shifter_srl_41_n134), .B2(
        dp_ex_stage_alu_shifter_srl_41_n137), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n93) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U133 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n26), .A2(
        dp_ex_stage_alu_shifter_srl_41_n93), .ZN(dp_ex_stage_alu_shifter_N161)
         );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U132 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n136), .A2(
        dp_ex_stage_alu_shifter_srl_41_n82), .B1(
        dp_ex_stage_alu_shifter_srl_41_n133), .B2(
        dp_ex_stage_alu_shifter_srl_41_n137), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n85) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U131 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n26), .A2(
        dp_ex_stage_alu_shifter_srl_41_n85), .ZN(dp_ex_stage_alu_shifter_N162)
         );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U130 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n26), .A2(
        dp_ex_stage_alu_shifter_srl_41_n135), .ZN(dp_ex_stage_alu_shifter_N163) );
  NOR3_X1 dp_ex_stage_alu_shifter_srl_41_U129 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n73), .A2(
        dp_ex_stage_alu_shifter_srl_41_n28), .A3(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_shifter_N164) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U128 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n134), .A2(
        dp_ex_stage_alu_shifter_srl_41_n81), .ZN(dp_ex_stage_alu_shifter_N165)
         );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U127 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n133), .A2(
        dp_ex_stage_alu_shifter_srl_41_n81), .ZN(dp_ex_stage_alu_shifter_N166)
         );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U126 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n32), .A2(
        dp_ex_stage_alu_shifter_srl_41_n78), .B1(
        dp_ex_stage_alu_shifter_srl_41_n56), .B2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n132) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U125 ( .A1(dp_ex_stage_alu_n69), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_alu_n44), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n131) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U124 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n55), .C1(
        dp_ex_stage_alu_shifter_srl_41_n22), .C2(
        dp_ex_stage_alu_shifter_srl_41_n54), .A(
        dp_ex_stage_alu_shifter_srl_41_n131), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n129) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U123 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n90), .A2(
        dp_ex_stage_alu_shifter_srl_41_n106), .B1(
        dp_ex_stage_alu_shifter_srl_41_n81), .B2(
        dp_ex_stage_alu_shifter_srl_41_n129), .C1(
        dp_ex_stage_alu_shifter_srl_41_n88), .C2(
        dp_ex_stage_alu_shifter_srl_41_n59), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n128) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U122 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n103), .B2(
        dp_ex_stage_alu_shifter_srl_41_n114), .C1(
        dp_ex_stage_alu_shifter_srl_41_n127), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n128), .ZN(dp_ex_stage_alu_shifter_N139) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U121 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n126), .A2(
        dp_ex_stage_alu_shifter_srl_41_n81), .ZN(dp_ex_stage_alu_shifter_N167)
         );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U120 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n81), .A2(
        dp_ex_stage_alu_shifter_srl_41_n125), .ZN(dp_ex_stage_alu_shifter_N168) );
  OAI22_X1 dp_ex_stage_alu_shifter_srl_41_U119 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n33), .A2(
        dp_ex_stage_alu_shifter_srl_41_n78), .B1(
        dp_ex_stage_alu_shifter_srl_41_n32), .B2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n124) );
  AOI22_X1 dp_ex_stage_alu_shifter_srl_41_U118 ( .A1(dp_ex_stage_alu_n52), 
        .A2(dp_ex_stage_alu_shifter_srl_41_n20), .B1(dp_ex_stage_alu_n69), 
        .B2(dp_ex_stage_alu_shifter_srl_41_n18), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n121) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U117 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n1), .B2(
        dp_ex_stage_alu_shifter_srl_41_n56), .C1(
        dp_ex_stage_alu_shifter_srl_41_n21), .C2(
        dp_ex_stage_alu_shifter_srl_41_n55), .A(
        dp_ex_stage_alu_shifter_srl_41_n121), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n117) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U116 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n90), .A2(
        dp_ex_stage_alu_shifter_srl_41_n101), .B1(
        dp_ex_stage_alu_shifter_srl_41_n81), .B2(
        dp_ex_stage_alu_shifter_srl_41_n117), .C1(
        dp_ex_stage_alu_shifter_srl_41_n88), .C2(
        dp_ex_stage_alu_shifter_srl_41_n60), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n116) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U115 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n98), .B2(
        dp_ex_stage_alu_shifter_srl_41_n114), .C1(
        dp_ex_stage_alu_shifter_srl_41_n115), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n116), .ZN(dp_ex_stage_alu_shifter_N140) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U114 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n80), .A2(
        dp_ex_stage_alu_shifter_srl_41_n57), .B1(
        dp_ex_stage_alu_shifter_srl_41_n88), .B2(
        dp_ex_stage_alu_shifter_srl_41_n95), .C1(
        dp_ex_stage_alu_shifter_srl_41_n90), .C2(
        dp_ex_stage_alu_shifter_srl_41_n96), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n113) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U113 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n111), .B2(
        dp_ex_stage_alu_shifter_srl_41_n84), .C1(
        dp_ex_stage_alu_shifter_srl_41_n112), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n113), .ZN(dp_ex_stage_alu_shifter_N141) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U112 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n80), .A2(
        dp_ex_stage_alu_shifter_srl_41_n58), .B1(
        dp_ex_stage_alu_shifter_srl_41_n88), .B2(
        dp_ex_stage_alu_shifter_srl_41_n87), .C1(
        dp_ex_stage_alu_shifter_srl_41_n90), .C2(
        dp_ex_stage_alu_shifter_srl_41_n89), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n110) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U111 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n108), .B2(
        dp_ex_stage_alu_shifter_srl_41_n84), .C1(
        dp_ex_stage_alu_shifter_srl_41_n109), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n110), .ZN(dp_ex_stage_alu_shifter_N142) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U110 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n80), .A2(
        dp_ex_stage_alu_shifter_srl_41_n59), .B1(
        dp_ex_stage_alu_shifter_srl_41_n88), .B2(
        dp_ex_stage_alu_shifter_srl_41_n106), .C1(
        dp_ex_stage_alu_shifter_srl_41_n90), .C2(
        dp_ex_stage_alu_shifter_srl_41_n107), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n105) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U109 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n103), .B2(
        dp_ex_stage_alu_shifter_srl_41_n84), .C1(
        dp_ex_stage_alu_shifter_srl_41_n104), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n105), .ZN(dp_ex_stage_alu_shifter_N143) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U108 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n80), .A2(
        dp_ex_stage_alu_shifter_srl_41_n60), .B1(
        dp_ex_stage_alu_shifter_srl_41_n88), .B2(
        dp_ex_stage_alu_shifter_srl_41_n101), .C1(
        dp_ex_stage_alu_shifter_srl_41_n90), .C2(
        dp_ex_stage_alu_shifter_srl_41_n102), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n100) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U107 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n98), .B2(
        dp_ex_stage_alu_shifter_srl_41_n84), .C1(
        dp_ex_stage_alu_shifter_srl_41_n99), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n100), .ZN(dp_ex_stage_alu_shifter_N144) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U106 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n80), .A2(
        dp_ex_stage_alu_shifter_srl_41_n95), .B1(
        dp_ex_stage_alu_shifter_srl_41_n88), .B2(
        dp_ex_stage_alu_shifter_srl_41_n96), .C1(
        dp_ex_stage_alu_shifter_srl_41_n90), .C2(
        dp_ex_stage_alu_shifter_srl_41_n97), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n94) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U105 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n92), .B2(
        dp_ex_stage_alu_shifter_srl_41_n84), .C1(
        dp_ex_stage_alu_shifter_srl_41_n93), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n94), .ZN(dp_ex_stage_alu_shifter_N145)
         );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U104 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n80), .A2(
        dp_ex_stage_alu_shifter_srl_41_n87), .B1(
        dp_ex_stage_alu_shifter_srl_41_n88), .B2(
        dp_ex_stage_alu_shifter_srl_41_n89), .C1(
        dp_ex_stage_alu_shifter_srl_41_n90), .C2(
        dp_ex_stage_alu_shifter_srl_41_n91), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n86) );
  OAI221_X1 dp_ex_stage_alu_shifter_srl_41_U103 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n83), .B2(
        dp_ex_stage_alu_shifter_srl_41_n84), .C1(
        dp_ex_stage_alu_shifter_srl_41_n85), .C2(
        dp_ex_stage_alu_shifter_srl_41_n29), .A(
        dp_ex_stage_alu_shifter_srl_41_n86), .ZN(dp_ex_stage_alu_shifter_N146)
         );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U102 ( .A(dp_ex_stage_muxA_out[31]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n53) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U101 ( .A(dp_ex_stage_alu_n1), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n52) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U100 ( .A(dp_ex_stage_muxA_out[27]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n51) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U99 ( .A(dp_ex_stage_muxA_out[26]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n50) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U98 ( .A(dp_ex_stage_muxA_out[25]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n49) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U97 ( .A(dp_ex_stage_muxA_out[24]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n48) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U96 ( .A(dp_ex_stage_muxA_out[23]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n47) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U95 ( .A(dp_ex_stage_muxA_out[21]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n46) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U94 ( .A(dp_ex_stage_muxA_out[18]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n45) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U93 ( .A(dp_ex_stage_muxA_out[17]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n44) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U92 ( .A(dp_ex_stage_alu_n38), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n43) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U91 ( .A(dp_ex_stage_alu_n29), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n42) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U90 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n42), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n41) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U89 ( .A(dp_ex_stage_muxA_out[14]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n40) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U88 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n40), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n39) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U87 ( .A(dp_ex_stage_muxA_out[12]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n38) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U86 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n38), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n37) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U85 ( .A(dp_ex_stage_alu_n33), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n36) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U84 ( .A(dp_ex_stage_alu_n74), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n35) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U83 ( .A(dp_ex_stage_alu_n72), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n34) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U82 ( .A(dp_ex_stage_alu_n71), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n33) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U81 ( .A(dp_ex_stage_alu_n34), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n32) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U80 ( .A(dp_ex_stage_alu_n69), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n31) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U79 ( .A(dp_ex_stage_alu_n44), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n30) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U78 ( .A(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n25) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U77 ( .A(dp_ex_stage_alu_n49), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n24) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U76 ( .A(dp_ex_stage_alu_n45), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n23) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U75 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n23), .A2(dp_ex_stage_alu_n46), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n122) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U74 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n163), .ZN(dp_ex_stage_alu_shifter_N149) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U73 ( .A(dp_ex_stage_alu_n52), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n54) );
  BUF_X2 dp_ex_stage_alu_shifter_srl_41_U72 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n122), .Z(
        dp_ex_stage_alu_shifter_srl_41_n20) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_srl_41_U71 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n122), .Z(
        dp_ex_stage_alu_shifter_srl_41_n19) );
  NOR2_X1 dp_ex_stage_alu_shifter_srl_41_U70 ( .A1(dp_ex_stage_alu_n45), .A2(
        dp_ex_stage_alu_n46), .ZN(dp_ex_stage_alu_shifter_srl_41_n123) );
  BUF_X2 dp_ex_stage_alu_shifter_srl_41_U69 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n123), .Z(
        dp_ex_stage_alu_shifter_srl_41_n18) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U68 ( .A(dp_ex_stage_alu_n78), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n56) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U67 ( .A(dp_ex_stage_alu_n70), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n55) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U66 ( .A(dp_ex_stage_muxA_out[29]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n74) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U65 ( .A(dp_ex_stage_muxA_out[19]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n68) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U64 ( .A(dp_ex_stage_muxA_out[30]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n75) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U63 ( .A(dp_ex_stage_muxA_out[20]), 
        .ZN(dp_ex_stage_alu_shifter_srl_41_n69) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U62 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n92), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n57) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U61 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n150), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n73) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U60 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n107), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n66) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U59 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n83), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n58) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U58 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n119), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n79) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U57 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n184), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n70) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U56 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n151), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n72) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U55 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n153), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n71) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U54 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n89), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n65) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U53 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n102), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n67) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U52 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n87), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n62) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U51 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n106), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n63) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U50 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n101), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n64) );
  BUF_X1 dp_ex_stage_alu_shifter_srl_41_U49 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n120), .Z(
        dp_ex_stage_alu_shifter_srl_41_n22) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U48 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n118), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n60) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U47 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n130), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n59) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U46 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n120), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n77) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U45 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n114), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n80) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U44 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n164), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n82) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U43 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n28), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n29) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U42 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n84), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n81) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_srl_41_U41 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_srl_41_n27)
         );
  CLKBUF_X1 dp_ex_stage_alu_shifter_srl_41_U40 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_srl_41_n26)
         );
  INV_X2 dp_ex_stage_alu_shifter_srl_41_U39 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n123), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n76) );
  INV_X2 dp_ex_stage_alu_shifter_srl_41_U38 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n19), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n78) );
  NAND3_X1 dp_ex_stage_alu_shifter_srl_41_U37 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n16), .A2(
        dp_ex_stage_alu_shifter_srl_41_n17), .A3(
        dp_ex_stage_alu_shifter_srl_41_n188), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n97) );
  OR2_X1 dp_ex_stage_alu_shifter_srl_41_U36 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n69), .A2(
        dp_ex_stage_alu_shifter_srl_41_n76), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n17) );
  OR2_X1 dp_ex_stage_alu_shifter_srl_41_U35 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n78), .A2(
        dp_ex_stage_alu_shifter_srl_41_n46), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n16) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U34 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n88), .A2(
        dp_ex_stage_alu_shifter_srl_41_n97), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n15) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U33 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n156), .A2(
        dp_ex_stage_alu_shifter_srl_41_n134), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n14) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U32 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n90), .A2(
        dp_ex_stage_alu_shifter_srl_41_n138), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n13) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U31 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n77), .A2(dp_ex_stage_alu_n74), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n12) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U30 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n79), .A2(dp_ex_stage_alu_n33), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n11) );
  AND3_X1 dp_ex_stage_alu_shifter_srl_41_U29 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n8), .A2(
        dp_ex_stage_alu_shifter_srl_41_n9), .A3(
        dp_ex_stage_alu_shifter_srl_41_n10), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n178) );
  NAND2_X1 dp_ex_stage_alu_shifter_srl_41_U28 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n88), .A2(
        dp_ex_stage_alu_shifter_srl_41_n57), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n10) );
  NAND2_X1 dp_ex_stage_alu_shifter_srl_41_U27 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n81), .A2(
        dp_ex_stage_alu_shifter_srl_41_n179), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n9) );
  NAND2_X1 dp_ex_stage_alu_shifter_srl_41_U26 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n90), .A2(
        dp_ex_stage_alu_shifter_srl_41_n95), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n8) );
  CLKBUF_X3 dp_ex_stage_alu_shifter_srl_41_U25 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n120), .Z(
        dp_ex_stage_alu_shifter_srl_41_n21) );
  NAND3_X1 dp_ex_stage_alu_shifter_srl_41_U24 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n6), .A2(
        dp_ex_stage_alu_shifter_srl_41_n7), .A3(
        dp_ex_stage_alu_shifter_srl_41_n186), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n134) );
  OR2_X1 dp_ex_stage_alu_shifter_srl_41_U23 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n21), .A2(
        dp_ex_stage_alu_shifter_srl_41_n75), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n7) );
  OR2_X1 dp_ex_stage_alu_shifter_srl_41_U22 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n119), .A2(
        dp_ex_stage_alu_shifter_srl_41_n53), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n6) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U21 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n139), .A2(
        dp_ex_stage_alu_shifter_srl_41_n137), .B1(
        dp_ex_stage_alu_shifter_srl_41_n125), .B2(
        dp_ex_stage_alu_shifter_srl_41_n140), .C1(
        dp_ex_stage_alu_shifter_srl_41_n141), .C2(
        dp_ex_stage_alu_shifter_srl_41_n82), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n99) );
  NAND3_X1 dp_ex_stage_alu_shifter_srl_41_U20 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n4), .A2(
        dp_ex_stage_alu_shifter_srl_41_n5), .A3(
        dp_ex_stage_alu_shifter_srl_41_n167), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n139) );
  OR2_X1 dp_ex_stage_alu_shifter_srl_41_U19 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n21), .A2(
        dp_ex_stage_alu_shifter_srl_41_n74), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n5) );
  OR2_X1 dp_ex_stage_alu_shifter_srl_41_U18 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n119), .A2(
        dp_ex_stage_alu_shifter_srl_41_n75), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n4) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U17 ( .A(dp_ex_stage_alu_n45), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n3) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U16 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n181), .A2(
        dp_ex_stage_alu_shifter_srl_41_n24), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n88) );
  AOI222_X1 dp_ex_stage_alu_shifter_srl_41_U15 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n138), .A2(
        dp_ex_stage_alu_shifter_srl_41_n137), .B1(
        dp_ex_stage_alu_shifter_srl_41_n134), .B2(
        dp_ex_stage_alu_shifter_srl_41_n140), .C1(
        dp_ex_stage_alu_shifter_srl_41_n97), .C2(
        dp_ex_stage_alu_shifter_srl_41_n82), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n112) );
  AND2_X1 dp_ex_stage_alu_shifter_srl_41_U14 ( .A1(dp_ex_stage_alu_n49), .A2(
        dp_ex_stage_alu_shifter_srl_41_n181), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n90) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U13 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n79), .B2(
        dp_ex_stage_alu_shifter_srl_41_n39), .C1(
        dp_ex_stage_alu_shifter_srl_41_n77), .C2(dp_ex_stage_alu_n231), .A(
        dp_ex_stage_alu_shifter_srl_41_n170), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n118) );
  NAND2_X2 dp_ex_stage_alu_shifter_srl_41_U12 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n82), .A2(
        dp_ex_stage_alu_shifter_srl_41_n29), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n84) );
  OR3_X1 dp_ex_stage_alu_shifter_srl_41_U11 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n13), .A2(
        dp_ex_stage_alu_shifter_srl_41_n14), .A3(
        dp_ex_stage_alu_shifter_srl_41_n15), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n2) );
  BUF_X1 dp_ex_stage_alu_shifter_srl_41_U10 ( .A(dp_ex_stage_alu_shifter_n116), 
        .Z(dp_ex_stage_alu_shifter_srl_41_n28) );
  NAND2_X1 dp_ex_stage_alu_shifter_srl_41_U9 ( .A1(dp_ex_stage_alu_n46), .A2(
        dp_ex_stage_alu_n45), .ZN(dp_ex_stage_alu_shifter_srl_41_n119) );
  INV_X1 dp_ex_stage_alu_shifter_srl_41_U8 ( .A(
        dp_ex_stage_alu_shifter_srl_41_n79), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n1) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U7 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n79), .B2(dp_ex_stage_alu_n71), .C1(
        dp_ex_stage_alu_shifter_srl_41_n77), .C2(dp_ex_stage_alu_n34), .A(
        dp_ex_stage_alu_shifter_srl_41_n149), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n108) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U6 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n79), .B2(dp_ex_stage_alu_n74), .C1(
        dp_ex_stage_alu_shifter_srl_41_n77), .C2(dp_ex_stage_alu_n72), .A(
        dp_ex_stage_alu_shifter_srl_41_n124), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n98) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U5 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n79), .B2(dp_ex_stage_alu_n34), .C1(
        dp_ex_stage_alu_shifter_srl_41_n77), .C2(dp_ex_stage_alu_n78), .A(
        dp_ex_stage_alu_shifter_srl_41_n189), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n111) );
  AOI221_X1 dp_ex_stage_alu_shifter_srl_41_U4 ( .B1(
        dp_ex_stage_alu_shifter_srl_41_n79), .B2(dp_ex_stage_alu_n72), .C1(
        dp_ex_stage_alu_shifter_srl_41_n77), .C2(dp_ex_stage_alu_n71), .A(
        dp_ex_stage_alu_shifter_srl_41_n132), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n103) );
  NOR3_X1 dp_ex_stage_alu_shifter_srl_41_U3 ( .A1(
        dp_ex_stage_alu_shifter_srl_41_n11), .A2(
        dp_ex_stage_alu_shifter_srl_41_n12), .A3(
        dp_ex_stage_alu_shifter_srl_41_n180), .ZN(
        dp_ex_stage_alu_shifter_srl_41_n92) );
  OAI22_X1 dp_ex_stage_alu_shifter_sra_39_U225 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n47), .A2(
        dp_ex_stage_alu_shifter_sra_39_n10), .B1(
        dp_ex_stage_alu_shifter_sra_39_n46), .B2(
        dp_ex_stage_alu_shifter_sra_39_n13), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n193) );
  NOR2_X1 dp_ex_stage_alu_shifter_sra_39_U224 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n17), .A2(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n131) );
  NAND2_X1 dp_ex_stage_alu_shifter_sra_39_U223 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n131), .A2(
        dp_ex_stage_alu_shifter_sra_39_n21), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n107) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U222 ( .A1(dp_ex_stage_alu_n240), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n113), .B1(
        dp_ex_stage_alu_shifter_sra_39_n37), .B2(
        dp_ex_stage_alu_shifter_sra_39_n114), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n192) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U221 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n10), .B2(
        dp_ex_stage_alu_shifter_sra_39_n36), .C1(
        dp_ex_stage_alu_shifter_sra_39_n63), .C2(
        dp_ex_stage_alu_shifter_sra_39_n12), .A(
        dp_ex_stage_alu_shifter_sra_39_n192), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n91) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U220 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n32), .A2(
        dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_alu_n38), .B2(
        dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n191) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U219 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n34), .C1(
        dp_ex_stage_alu_shifter_sra_39_n62), .C2(
        dp_ex_stage_alu_shifter_sra_39_n74), .A(
        dp_ex_stage_alu_shifter_sra_39_n191), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n90) );
  AND2_X1 dp_ex_stage_alu_shifter_sra_39_U218 ( .A1(dp_ex_stage_alu_n49), .A2(
        dp_ex_stage_alu_n31), .ZN(dp_ex_stage_alu_shifter_sra_39_n155) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U217 ( .A1(dp_ex_stage_muxA_out[29]), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_alu_n1), .B2(
        dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n190) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U216 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n70), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n45), .A(
        dp_ex_stage_alu_shifter_sra_39_n190), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n134) );
  AND2_X1 dp_ex_stage_alu_shifter_sra_39_U215 ( .A1(dp_ex_stage_alu_n31), .A2(
        dp_ex_stage_alu_shifter_sra_39_n17), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n141) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U214 ( .A1(dp_ex_stage_muxA_out[25]), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n14), .B1(dp_ex_stage_muxA_out[24]), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n189) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U213 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n155), .A2(
        dp_ex_stage_alu_shifter_sra_39_n134), .B1(
        dp_ex_stage_alu_shifter_sra_39_n141), .B2(
        dp_ex_stage_alu_shifter_sra_39_n135), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n188) );
  AND2_X1 dp_ex_stage_alu_shifter_sra_39_U212 ( .A1(dp_ex_stage_alu_n31), .A2(
        dp_ex_stage_alu_shifter_sra_39_n22), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n185) );
  AND2_X1 dp_ex_stage_alu_shifter_sra_39_U211 ( .A1(dp_ex_stage_alu_n49), .A2(
        dp_ex_stage_alu_shifter_sra_39_n185), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n85) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U210 ( .A1(dp_ex_stage_alu_n231), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n73), .B1(
        dp_ex_stage_alu_shifter_sra_39_n30), .B2(
        dp_ex_stage_alu_shifter_sra_39_n15), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n187) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U209 ( .A1(dp_ex_stage_alu_n76), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n14), .B1(
        dp_ex_stage_alu_shifter_N202), .B2(dp_ex_stage_alu_shifter_sra_39_n75), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n186) );
  OAI22_X1 dp_ex_stage_alu_shifter_sra_39_U208 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n27), .A2(
        dp_ex_stage_alu_shifter_sra_39_n10), .B1(
        dp_ex_stage_alu_shifter_sra_39_n26), .B2(
        dp_ex_stage_alu_shifter_sra_39_n13), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n184) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U207 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n85), .A2(
        dp_ex_stage_alu_shifter_sra_39_n53), .B1(
        dp_ex_stage_alu_shifter_sra_39_n77), .B2(
        dp_ex_stage_alu_shifter_sra_39_n183), .C1(
        dp_ex_stage_alu_shifter_sra_39_n83), .C2(
        dp_ex_stage_alu_shifter_sra_39_n49), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n182) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U206 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n104), .B2(
        dp_ex_stage_alu_shifter_sra_39_n107), .C1(
        dp_ex_stage_alu_shifter_sra_39_n158), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n182), .ZN(dp_ex_stage_alu_shifter_N105) );
  OAI22_X1 dp_ex_stage_alu_shifter_sra_39_U205 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n29), .A2(
        dp_ex_stage_alu_shifter_sra_39_n10), .B1(
        dp_ex_stage_alu_shifter_sra_39_n28), .B2(
        dp_ex_stage_alu_shifter_sra_39_n13), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n181) );
  MUX2_X1 dp_ex_stage_alu_shifter_sra_39_U204 ( .A(dp_ex_stage_muxA_out[30]), 
        .B(dp_ex_stage_alu_shifter_N136), .S(
        dp_ex_stage_alu_shifter_sra_39_n12), .Z(
        dp_ex_stage_alu_shifter_sra_39_n142) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U203 ( .A1(dp_ex_stage_muxA_out[27]), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_muxA_out[26]), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n180) );
  NAND2_X1 dp_ex_stage_alu_shifter_sra_39_U202 ( .A1(
        dp_ex_stage_alu_shifter_N136), .A2(dp_ex_stage_alu_n31), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n154) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U201 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n142), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n138), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n71), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n129) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U200 ( .A1(dp_ex_stage_alu_n29), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n14), .B1(dp_ex_stage_muxA_out[14]), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n15), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n179) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U199 ( .A1(dp_ex_stage_muxA_out[20]), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n113), .B1(
        dp_ex_stage_alu_shifter_sra_39_n35), .B2(
        dp_ex_stage_alu_shifter_sra_39_n114), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n178) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U198 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n62), .B2(
        dp_ex_stage_alu_shifter_sra_39_n10), .C1(
        dp_ex_stage_alu_shifter_sra_39_n34), .C2(
        dp_ex_stage_alu_shifter_sra_39_n12), .A(
        dp_ex_stage_alu_shifter_sra_39_n178), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n100) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U197 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n37), .A2(
        dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_alu_n240), .B2(
        dp_ex_stage_alu_shifter_sra_39_n15), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n177) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U196 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n39), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n40), .A(
        dp_ex_stage_alu_shifter_sra_39_n177), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n139) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U195 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n57), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n100), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n139), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n176) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U194 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n123), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n129), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n176), .ZN(dp_ex_stage_alu_shifter_N115) );
  OAI22_X1 dp_ex_stage_alu_shifter_sra_39_U193 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n31), .A2(
        dp_ex_stage_alu_shifter_sra_39_n10), .B1(
        dp_ex_stage_alu_shifter_sra_39_n29), .B2(
        dp_ex_stage_alu_shifter_sra_39_n13), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n175) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U192 ( .A1(dp_ex_stage_alu_n1), .A2(
        dp_ex_stage_alu_shifter_sra_39_n14), .B1(dp_ex_stage_muxA_out[27]), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n174) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U191 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n68), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n70), .A(
        dp_ex_stage_alu_shifter_sra_39_n174), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n136) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U190 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n17), .B2(
        dp_ex_stage_alu_shifter_sra_39_n45), .A(
        dp_ex_stage_alu_shifter_sra_39_n154), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n162) );
  AOI21_X1 dp_ex_stage_alu_shifter_sra_39_U189 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n136), .B2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n162), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n128) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U188 ( .A1(dp_ex_stage_alu_n38), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_alu_n29), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n173) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U187 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n35), .A2(
        dp_ex_stage_alu_shifter_sra_39_n113), .B1(dp_ex_stage_alu_n240), .B2(
        dp_ex_stage_alu_shifter_sra_39_n114), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n172) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U186 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n63), .B2(
        dp_ex_stage_alu_shifter_sra_39_n10), .C1(
        dp_ex_stage_alu_shifter_sra_39_n62), .C2(
        dp_ex_stage_alu_shifter_sra_39_n13), .A(
        dp_ex_stage_alu_shifter_sra_39_n172), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n96) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U185 ( .A1(dp_ex_stage_muxA_out[24]), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n14), .B1(
        dp_ex_stage_alu_shifter_sra_39_n37), .B2(
        dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n171) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U184 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n95), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n96), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n137), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n170) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U183 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n111), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n128), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n170), .ZN(dp_ex_stage_alu_shifter_N116) );
  AOI21_X1 dp_ex_stage_alu_shifter_sra_39_U182 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n7), .B2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n162), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n127) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U181 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n90), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n91), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n135), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n169) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U180 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n168), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n127), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n169), .ZN(dp_ex_stage_alu_shifter_N117) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U179 ( .A1(dp_ex_stage_muxA_out[14]), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n14), .B1(dp_ex_stage_alu_n231), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n15), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n167) );
  OAI222_X1 dp_ex_stage_alu_shifter_sra_39_U178 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n13), .A2(
        dp_ex_stage_alu_shifter_sra_39_n68), .B1(
        dp_ex_stage_alu_shifter_sra_39_n10), .B2(
        dp_ex_stage_alu_shifter_sra_39_n70), .C1(
        dp_ex_stage_alu_shifter_sra_39_n3), .C2(
        dp_ex_stage_alu_shifter_sra_39_n45), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n130) );
  AOI21_X1 dp_ex_stage_alu_shifter_sra_39_U177 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n130), .B2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n162), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n126) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U176 ( .A1(dp_ex_stage_muxA_out[18]), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n14), .B1(
        dp_ex_stage_alu_shifter_sra_39_n32), .B2(
        dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n166) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U175 ( .A1(dp_ex_stage_alu_n240), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n14), .B1(
        dp_ex_stage_alu_shifter_sra_39_n35), .B2(
        dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n165) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U174 ( .A1(dp_ex_stage_muxA_out[26]), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_muxA_out[25]), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n15), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n164) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U173 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n42), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n43), .A(
        dp_ex_stage_alu_shifter_sra_39_n164), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n132) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U172 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n84), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n86), .C1(
        dp_ex_stage_alu_shifter_sra_39_n132), .C2(
        dp_ex_stage_alu_shifter_sra_39_n85), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n163) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U171 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n151), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n126), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n163), .ZN(dp_ex_stage_alu_shifter_N118) );
  AOI21_X1 dp_ex_stage_alu_shifter_sra_39_U170 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n142), .B2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n162), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n118) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U169 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n100), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n139), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n138), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n161) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U168 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n160), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n118), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n161), .ZN(dp_ex_stage_alu_shifter_N119) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U167 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n85), .B2(
        dp_ex_stage_alu_shifter_sra_39_n136), .C1(
        dp_ex_stage_alu_shifter_sra_39_n83), .C2(
        dp_ex_stage_alu_shifter_sra_39_n137), .A(
        dp_ex_stage_alu_shifter_sra_39_n72), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n159) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U166 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n61), .B2(
        dp_ex_stage_alu_shifter_sra_39_n107), .C1(
        dp_ex_stage_alu_shifter_sra_39_n59), .C2(
        dp_ex_stage_alu_shifter_sra_39_n80), .A(
        dp_ex_stage_alu_shifter_sra_39_n159), .ZN(dp_ex_stage_alu_shifter_N120) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U165 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n20), .B2(
        dp_ex_stage_alu_shifter_sra_39_n158), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N121) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U164 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n155), .A2(
        dp_ex_stage_alu_shifter_sra_39_n130), .B1(
        dp_ex_stage_alu_shifter_sra_39_n132), .B2(
        dp_ex_stage_alu_shifter_sra_39_n141), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n157) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U163 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n20), .B2(
        dp_ex_stage_alu_shifter_sra_39_n146), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N122) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U162 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n131), .A2(
        dp_ex_stage_alu_shifter_sra_39_n139), .B1(
        dp_ex_stage_alu_shifter_sra_39_n133), .B2(
        dp_ex_stage_alu_shifter_sra_39_n100), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n156) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U161 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n142), .B2(
        dp_ex_stage_alu_shifter_sra_39_n155), .C1(
        dp_ex_stage_alu_shifter_sra_39_n138), .C2(
        dp_ex_stage_alu_shifter_sra_39_n141), .A(
        dp_ex_stage_alu_shifter_sra_39_n60), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n120) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U160 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n20), .B2(
        dp_ex_stage_alu_shifter_sra_39_n120), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N123) );
  NOR2_X1 dp_ex_stage_alu_shifter_sra_39_U159 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n154), .A2(
        dp_ex_stage_alu_shifter_sra_39_n17), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n143) );
  AOI21_X1 dp_ex_stage_alu_shifter_sra_39_U158 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n141), .B2(
        dp_ex_stage_alu_shifter_sra_39_n136), .A(
        dp_ex_stage_alu_shifter_sra_39_n143), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n153) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U157 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n19), .B2(
        dp_ex_stage_alu_shifter_sra_39_n108), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N124) );
  OAI22_X1 dp_ex_stage_alu_shifter_sra_39_U156 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n48), .A2(
        dp_ex_stage_alu_shifter_sra_39_n10), .B1(
        dp_ex_stage_alu_shifter_sra_39_n47), .B2(
        dp_ex_stage_alu_shifter_sra_39_n12), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n152) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U155 ( .A1(dp_ex_stage_alu_n44), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_alu_n76), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n150) );
  OAI22_X1 dp_ex_stage_alu_shifter_sra_39_U154 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n28), .A2(
        dp_ex_stage_alu_shifter_sra_39_n10), .B1(
        dp_ex_stage_alu_shifter_sra_39_n27), .B2(
        dp_ex_stage_alu_shifter_sra_39_n13), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n149) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U153 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n85), .A2(
        dp_ex_stage_alu_shifter_sra_39_n55), .B1(
        dp_ex_stage_alu_shifter_sra_39_n77), .B2(
        dp_ex_stage_alu_shifter_sra_39_n148), .C1(
        dp_ex_stage_alu_shifter_sra_39_n83), .C2(
        dp_ex_stage_alu_shifter_sra_39_n50), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n147) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U152 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n101), .B2(
        dp_ex_stage_alu_shifter_sra_39_n107), .C1(
        dp_ex_stage_alu_shifter_sra_39_n146), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n147), .ZN(dp_ex_stage_alu_shifter_N106) );
  AOI21_X1 dp_ex_stage_alu_shifter_sra_39_U151 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n141), .B2(
        dp_ex_stage_alu_shifter_sra_39_n134), .A(
        dp_ex_stage_alu_shifter_sra_39_n143), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n145) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U150 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n19), .B2(
        dp_ex_stage_alu_shifter_sra_39_n105), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N125) );
  AOI21_X1 dp_ex_stage_alu_shifter_sra_39_U149 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n141), .B2(
        dp_ex_stage_alu_shifter_sra_39_n130), .A(
        dp_ex_stage_alu_shifter_sra_39_n143), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n144) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U148 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n19), .B2(
        dp_ex_stage_alu_shifter_sra_39_n102), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N126) );
  AOI21_X1 dp_ex_stage_alu_shifter_sra_39_U147 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n141), .B2(
        dp_ex_stage_alu_shifter_sra_39_n142), .A(
        dp_ex_stage_alu_shifter_sra_39_n143), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n140) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U146 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n19), .B2(
        dp_ex_stage_alu_shifter_sra_39_n98), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N127) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U145 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n19), .B2(
        dp_ex_stage_alu_shifter_sra_39_n93), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N128) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U144 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n19), .B2(
        dp_ex_stage_alu_shifter_sra_39_n88), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N129) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U143 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n19), .B2(
        dp_ex_stage_alu_shifter_sra_39_n81), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N130) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U142 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n18), .B2(
        dp_ex_stage_alu_shifter_sra_39_n129), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N131) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U141 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n18), .B2(
        dp_ex_stage_alu_shifter_sra_39_n128), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N132) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U140 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n18), .B2(
        dp_ex_stage_alu_shifter_sra_39_n127), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N133) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U139 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n18), .B2(
        dp_ex_stage_alu_shifter_sra_39_n126), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N134) );
  OAI22_X1 dp_ex_stage_alu_shifter_sra_39_U138 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n25), .A2(
        dp_ex_stage_alu_shifter_sra_39_n10), .B1(
        dp_ex_stage_alu_shifter_sra_39_n48), .B2(
        dp_ex_stage_alu_shifter_sra_39_n12), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n125) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U137 ( .A1(dp_ex_stage_alu_n69), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_alu_n44), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n124) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U136 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n85), .A2(
        dp_ex_stage_alu_shifter_sra_39_n57), .B1(
        dp_ex_stage_alu_shifter_sra_39_n77), .B2(
        dp_ex_stage_alu_shifter_sra_39_n122), .C1(
        dp_ex_stage_alu_shifter_sra_39_n83), .C2(
        dp_ex_stage_alu_shifter_sra_39_n51), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n121) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U135 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n97), .B2(
        dp_ex_stage_alu_shifter_sra_39_n107), .C1(
        dp_ex_stage_alu_shifter_sra_39_n120), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n121), .ZN(dp_ex_stage_alu_shifter_N107) );
  OAI21_X1 dp_ex_stage_alu_shifter_sra_39_U134 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n18), .B2(
        dp_ex_stage_alu_shifter_sra_39_n118), .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(dp_ex_stage_alu_shifter_N135) );
  OAI22_X1 dp_ex_stage_alu_shifter_sra_39_U133 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n26), .A2(
        dp_ex_stage_alu_shifter_sra_39_n10), .B1(
        dp_ex_stage_alu_shifter_sra_39_n25), .B2(
        dp_ex_stage_alu_shifter_sra_39_n13), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n115) );
  AOI22_X1 dp_ex_stage_alu_shifter_sra_39_U132 ( .A1(dp_ex_stage_alu_n52), 
        .A2(dp_ex_stage_alu_shifter_sra_39_n73), .B1(dp_ex_stage_alu_n69), 
        .B2(dp_ex_stage_alu_shifter_sra_39_n75), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n112) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U131 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n85), .A2(
        dp_ex_stage_alu_shifter_sra_39_n95), .B1(
        dp_ex_stage_alu_shifter_sra_39_n77), .B2(
        dp_ex_stage_alu_shifter_sra_39_n110), .C1(
        dp_ex_stage_alu_shifter_sra_39_n83), .C2(
        dp_ex_stage_alu_shifter_sra_39_n52), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n109) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U130 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n92), .B2(
        dp_ex_stage_alu_shifter_sra_39_n107), .C1(
        dp_ex_stage_alu_shifter_sra_39_n108), .C2(
        dp_ex_stage_alu_shifter_sra_39_n22), .A(
        dp_ex_stage_alu_shifter_sra_39_n109), .ZN(dp_ex_stage_alu_shifter_N108) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U129 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n49), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n53), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n90), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n106) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U128 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n104), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n105), .C2(
        dp_ex_stage_alu_shifter_sra_39_n22), .A(
        dp_ex_stage_alu_shifter_sra_39_n106), .ZN(dp_ex_stage_alu_shifter_N109) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U127 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n50), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n55), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n84), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n103) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U126 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n101), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n102), .C2(
        dp_ex_stage_alu_shifter_sra_39_n22), .A(
        dp_ex_stage_alu_shifter_sra_39_n103), .ZN(dp_ex_stage_alu_shifter_N110) );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U125 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n51), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n57), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n100), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n99) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U124 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n97), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n98), .C2(
        dp_ex_stage_alu_shifter_sra_39_n22), .A(
        dp_ex_stage_alu_shifter_sra_39_n99), .ZN(dp_ex_stage_alu_shifter_N111)
         );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U123 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n52), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n95), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n96), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n94) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U122 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n92), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n93), .C2(
        dp_ex_stage_alu_shifter_sra_39_n22), .A(
        dp_ex_stage_alu_shifter_sra_39_n94), .ZN(dp_ex_stage_alu_shifter_N112)
         );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U121 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n53), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n90), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n91), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n89) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U120 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n87), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n88), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n89), .ZN(dp_ex_stage_alu_shifter_N113)
         );
  AOI222_X1 dp_ex_stage_alu_shifter_sra_39_U119 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n78), .A2(
        dp_ex_stage_alu_shifter_sra_39_n55), .B1(
        dp_ex_stage_alu_shifter_sra_39_n83), .B2(
        dp_ex_stage_alu_shifter_sra_39_n84), .C1(
        dp_ex_stage_alu_shifter_sra_39_n85), .C2(
        dp_ex_stage_alu_shifter_sra_39_n86), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n82) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U118 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n79), .B2(
        dp_ex_stage_alu_shifter_sra_39_n80), .C1(
        dp_ex_stage_alu_shifter_sra_39_n81), .C2(
        dp_ex_stage_alu_shifter_sra_39_n21), .A(
        dp_ex_stage_alu_shifter_sra_39_n82), .ZN(dp_ex_stage_alu_shifter_N114)
         );
  INV_X2 dp_ex_stage_alu_shifter_sra_39_U117 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n113), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n76) );
  INV_X2 dp_ex_stage_alu_shifter_sra_39_U116 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n114), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n74) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U115 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n45), .ZN(dp_ex_stage_alu_shifter_N136)
         );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U114 ( .A(dp_ex_stage_alu_n1), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n43) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U113 ( .A(dp_ex_stage_muxA_out[27]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n42) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U112 ( .A(dp_ex_stage_muxA_out[26]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n41) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U111 ( .A(dp_ex_stage_muxA_out[25]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n40) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U110 ( .A(dp_ex_stage_muxA_out[24]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n39) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U109 ( .A(dp_ex_stage_muxA_out[23]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n38) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U108 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n38), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n37) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U107 ( .A(dp_ex_stage_muxA_out[21]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n36) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U106 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n36), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n35) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U105 ( .A(dp_ex_stage_muxA_out[18]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n34) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U104 ( .A(dp_ex_stage_muxA_out[17]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n33) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U103 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n33), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n32) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U102 ( .A(dp_ex_stage_muxA_out[12]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n31) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U101 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n31), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n30) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U100 ( .A(dp_ex_stage_alu_n33), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n29) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U99 ( .A(dp_ex_stage_alu_n74), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n28) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U98 ( .A(dp_ex_stage_alu_n72), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n27) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U97 ( .A(dp_ex_stage_alu_n71), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n26) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U96 ( .A(dp_ex_stage_alu_n34), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n25) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U95 ( .A(dp_ex_stage_alu_n69), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n24) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U94 ( .A(dp_ex_stage_alu_n44), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n23) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U93 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n18), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n22) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U92 ( .A(dp_ex_stage_alu_n49), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n17) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U91 ( .A(dp_ex_stage_alu_n45), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n16) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U90 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n160), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n57) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U89 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n168), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n53) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U88 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n167), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n56) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U87 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n151), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n55) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U86 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n179), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n58) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U85 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n187), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n54) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U84 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n156), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n60) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U83 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n153), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n65) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U82 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n157), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n64) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U81 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n11), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n15) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U80 ( .A(dp_ex_stage_alu_n52), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n46) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U79 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n9), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n73) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U78 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n9), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n14) );
  NAND2_X1 dp_ex_stage_alu_shifter_sra_39_U77 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n16), .A2(
        dp_ex_stage_alu_shifter_sra_39_n4), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n117) );
  BUF_X1 dp_ex_stage_alu_shifter_sra_39_U76 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n117), .Z(
        dp_ex_stage_alu_shifter_sra_39_n12) );
  NAND2_X1 dp_ex_stage_alu_shifter_sra_39_U75 ( .A1(dp_ex_stage_alu_n45), .A2(
        dp_ex_stage_alu_shifter_sra_39_n3), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n116) );
  CLKBUF_X3 dp_ex_stage_alu_shifter_sra_39_U74 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n116), .Z(
        dp_ex_stage_alu_shifter_sra_39_n10) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U73 ( .A(dp_ex_stage_alu_n78), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n48) );
  BUF_X1 dp_ex_stage_alu_shifter_sra_39_U72 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n116), .Z(
        dp_ex_stage_alu_shifter_sra_39_n9) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U71 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_muxA_out[14]), 
        .C1(dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_alu_n29), 
        .A(dp_ex_stage_alu_shifter_sra_39_n54), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n168) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U70 ( .A(dp_ex_stage_alu_n70), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n47) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U69 ( .A(dp_ex_stage_muxA_out[30]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n70) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U68 ( .A(dp_ex_stage_muxA_out[20]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n63) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U67 ( .A(dp_ex_stage_muxA_out[29]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n68) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U66 ( .A(dp_ex_stage_muxA_out[19]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n62) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U65 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n38), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(
        dp_ex_stage_alu_shifter_sra_39_n32), .A(
        dp_ex_stage_alu_shifter_sra_39_n58), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n160) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U64 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n144), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n67) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U63 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n140), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n69) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U62 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n145), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n66) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U61 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n154), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n71) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U60 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n95), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n59) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U59 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n79), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n50) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U58 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n111), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n52) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U57 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n87), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n49) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U56 ( .A(dp_ex_stage_muxA_out[31]), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n45) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U55 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n119), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n72) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U54 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n96), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n61) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U53 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n123), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n51) );
  BUF_X2 dp_ex_stage_alu_shifter_sra_39_U52 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n117), .Z(
        dp_ex_stage_alu_shifter_sra_39_n13) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U51 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n80), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n77) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U50 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n107), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n78) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U49 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n18), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n21) );
  NAND2_X1 dp_ex_stage_alu_shifter_sra_39_U48 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n20), .A2(dp_ex_stage_alu_shifter_N136), 
        .ZN(dp_ex_stage_alu_shifter_sra_39_n119) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_sra_39_U47 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_sra_39_n20)
         );
  CLKBUF_X1 dp_ex_stage_alu_shifter_sra_39_U46 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_sra_39_n19)
         );
  BUF_X2 dp_ex_stage_alu_shifter_sra_39_U45 ( .A(dp_ex_stage_alu_shifter_n116), 
        .Z(dp_ex_stage_alu_shifter_sra_39_n18) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_sra_39_U44 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n135), .Z(
        dp_ex_stage_alu_shifter_sra_39_n8) );
  BUF_X1 dp_ex_stage_alu_shifter_sra_39_U43 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n134), .Z(
        dp_ex_stage_alu_shifter_sra_39_n7) );
  NAND2_X1 dp_ex_stage_alu_shifter_sra_39_U42 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n90), .A2(
        dp_ex_stage_alu_shifter_sra_39_n133), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n6) );
  NAND2_X1 dp_ex_stage_alu_shifter_sra_39_U41 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n91), .A2(
        dp_ex_stage_alu_shifter_sra_39_n131), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n5) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U40 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n86), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n84), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n64), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n146) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U39 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n137), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n96), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n65), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n108) );
  OAI221_X4 dp_ex_stage_alu_shifter_sra_39_U38 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n47), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n48), .A(
        dp_ex_stage_alu_shifter_sra_39_n112), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n110) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U37 ( .A(dp_ex_stage_alu_n46), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n4) );
  INV_X1 dp_ex_stage_alu_shifter_sra_39_U36 ( .A(dp_ex_stage_alu_n46), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n3) );
  NOR2_X2 dp_ex_stage_alu_shifter_sra_39_U35 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n16), .A2(
        dp_ex_stage_alu_shifter_sra_39_n3), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n114) );
  AND3_X1 dp_ex_stage_alu_shifter_sra_39_U34 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n5), .A2(
        dp_ex_stage_alu_shifter_sra_39_n6), .A3(
        dp_ex_stage_alu_shifter_sra_39_n188), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n158) );
  INV_X2 dp_ex_stage_alu_shifter_sra_39_U33 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n11), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n75) );
  NAND3_X1 dp_ex_stage_alu_shifter_sra_39_U32 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n1), .A2(
        dp_ex_stage_alu_shifter_sra_39_n2), .A3(
        dp_ex_stage_alu_shifter_sra_39_n189), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n135) );
  OR2_X1 dp_ex_stage_alu_shifter_sra_39_U31 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n74), .A2(
        dp_ex_stage_alu_shifter_sra_39_n42), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n2) );
  OR2_X1 dp_ex_stage_alu_shifter_sra_39_U30 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n76), .A2(
        dp_ex_stage_alu_shifter_sra_39_n41), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n1) );
  NOR2_X2 dp_ex_stage_alu_shifter_sra_39_U29 ( .A1(dp_ex_stage_alu_n49), .A2(
        dp_ex_stage_alu_n31), .ZN(dp_ex_stage_alu_shifter_sra_39_n133) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U28 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n130), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n132), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n71), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n81) );
  NAND2_X1 dp_ex_stage_alu_shifter_sra_39_U27 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n133), .A2(
        dp_ex_stage_alu_shifter_sra_39_n21), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n80) );
  AND2_X1 dp_ex_stage_alu_shifter_sra_39_U26 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n185), .A2(
        dp_ex_stage_alu_shifter_sra_39_n17), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n83) );
  NOR2_X2 dp_ex_stage_alu_shifter_sra_39_U25 ( .A1(
        dp_ex_stage_alu_shifter_sra_39_n4), .A2(dp_ex_stage_alu_n45), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n113) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U24 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n23), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n24), .A(
        dp_ex_stage_alu_shifter_sra_39_n186), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n183) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U23 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n34), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_alu_n71), .A(
        dp_ex_stage_alu_shifter_sra_39_n152), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n101) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U22 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n24), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n46), .A(
        dp_ex_stage_alu_shifter_sra_39_n150), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n148) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U21 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n46), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n47), .A(
        dp_ex_stage_alu_shifter_sra_39_n124), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n122) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U20 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n72), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_alu_n74), .A(
        dp_ex_stage_alu_shifter_sra_39_n115), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n92) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U19 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n8), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n91), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n66), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n105) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U18 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n132), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n86), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n67), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n102) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U17 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n138), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n139), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n69), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n98) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U16 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n136), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n137), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n71), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n93) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U15 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n7), .B2(
        dp_ex_stage_alu_shifter_sra_39_n131), .C1(
        dp_ex_stage_alu_shifter_sra_39_n8), .C2(
        dp_ex_stage_alu_shifter_sra_39_n133), .A(
        dp_ex_stage_alu_shifter_sra_39_n71), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n88) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U14 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n231), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_muxA_out[14]), 
        .A(dp_ex_stage_alu_shifter_sra_39_n175), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n111) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U13 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n62), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n63), .A(
        dp_ex_stage_alu_shifter_sra_39_n166), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n84) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U12 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n33), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n34), .A(
        dp_ex_stage_alu_shifter_sra_39_n173), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n95) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U11 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n40), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n41), .A(
        dp_ex_stage_alu_shifter_sra_39_n171), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n137) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U10 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n78), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_alu_n34), .A(
        dp_ex_stage_alu_shifter_sra_39_n193), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n104) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U9 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n71), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_alu_n72), .A(
        dp_ex_stage_alu_shifter_sra_39_n125), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n97) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U8 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n74), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_alu_n33), .A(
        dp_ex_stage_alu_shifter_sra_39_n184), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n87) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U7 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n33), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(
        dp_ex_stage_alu_shifter_sra_39_n30), .A(
        dp_ex_stage_alu_shifter_sra_39_n149), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n79) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U6 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(
        dp_ex_stage_alu_shifter_sra_39_n30), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_alu_n231), .A(
        dp_ex_stage_alu_shifter_sra_39_n181), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n123) );
  AOI221_X1 dp_ex_stage_alu_shifter_sra_39_U5 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n113), .B2(dp_ex_stage_alu_n29), .C1(
        dp_ex_stage_alu_shifter_sra_39_n114), .C2(dp_ex_stage_alu_n38), .A(
        dp_ex_stage_alu_shifter_sra_39_n56), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n151) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U4 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n38), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n39), .A(
        dp_ex_stage_alu_shifter_sra_39_n165), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n86) );
  OAI221_X1 dp_ex_stage_alu_shifter_sra_39_U3 ( .B1(
        dp_ex_stage_alu_shifter_sra_39_n76), .B2(
        dp_ex_stage_alu_shifter_sra_39_n43), .C1(
        dp_ex_stage_alu_shifter_sra_39_n74), .C2(
        dp_ex_stage_alu_shifter_sra_39_n68), .A(
        dp_ex_stage_alu_shifter_sra_39_n180), .ZN(
        dp_ex_stage_alu_shifter_sra_39_n138) );
  BUF_X1 dp_ex_stage_alu_shifter_sra_39_U2 ( .A(
        dp_ex_stage_alu_shifter_sra_39_n117), .Z(
        dp_ex_stage_alu_shifter_sra_39_n11) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U16 ( .A(dp_ex_stage_alu_n31), .Z(
        dp_ex_stage_alu_shifter_rol_32_n10) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U15 ( .A(dp_ex_stage_alu_n31), .Z(
        dp_ex_stage_alu_shifter_rol_32_n11) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U14 ( .A(dp_ex_stage_alu_n31), .Z(
        dp_ex_stage_alu_shifter_rol_32_n12) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U13 ( .A(dp_ex_stage_alu_n49), .Z(
        dp_ex_stage_alu_shifter_rol_32_n7) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U12 ( .A(dp_ex_stage_alu_n49), .Z(
        dp_ex_stage_alu_shifter_rol_32_n8) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U11 ( .A(dp_ex_stage_alu_n49), .Z(
        dp_ex_stage_alu_shifter_rol_32_n9) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U10 ( .A(dp_ex_stage_alu_shifter_n5), .Z(dp_ex_stage_alu_shifter_rol_32_n4) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U9 ( .A(dp_ex_stage_alu_shifter_n5), 
        .Z(dp_ex_stage_alu_shifter_rol_32_n5) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U8 ( .A(dp_ex_stage_alu_shifter_n5), 
        .Z(dp_ex_stage_alu_shifter_rol_32_n6) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U7 ( .A(dp_ex_stage_alu_shifter_n3), 
        .Z(dp_ex_stage_alu_shifter_rol_32_n3) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U6 ( .A(dp_ex_stage_alu_shifter_n3), 
        .Z(dp_ex_stage_alu_shifter_rol_32_n2) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U5 ( .A(dp_ex_stage_alu_shifter_n3), 
        .Z(dp_ex_stage_alu_shifter_rol_32_n1) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U4 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_rol_32_n15)
         );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U3 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_rol_32_n13)
         );
  CLKBUF_X1 dp_ex_stage_alu_shifter_rol_32_U2 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_rol_32_n14)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_0_0 ( .A(
        dp_ex_stage_alu_shifter_N202), .B(dp_ex_stage_alu_shifter_n1), .S(
        dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__0_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_1 ( .A(dp_ex_stage_alu_n76), .B(
        dp_ex_stage_alu_shifter_N202), .S(dp_ex_stage_alu_shifter_rol_32_n1), 
        .Z(dp_ex_stage_alu_shifter_rol_32_ML_int_1__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_2 ( .A(dp_ex_stage_alu_n44), .B(
        dp_ex_stage_alu_n76), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_3 ( .A(dp_ex_stage_alu_n69), .B(
        dp_ex_stage_alu_n44), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_4 ( .A(dp_ex_stage_alu_n52), .B(
        dp_ex_stage_alu_n69), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_5 ( .A(dp_ex_stage_alu_n70), .B(
        dp_ex_stage_alu_n52), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_6 ( .A(dp_ex_stage_alu_n78), .B(
        dp_ex_stage_alu_n70), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_7 ( .A(dp_ex_stage_alu_n34), .B(
        dp_ex_stage_alu_n78), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_8 ( .A(dp_ex_stage_alu_n71), .B(
        dp_ex_stage_alu_n34), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_9 ( .A(dp_ex_stage_alu_n72), .B(
        dp_ex_stage_alu_n71), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_10 ( .A(dp_ex_stage_alu_n74), 
        .B(dp_ex_stage_alu_n72), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_11 ( .A(dp_ex_stage_alu_n33), 
        .B(dp_ex_stage_alu_n74), .S(dp_ex_stage_alu_shifter_rol_32_n1), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_12 ( .A(dp_ex_stage_muxA_out[12]), .B(dp_ex_stage_alu_n33), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_13 ( .A(dp_ex_stage_alu_n231), 
        .B(dp_ex_stage_muxA_out[12]), .S(dp_ex_stage_alu_shifter_rol_32_n2), 
        .Z(dp_ex_stage_alu_shifter_rol_32_ML_int_1__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_14 ( .A(dp_ex_stage_muxA_out[14]), .B(dp_ex_stage_alu_n231), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_15 ( .A(dp_ex_stage_alu_n29), 
        .B(dp_ex_stage_muxA_out[14]), .S(dp_ex_stage_alu_shifter_rol_32_n2), 
        .Z(dp_ex_stage_alu_shifter_rol_32_ML_int_1__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_16 ( .A(dp_ex_stage_alu_n38), 
        .B(dp_ex_stage_alu_n29), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_17 ( .A(dp_ex_stage_muxA_out[17]), .B(dp_ex_stage_alu_n38), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_18 ( .A(dp_ex_stage_muxA_out[18]), .B(dp_ex_stage_muxA_out[17]), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_19 ( .A(dp_ex_stage_muxA_out[19]), .B(dp_ex_stage_muxA_out[18]), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_20 ( .A(dp_ex_stage_muxA_out[20]), .B(dp_ex_stage_muxA_out[19]), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_21 ( .A(dp_ex_stage_muxA_out[21]), .B(dp_ex_stage_muxA_out[20]), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_22 ( .A(dp_ex_stage_alu_n240), 
        .B(dp_ex_stage_muxA_out[21]), .S(dp_ex_stage_alu_shifter_rol_32_n2), 
        .Z(dp_ex_stage_alu_shifter_rol_32_ML_int_1__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_23 ( .A(dp_ex_stage_muxA_out[23]), .B(dp_ex_stage_alu_n240), .S(dp_ex_stage_alu_shifter_rol_32_n2), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_24 ( .A(
        dp_ex_stage_alu_shifter_n94), .B(dp_ex_stage_muxA_out[23]), .S(
        dp_ex_stage_alu_shifter_rol_32_n3), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_25 ( .A(
        dp_ex_stage_alu_shifter_n7), .B(dp_ex_stage_alu_shifter_n94), .S(
        dp_ex_stage_alu_shifter_rol_32_n3), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_26 ( .A(
        dp_ex_stage_alu_shifter_n11), .B(dp_ex_stage_alu_shifter_n7), .S(
        dp_ex_stage_alu_shifter_rol_32_n3), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_27 ( .A(
        dp_ex_stage_alu_shifter_n12), .B(dp_ex_stage_alu_shifter_n11), .S(
        dp_ex_stage_alu_shifter_rol_32_n3), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_28 ( .A(dp_ex_stage_alu_n1), .B(
        dp_ex_stage_alu_shifter_n12), .S(dp_ex_stage_alu_shifter_rol_32_n3), 
        .Z(dp_ex_stage_alu_shifter_rol_32_ML_int_1__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_29 ( .A(dp_ex_stage_muxA_out[29]), .B(dp_ex_stage_alu_n1), .S(dp_ex_stage_alu_shifter_rol_32_n3), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_30 ( .A(dp_ex_stage_muxA_out[30]), .B(dp_ex_stage_muxA_out[29]), .S(dp_ex_stage_alu_shifter_rol_32_n3), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_0_31 ( .A(
        dp_ex_stage_alu_shifter_n1), .B(dp_ex_stage_muxA_out[30]), .S(
        dp_ex_stage_alu_shifter_rol_32_n3), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_1_0 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__0_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__30_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__0_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_1_1 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__1_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__31_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_2 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__2_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__0_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_3 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__3_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__1_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_4 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__4_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__2_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_5 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__5_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__3_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_6 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__6_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__4_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_7 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__7_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__5_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_8 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__8_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__6_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_9 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__9_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__7_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_10 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__10_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__8_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_11 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__11_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__9_), .S(
        dp_ex_stage_alu_shifter_rol_32_n4), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_12 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__12_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__10_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_13 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__13_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__11_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_14 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__14_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__12_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_15 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__15_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__13_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_16 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__16_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__14_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_17 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__17_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__15_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_18 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__18_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__16_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_19 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__19_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__17_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_20 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__20_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__18_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_21 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__21_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__19_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_22 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__22_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__20_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_23 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__23_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__21_), .S(
        dp_ex_stage_alu_shifter_rol_32_n5), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_24 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__24_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__22_), .S(
        dp_ex_stage_alu_shifter_rol_32_n6), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_25 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__25_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__23_), .S(
        dp_ex_stage_alu_shifter_rol_32_n6), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_26 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__26_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__24_), .S(
        dp_ex_stage_alu_shifter_rol_32_n6), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_27 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__27_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__25_), .S(
        dp_ex_stage_alu_shifter_rol_32_n6), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_28 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__28_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__26_), .S(
        dp_ex_stage_alu_shifter_rol_32_n6), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_29 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__29_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__27_), .S(
        dp_ex_stage_alu_shifter_rol_32_n6), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_30 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__30_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__28_), .S(
        dp_ex_stage_alu_shifter_rol_32_n6), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_1_31 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__31_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_1__29_), .S(
        dp_ex_stage_alu_shifter_rol_32_n6), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_2_0 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__0_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__28_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__0_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_2_1 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__1_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__29_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_2_2 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__2_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__30_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_2_3 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__3_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__31_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_4 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__4_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__0_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_5 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__5_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__1_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_6 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__6_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__2_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_7 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__7_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__3_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_8 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__8_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__4_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_9 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__9_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__5_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_10 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__10_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__6_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_11 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__11_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__7_), .S(
        dp_ex_stage_alu_shifter_rol_32_n7), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_12 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__12_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__8_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_13 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__13_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__9_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_14 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__14_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__10_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_15 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__15_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__11_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_16 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__16_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__12_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_17 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__17_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__13_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_18 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__18_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__14_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_19 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__19_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__15_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_20 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__20_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__16_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_21 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__21_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__17_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_22 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__22_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__18_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_23 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__23_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__19_), .S(
        dp_ex_stage_alu_shifter_rol_32_n8), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_24 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__24_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__20_), .S(
        dp_ex_stage_alu_shifter_rol_32_n9), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_25 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__25_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__21_), .S(
        dp_ex_stage_alu_shifter_rol_32_n9), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_26 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__26_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__22_), .S(
        dp_ex_stage_alu_shifter_rol_32_n9), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_27 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__27_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__23_), .S(
        dp_ex_stage_alu_shifter_rol_32_n9), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_28 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__28_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__24_), .S(
        dp_ex_stage_alu_shifter_rol_32_n9), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_29 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__29_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__25_), .S(
        dp_ex_stage_alu_shifter_rol_32_n9), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_30 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__30_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__26_), .S(
        dp_ex_stage_alu_shifter_rol_32_n9), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_2_31 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__31_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_2__27_), .S(
        dp_ex_stage_alu_shifter_rol_32_n9), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_3_0 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__0_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__24_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__0_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_3_1 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__1_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__25_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_3_2 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__2_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__26_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_3_3 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__3_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__27_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_3_4 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__4_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__28_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_3_5 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__5_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__29_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_3_6 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__6_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__30_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_3_7 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__7_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__31_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_8 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__8_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__0_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_9 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__9_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__1_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_10 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__10_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__2_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_11 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__11_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__3_), .S(
        dp_ex_stage_alu_shifter_rol_32_n10), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_12 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__12_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__4_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_13 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__13_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__5_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_14 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__14_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__6_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_15 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__15_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__7_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_16 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__16_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__8_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_17 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__17_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__9_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_18 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__18_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__10_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_19 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__19_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__11_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_20 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__20_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__12_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_21 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__21_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__13_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_22 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__22_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__14_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_23 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__23_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__15_), .S(
        dp_ex_stage_alu_shifter_rol_32_n11), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_24 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__24_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__16_), .S(
        dp_ex_stage_alu_shifter_rol_32_n12), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_25 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__25_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__17_), .S(
        dp_ex_stage_alu_shifter_rol_32_n12), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_26 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__26_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__18_), .S(
        dp_ex_stage_alu_shifter_rol_32_n12), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_27 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__27_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__19_), .S(
        dp_ex_stage_alu_shifter_rol_32_n12), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_28 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__28_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__20_), .S(
        dp_ex_stage_alu_shifter_rol_32_n12), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_29 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__29_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__21_), .S(
        dp_ex_stage_alu_shifter_rol_32_n12), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_30 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__30_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__22_), .S(
        dp_ex_stage_alu_shifter_rol_32_n12), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_3_31 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__31_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_3__23_), .S(
        dp_ex_stage_alu_shifter_rol_32_n12), .Z(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_0 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__0_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__16_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N39)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_1 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__1_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__17_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N40)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_2 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__2_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__18_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N41)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_3 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__3_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__19_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N42)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_4 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__4_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__20_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N43)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_5 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__5_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__21_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N44)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_6 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__6_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__22_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N45)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_7 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__7_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__23_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N46)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_8 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__8_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__24_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N47)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_9 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__9_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__25_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N48)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_10 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__10_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__26_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N49)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_11 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__11_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__27_), .S(
        dp_ex_stage_alu_shifter_rol_32_n13), .Z(dp_ex_stage_alu_shifter_N50)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_12 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__12_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__28_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N51)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_13 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__13_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__29_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N52)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_14 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__14_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__30_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N53)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M0_4_15 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__15_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__31_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N54)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_16 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__16_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__0_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N55)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_17 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__17_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__1_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N56)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_18 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__18_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__2_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N57)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_19 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__19_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__3_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N58)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_20 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__20_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__4_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N59)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_21 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__21_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__5_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N60)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_22 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__22_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__6_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N61)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_23 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__23_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__7_), .S(
        dp_ex_stage_alu_shifter_rol_32_n14), .Z(dp_ex_stage_alu_shifter_N62)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_24 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__24_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__8_), .S(
        dp_ex_stage_alu_shifter_rol_32_n15), .Z(dp_ex_stage_alu_shifter_N63)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_25 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__25_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__9_), .S(
        dp_ex_stage_alu_shifter_rol_32_n15), .Z(dp_ex_stage_alu_shifter_N64)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_26 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__26_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__10_), .S(
        dp_ex_stage_alu_shifter_rol_32_n15), .Z(dp_ex_stage_alu_shifter_N65)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_27 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__27_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__11_), .S(
        dp_ex_stage_alu_shifter_rol_32_n15), .Z(dp_ex_stage_alu_shifter_N66)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_28 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__28_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__12_), .S(
        dp_ex_stage_alu_shifter_rol_32_n15), .Z(dp_ex_stage_alu_shifter_N67)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_29 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__29_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__13_), .S(
        dp_ex_stage_alu_shifter_rol_32_n15), .Z(dp_ex_stage_alu_shifter_N68)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_30 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__30_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__14_), .S(
        dp_ex_stage_alu_shifter_rol_32_n15), .Z(dp_ex_stage_alu_shifter_N69)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_rol_32_M1_4_31 ( .A(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__31_), .B(
        dp_ex_stage_alu_shifter_rol_32_ML_int_4__15_), .S(
        dp_ex_stage_alu_shifter_rol_32_n15), .Z(dp_ex_stage_alu_shifter_N70)
         );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U16 ( .A(dp_ex_stage_alu_n31), .Z(
        dp_ex_stage_alu_shifter_ror_30_n10) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U15 ( .A(dp_ex_stage_alu_n31), .Z(
        dp_ex_stage_alu_shifter_ror_30_n11) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U14 ( .A(dp_ex_stage_alu_n31), .Z(
        dp_ex_stage_alu_shifter_ror_30_n12) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U13 ( .A(dp_ex_stage_alu_n49), .Z(
        dp_ex_stage_alu_shifter_ror_30_n7) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U12 ( .A(dp_ex_stage_alu_n49), .Z(
        dp_ex_stage_alu_shifter_ror_30_n8) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U11 ( .A(dp_ex_stage_alu_n49), .Z(
        dp_ex_stage_alu_shifter_ror_30_n9) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U10 ( .A(dp_ex_stage_alu_shifter_n5), .Z(dp_ex_stage_alu_shifter_ror_30_n4) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U9 ( .A(dp_ex_stage_alu_shifter_n5), 
        .Z(dp_ex_stage_alu_shifter_ror_30_n5) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U8 ( .A(dp_ex_stage_alu_shifter_n5), 
        .Z(dp_ex_stage_alu_shifter_ror_30_n6) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U7 ( .A(dp_ex_stage_alu_shifter_n3), 
        .Z(dp_ex_stage_alu_shifter_ror_30_n3) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U6 ( .A(dp_ex_stage_alu_shifter_n3), 
        .Z(dp_ex_stage_alu_shifter_ror_30_n1) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U5 ( .A(dp_ex_stage_alu_shifter_n3), 
        .Z(dp_ex_stage_alu_shifter_ror_30_n2) );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U4 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_ror_30_n15)
         );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U3 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_ror_30_n13)
         );
  CLKBUF_X1 dp_ex_stage_alu_shifter_ror_30_U2 ( .A(
        dp_ex_stage_alu_shifter_n116), .Z(dp_ex_stage_alu_shifter_ror_30_n14)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_0 ( .A(
        dp_ex_stage_alu_shifter_N202), .B(dp_ex_stage_alu_n76), .S(
        dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__0_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_1_0 ( .A(dp_ex_stage_alu_n76), 
        .B(dp_ex_stage_alu_n44), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_2_0 ( .A(dp_ex_stage_alu_n44), 
        .B(dp_ex_stage_alu_n69), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_3_0 ( .A(dp_ex_stage_alu_n69), 
        .B(dp_ex_stage_alu_n52), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_4_0 ( .A(dp_ex_stage_alu_n52), 
        .B(dp_ex_stage_alu_n70), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_5_0 ( .A(dp_ex_stage_alu_n70), 
        .B(dp_ex_stage_alu_n78), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_6_0 ( .A(dp_ex_stage_alu_n78), 
        .B(dp_ex_stage_alu_n34), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_7_0 ( .A(dp_ex_stage_alu_n34), 
        .B(dp_ex_stage_alu_n71), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_8_0 ( .A(dp_ex_stage_alu_n71), 
        .B(dp_ex_stage_alu_n72), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_9_0 ( .A(dp_ex_stage_alu_n72), 
        .B(dp_ex_stage_alu_n74), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_10_0 ( .A(dp_ex_stage_alu_n74), 
        .B(dp_ex_stage_alu_n33), .S(dp_ex_stage_alu_shifter_ror_30_n1), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_11_0 ( .A(dp_ex_stage_alu_n33), 
        .B(dp_ex_stage_muxA_out[12]), .S(dp_ex_stage_alu_shifter_ror_30_n1), 
        .Z(dp_ex_stage_alu_shifter_ror_30_MR_int_1__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_12_0 ( .A(
        dp_ex_stage_muxA_out[12]), .B(dp_ex_stage_alu_n231), .S(
        dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_13_0 ( .A(dp_ex_stage_alu_n231), 
        .B(dp_ex_stage_muxA_out[14]), .S(dp_ex_stage_alu_shifter_ror_30_n2), 
        .Z(dp_ex_stage_alu_shifter_ror_30_MR_int_1__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_14_0 ( .A(
        dp_ex_stage_muxA_out[14]), .B(dp_ex_stage_alu_n29), .S(
        dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_15_0 ( .A(dp_ex_stage_alu_n29), 
        .B(dp_ex_stage_alu_n38), .S(dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_16_0 ( .A(dp_ex_stage_alu_n38), 
        .B(dp_ex_stage_muxA_out[17]), .S(dp_ex_stage_alu_shifter_ror_30_n2), 
        .Z(dp_ex_stage_alu_shifter_ror_30_MR_int_1__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_17_0 ( .A(
        dp_ex_stage_muxA_out[17]), .B(dp_ex_stage_muxA_out[18]), .S(
        dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_18_0 ( .A(
        dp_ex_stage_muxA_out[18]), .B(dp_ex_stage_muxA_out[19]), .S(
        dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_19_0 ( .A(
        dp_ex_stage_muxA_out[19]), .B(dp_ex_stage_muxA_out[20]), .S(
        dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_20_0 ( .A(
        dp_ex_stage_muxA_out[20]), .B(dp_ex_stage_muxA_out[21]), .S(
        dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_21_0 ( .A(
        dp_ex_stage_muxA_out[21]), .B(dp_ex_stage_alu_n240), .S(
        dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_22_0 ( .A(dp_ex_stage_alu_n240), 
        .B(dp_ex_stage_muxA_out[23]), .S(dp_ex_stage_alu_shifter_ror_30_n2), 
        .Z(dp_ex_stage_alu_shifter_ror_30_MR_int_1__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_23_0 ( .A(
        dp_ex_stage_muxA_out[23]), .B(dp_ex_stage_alu_shifter_n94), .S(
        dp_ex_stage_alu_shifter_ror_30_n2), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_24_0 ( .A(
        dp_ex_stage_alu_shifter_n94), .B(dp_ex_stage_alu_shifter_n7), .S(
        dp_ex_stage_alu_shifter_ror_30_n3), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_25_0 ( .A(
        dp_ex_stage_alu_shifter_n7), .B(dp_ex_stage_alu_shifter_n11), .S(
        dp_ex_stage_alu_shifter_ror_30_n3), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_26_0 ( .A(
        dp_ex_stage_alu_shifter_n11), .B(dp_ex_stage_alu_shifter_n12), .S(
        dp_ex_stage_alu_shifter_ror_30_n3), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_27_0 ( .A(
        dp_ex_stage_alu_shifter_n12), .B(dp_ex_stage_alu_n1), .S(
        dp_ex_stage_alu_shifter_ror_30_n3), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_28_0 ( .A(dp_ex_stage_alu_n1), 
        .B(dp_ex_stage_muxA_out[29]), .S(dp_ex_stage_alu_shifter_ror_30_n3), 
        .Z(dp_ex_stage_alu_shifter_ror_30_MR_int_1__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_29_0 ( .A(
        dp_ex_stage_muxA_out[29]), .B(dp_ex_stage_muxA_out[30]), .S(
        dp_ex_stage_alu_shifter_ror_30_n3), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_30_0 ( .A(
        dp_ex_stage_muxA_out[30]), .B(dp_ex_stage_alu_shifter_n1), .S(
        dp_ex_stage_alu_shifter_ror_30_n3), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_0_31_0 ( .A(
        dp_ex_stage_alu_shifter_n1), .B(dp_ex_stage_alu_shifter_N202), .S(
        dp_ex_stage_alu_shifter_ror_30_n3), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__0_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__2_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__0_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_1 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__1_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__3_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_2_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__2_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__4_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_3_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__3_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__5_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_4_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__4_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__6_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_5_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__5_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__7_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_6_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__6_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__8_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_7_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__7_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__9_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_8_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__8_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__10_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_9_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__9_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__11_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_10_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__10_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__12_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_11_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__11_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__13_), .S(
        dp_ex_stage_alu_shifter_ror_30_n4), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_12_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__12_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__14_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_13_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__13_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__15_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_14_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__14_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__16_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_15_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__15_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__17_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_16_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__16_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__18_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_17_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__17_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__19_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_18_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__18_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__20_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_19_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__19_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__21_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_20_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__20_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__22_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_21_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__21_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__23_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_22_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__22_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__24_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_23_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__23_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__25_), .S(
        dp_ex_stage_alu_shifter_ror_30_n5), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_24_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__24_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__26_), .S(
        dp_ex_stage_alu_shifter_ror_30_n6), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_25_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__25_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__27_), .S(
        dp_ex_stage_alu_shifter_ror_30_n6), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_26_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__26_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__28_), .S(
        dp_ex_stage_alu_shifter_ror_30_n6), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_27_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__27_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__29_), .S(
        dp_ex_stage_alu_shifter_ror_30_n6), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_28_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__28_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__30_), .S(
        dp_ex_stage_alu_shifter_ror_30_n6), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_29_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__29_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__31_), .S(
        dp_ex_stage_alu_shifter_ror_30_n6), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_30_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__30_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__0_), .S(
        dp_ex_stage_alu_shifter_ror_30_n6), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_1_31_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__31_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_1__1_), .S(
        dp_ex_stage_alu_shifter_ror_30_n6), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__0_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__4_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__0_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_1 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__1_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__5_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_2 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__2_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__6_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_3 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__3_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__7_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_4_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__4_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__8_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_5_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__5_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__9_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_6_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__6_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__10_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_7_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__7_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__11_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_8_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__8_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__12_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_9_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__9_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__13_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_10_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__10_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__14_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_11_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__11_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__15_), .S(
        dp_ex_stage_alu_shifter_ror_30_n7), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_12_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__12_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__16_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_13_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__13_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__17_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_14_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__14_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__18_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_15_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__15_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__19_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_16_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__16_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__20_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_17_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__17_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__21_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_18_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__18_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__22_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_19_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__19_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__23_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_20_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__20_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__24_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_21_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__21_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__25_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_22_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__22_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__26_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_23_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__23_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__27_), .S(
        dp_ex_stage_alu_shifter_ror_30_n8), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_24_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__24_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__28_), .S(
        dp_ex_stage_alu_shifter_ror_30_n9), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_25_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__25_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__29_), .S(
        dp_ex_stage_alu_shifter_ror_30_n9), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_26_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__26_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__30_), .S(
        dp_ex_stage_alu_shifter_ror_30_n9), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_27_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__27_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__31_), .S(
        dp_ex_stage_alu_shifter_ror_30_n9), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_28_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__28_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__0_), .S(
        dp_ex_stage_alu_shifter_ror_30_n9), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_29_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__29_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__1_), .S(
        dp_ex_stage_alu_shifter_ror_30_n9), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_30_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__30_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__2_), .S(
        dp_ex_stage_alu_shifter_ror_30_n9), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_2_31_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__31_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_2__3_), .S(
        dp_ex_stage_alu_shifter_ror_30_n9), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__0_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__8_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__0_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_1 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__1_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__9_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__1_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_2 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__2_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__10_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__2_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_3 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__3_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__11_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__3_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_4 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__4_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__12_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__4_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_5 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__5_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__13_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__5_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_6 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__6_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__14_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__6_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_7 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__7_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__15_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__7_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_8_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__8_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__16_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__8_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_9_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__9_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__17_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__9_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_10_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__10_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__18_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__10_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_11_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__11_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__19_), .S(
        dp_ex_stage_alu_shifter_ror_30_n10), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__11_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_12_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__12_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__20_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__12_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_13_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__13_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__21_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__13_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_14_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__14_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__22_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__14_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_15_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__15_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__23_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__15_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_16_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__16_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__24_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__16_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_17_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__17_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__25_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__17_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_18_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__18_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__26_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__18_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_19_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__19_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__27_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__19_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_20_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__20_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__28_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__20_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_21_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__21_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__29_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__21_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_22_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__22_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__30_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__22_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_23_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__23_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__31_), .S(
        dp_ex_stage_alu_shifter_ror_30_n11), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__23_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_24_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__24_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__0_), .S(
        dp_ex_stage_alu_shifter_ror_30_n12), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__24_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_25_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__25_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__1_), .S(
        dp_ex_stage_alu_shifter_ror_30_n12), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__25_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_26_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__26_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__2_), .S(
        dp_ex_stage_alu_shifter_ror_30_n12), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__26_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_27_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__27_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__3_), .S(
        dp_ex_stage_alu_shifter_ror_30_n12), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__27_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_28_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__28_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__4_), .S(
        dp_ex_stage_alu_shifter_ror_30_n12), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__28_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_29_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__29_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__5_), .S(
        dp_ex_stage_alu_shifter_ror_30_n12), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__29_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_30_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__30_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__6_), .S(
        dp_ex_stage_alu_shifter_ror_30_n12), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__30_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_3_31_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__31_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_3__7_), .S(
        dp_ex_stage_alu_shifter_ror_30_n12), .Z(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__31_) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_0 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__0_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__16_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N7) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_1 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__1_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__17_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N8) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_2 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__2_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__18_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N9) );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_3 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__3_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__19_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N10)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_4 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__4_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__20_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N11)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_5 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__5_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__21_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N12)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_6 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__6_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__22_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N13)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_7 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__7_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__23_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N14)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_8 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__8_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__24_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N15)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_9 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__9_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__25_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N16)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_10 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__10_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__26_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N17)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_11 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__11_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__27_), .S(
        dp_ex_stage_alu_shifter_ror_30_n13), .Z(dp_ex_stage_alu_shifter_N18)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_12 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__12_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__28_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N19)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_13 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__13_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__29_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N20)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_14 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__14_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__30_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N21)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_15 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__15_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__31_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N22)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_16 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__16_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__0_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N23)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_17 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__17_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__1_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N24)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_18 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__18_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__2_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N25)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_19 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__19_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__3_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N26)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_20 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__20_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__4_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N27)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_21 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__21_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__5_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N28)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_22 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__22_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__6_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N29)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_23 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__23_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__7_), .S(
        dp_ex_stage_alu_shifter_ror_30_n14), .Z(dp_ex_stage_alu_shifter_N30)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_24 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__24_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__8_), .S(
        dp_ex_stage_alu_shifter_ror_30_n15), .Z(dp_ex_stage_alu_shifter_N31)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_25 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__25_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__9_), .S(
        dp_ex_stage_alu_shifter_ror_30_n15), .Z(dp_ex_stage_alu_shifter_N32)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_26 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__26_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__10_), .S(
        dp_ex_stage_alu_shifter_ror_30_n15), .Z(dp_ex_stage_alu_shifter_N33)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_27 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__27_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__11_), .S(
        dp_ex_stage_alu_shifter_ror_30_n15), .Z(dp_ex_stage_alu_shifter_N34)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_28 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__28_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__12_), .S(
        dp_ex_stage_alu_shifter_ror_30_n15), .Z(dp_ex_stage_alu_shifter_N35)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_29 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__29_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__13_), .S(
        dp_ex_stage_alu_shifter_ror_30_n15), .Z(dp_ex_stage_alu_shifter_N36)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_30 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__30_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__14_), .S(
        dp_ex_stage_alu_shifter_ror_30_n15), .Z(dp_ex_stage_alu_shifter_N37)
         );
  MUX2_X1 dp_ex_stage_alu_shifter_ror_30_M1_4_31 ( .A(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__31_), .B(
        dp_ex_stage_alu_shifter_ror_30_MR_int_4__15_), .S(
        dp_ex_stage_alu_shifter_ror_30_n15), .Z(dp_ex_stage_alu_shifter_N38)
         );
  INV_X1 dp_ex_stage_alu_r61_U225 ( .A(dp_ex_stage_alu_r61_n91), .ZN(
        dp_ex_stage_alu_r61_n218) );
  INV_X1 dp_ex_stage_alu_r61_U224 ( .A(dp_ex_stage_alu_r61_n51), .ZN(
        dp_ex_stage_alu_r61_n219) );
  INV_X1 dp_ex_stage_alu_r61_U223 ( .A(dp_ex_stage_alu_r61_n45), .ZN(
        dp_ex_stage_alu_r61_n216) );
  NAND3_X1 dp_ex_stage_alu_r61_U222 ( .A1(dp_ex_stage_alu_r61_n155), .A2(
        dp_ex_stage_alu_r61_n147), .A3(dp_ex_stage_alu_r61_n216), .ZN(
        dp_ex_stage_alu_r61_n212) );
  NAND3_X1 dp_ex_stage_alu_r61_U221 ( .A1(dp_ex_stage_alu_r61_n211), .A2(
        dp_ex_stage_alu_r61_n212), .A3(dp_ex_stage_alu_r61_n213), .ZN(
        dp_ex_stage_alu_r61_n122) );
  INV_X1 dp_ex_stage_alu_r61_U220 ( .A(dp_ex_stage_alu_r61_n75), .ZN(
        dp_ex_stage_alu_r61_n207) );
  INV_X1 dp_ex_stage_alu_r61_U219 ( .A(dp_ex_stage_alu_r61_n88), .ZN(
        dp_ex_stage_alu_r61_n208) );
  INV_X1 dp_ex_stage_alu_r61_U218 ( .A(dp_ex_stage_alu_r61_n82), .ZN(
        dp_ex_stage_alu_r61_n204) );
  NAND3_X1 dp_ex_stage_alu_r61_U217 ( .A1(dp_ex_stage_alu_r61_n186), .A2(
        dp_ex_stage_alu_r61_n193), .A3(dp_ex_stage_alu_r61_n204), .ZN(
        dp_ex_stage_alu_r61_n202) );
  NAND3_X1 dp_ex_stage_alu_r61_U216 ( .A1(dp_ex_stage_alu_r61_n201), .A2(
        dp_ex_stage_alu_r61_n202), .A3(dp_ex_stage_alu_r61_n203), .ZN(
        dp_ex_stage_alu_r61_n166) );
  INV_X1 dp_ex_stage_alu_r61_U215 ( .A(dp_ex_stage_alu_r61_n193), .ZN(
        dp_ex_stage_alu_r61_n192) );
  INV_X1 dp_ex_stage_alu_r61_U214 ( .A(dp_ex_stage_alu_r61_n161), .ZN(
        dp_ex_stage_alu_r61_n179) );
  INV_X1 dp_ex_stage_alu_r61_U213 ( .A(dp_ex_stage_alu_r61_n87), .ZN(
        dp_ex_stage_alu_r61_n164) );
  INV_X1 dp_ex_stage_alu_r61_U212 ( .A(dp_ex_stage_alu_r61_n92), .ZN(
        dp_ex_stage_alu_r61_n165) );
  INV_X1 dp_ex_stage_alu_r61_U211 ( .A(dp_ex_stage_alu_r61_n86), .ZN(
        dp_ex_stage_alu_r61_n163) );
  NAND3_X1 dp_ex_stage_alu_r61_U210 ( .A1(dp_ex_stage_alu_r61_n2), .A2(
        dp_ex_stage_alu_r61_n162), .A3(dp_ex_stage_alu_r61_n163), .ZN(
        dp_ex_stage_alu_r61_n157) );
  INV_X1 dp_ex_stage_alu_r61_U209 ( .A(dp_ex_stage_alu_r61_n93), .ZN(
        dp_ex_stage_alu_r61_n160) );
  INV_X1 dp_ex_stage_alu_r61_U208 ( .A(dp_ex_stage_alu_r61_n155), .ZN(
        dp_ex_stage_alu_r61_n154) );
  INV_X1 dp_ex_stage_alu_r61_U207 ( .A(dp_ex_stage_alu_r61_n147), .ZN(
        dp_ex_stage_alu_r61_n146) );
  NAND3_X1 dp_ex_stage_alu_r61_U206 ( .A1(dp_ex_stage_alu_r61_n142), .A2(
        dp_ex_stage_alu_r61_n143), .A3(dp_ex_stage_alu_r61_n144), .ZN(
        dp_ex_stage_alu_r61_n141) );
  INV_X1 dp_ex_stage_alu_r61_U205 ( .A(dp_ex_stage_alu_r61_n117), .ZN(
        dp_ex_stage_alu_r61_n137) );
  INV_X1 dp_ex_stage_alu_r61_U204 ( .A(dp_ex_stage_alu_r61_n118), .ZN(
        dp_ex_stage_alu_r61_n129) );
  INV_X1 dp_ex_stage_alu_r61_U203 ( .A(dp_ex_stage_alu_r61_n50), .ZN(
        dp_ex_stage_alu_r61_n121) );
  NAND2_X1 dp_ex_stage_alu_r61_U202 ( .A1(dp_ex_stage_alu_r61_n117), .A2(
        dp_ex_stage_alu_r61_n121), .ZN(dp_ex_stage_alu_r61_n119) );
  NAND2_X1 dp_ex_stage_alu_r61_U201 ( .A1(dp_ex_stage_alu_r61_n119), .A2(
        dp_ex_stage_alu_r61_n120), .ZN(dp_ex_stage_alu_r61_n114) );
  NAND2_X1 dp_ex_stage_alu_r61_U200 ( .A1(dp_ex_stage_alu_r61_n97), .A2(
        dp_ex_stage_alu_r61_n98), .ZN(dp_ex_stage_alu_r61_n96) );
  NAND4_X1 dp_ex_stage_alu_r61_U199 ( .A1(dp_ex_stage_alu_r61_n67), .A2(
        dp_ex_stage_alu_r61_n68), .A3(dp_ex_stage_alu_r61_n69), .A4(
        dp_ex_stage_alu_r61_n70), .ZN(dp_ex_stage_alu_r61_n34) );
  XNOR2_X1 dp_ex_stage_alu_r61_U198 ( .A(dp_ex_stage_muxB_out[31]), .B(
        dp_ex_stage_alu_r61_n31), .ZN(dp_ex_stage_alu_r61_n60) );
  NAND2_X1 dp_ex_stage_alu_r61_U197 ( .A1(dp_ex_stage_alu_r61_n60), .A2(
        dp_ex_stage_alu_r61_n61), .ZN(dp_ex_stage_alu_r61_n59) );
  INV_X1 dp_ex_stage_alu_r61_U196 ( .A(dp_ex_stage_alu_N18), .ZN(
        dp_ex_stage_alu_N19) );
  INV_X1 dp_ex_stage_alu_r61_U195 ( .A(dp_ex_stage_muxA_out[31]), .ZN(
        dp_ex_stage_alu_r61_n32) );
  INV_X1 dp_ex_stage_alu_r61_U194 ( .A(dp_ex_stage_alu_r61_n32), .ZN(
        dp_ex_stage_alu_r61_n31) );
  INV_X1 dp_ex_stage_alu_r61_U193 ( .A(dp_ex_stage_alu_n247), .ZN(
        dp_ex_stage_alu_r61_n30) );
  INV_X1 dp_ex_stage_alu_r61_U192 ( .A(dp_ex_stage_muxA_out[27]), .ZN(
        dp_ex_stage_alu_r61_n29) );
  INV_X1 dp_ex_stage_alu_r61_U191 ( .A(dp_ex_stage_muxA_out[26]), .ZN(
        dp_ex_stage_alu_r61_n28) );
  INV_X1 dp_ex_stage_alu_r61_U190 ( .A(dp_ex_stage_muxA_out[25]), .ZN(
        dp_ex_stage_alu_r61_n27) );
  INV_X1 dp_ex_stage_alu_r61_U189 ( .A(dp_ex_stage_muxA_out[24]), .ZN(
        dp_ex_stage_alu_r61_n26) );
  INV_X1 dp_ex_stage_alu_r61_U188 ( .A(dp_ex_stage_muxA_out[23]), .ZN(
        dp_ex_stage_alu_r61_n25) );
  INV_X1 dp_ex_stage_alu_r61_U187 ( .A(dp_ex_stage_muxA_out[22]), .ZN(
        dp_ex_stage_alu_r61_n24) );
  INV_X1 dp_ex_stage_alu_r61_U186 ( .A(dp_ex_stage_muxA_out[21]), .ZN(
        dp_ex_stage_alu_r61_n23) );
  INV_X1 dp_ex_stage_alu_r61_U185 ( .A(dp_ex_stage_muxA_out[18]), .ZN(
        dp_ex_stage_alu_r61_n22) );
  INV_X1 dp_ex_stage_alu_r61_U184 ( .A(dp_ex_stage_muxA_out[17]), .ZN(
        dp_ex_stage_alu_r61_n21) );
  INV_X1 dp_ex_stage_alu_r61_U183 ( .A(dp_ex_stage_muxA_out[16]), .ZN(
        dp_ex_stage_alu_r61_n20) );
  INV_X1 dp_ex_stage_alu_r61_U182 ( .A(dp_ex_stage_muxA_out[15]), .ZN(
        dp_ex_stage_alu_r61_n19) );
  INV_X1 dp_ex_stage_alu_r61_U181 ( .A(dp_ex_stage_muxA_out[14]), .ZN(
        dp_ex_stage_alu_r61_n18) );
  INV_X1 dp_ex_stage_alu_r61_U180 ( .A(dp_ex_stage_muxA_out[13]), .ZN(
        dp_ex_stage_alu_r61_n17) );
  INV_X1 dp_ex_stage_alu_r61_U179 ( .A(dp_ex_stage_muxA_out[12]), .ZN(
        dp_ex_stage_alu_r61_n16) );
  INV_X1 dp_ex_stage_alu_r61_U178 ( .A(dp_ex_stage_muxA_out[11]), .ZN(
        dp_ex_stage_alu_r61_n15) );
  INV_X1 dp_ex_stage_alu_r61_U177 ( .A(dp_ex_stage_alu_n30), .ZN(
        dp_ex_stage_alu_r61_n14) );
  INV_X1 dp_ex_stage_alu_r61_U176 ( .A(dp_ex_stage_muxA_out[9]), .ZN(
        dp_ex_stage_alu_r61_n13) );
  INV_X1 dp_ex_stage_alu_r61_U175 ( .A(dp_ex_stage_muxA_out[8]), .ZN(
        dp_ex_stage_alu_r61_n12) );
  INV_X1 dp_ex_stage_alu_r61_U174 ( .A(dp_ex_stage_muxA_out[7]), .ZN(
        dp_ex_stage_alu_r61_n11) );
  INV_X1 dp_ex_stage_alu_r61_U173 ( .A(dp_ex_stage_muxA_out[3]), .ZN(
        dp_ex_stage_alu_r61_n10) );
  INV_X1 dp_ex_stage_alu_r61_U172 ( .A(dp_ex_stage_muxA_out[2]), .ZN(
        dp_ex_stage_alu_r61_n9) );
  INV_X1 dp_ex_stage_alu_r61_U171 ( .A(dp_ex_stage_alu_n22), .ZN(
        dp_ex_stage_alu_r61_n8) );
  INV_X1 dp_ex_stage_alu_r61_U170 ( .A(dp_ex_stage_alu_n50), .ZN(
        dp_ex_stage_alu_r61_n7) );
  NAND2_X1 dp_ex_stage_alu_r61_U169 ( .A1(dp_ex_stage_alu_n77), .A2(
        dp_ex_stage_alu_r61_n10), .ZN(dp_ex_stage_alu_r61_n76) );
  NOR2_X1 dp_ex_stage_alu_r61_U168 ( .A1(dp_ex_stage_alu_n77), .A2(
        dp_ex_stage_alu_r61_n10), .ZN(dp_ex_stage_alu_r61_n187) );
  NOR2_X1 dp_ex_stage_alu_r61_U167 ( .A1(dp_ex_stage_alu_n46), .A2(
        dp_ex_stage_alu_r61_n66), .ZN(dp_ex_stage_alu_r61_n199) );
  NAND2_X1 dp_ex_stage_alu_r61_U166 ( .A1(dp_ex_stage_alu_n46), .A2(
        dp_ex_stage_alu_r61_n66), .ZN(dp_ex_stage_alu_r61_n200) );
  NAND2_X1 dp_ex_stage_alu_r61_U165 ( .A1(dp_ex_stage_alu_n46), .A2(
        dp_ex_stage_alu_r61_n66), .ZN(dp_ex_stage_alu_r61_n63) );
  OAI21_X1 dp_ex_stage_alu_r61_U164 ( .B1(dp_ex_stage_alu_r61_n167), .B2(
        dp_ex_stage_alu_r61_n166), .A(dp_ex_stage_alu_r61_n168), .ZN(
        dp_ex_stage_alu_r61_n139) );
  AOI21_X1 dp_ex_stage_alu_r61_U163 ( .B1(dp_ex_stage_alu_r61_n139), .B2(
        dp_ex_stage_alu_r61_n140), .A(dp_ex_stage_alu_r61_n141), .ZN(
        dp_ex_stage_alu_r61_n123) );
  OAI21_X1 dp_ex_stage_alu_r61_U162 ( .B1(dp_ex_stage_alu_r61_n123), .B2(
        dp_ex_stage_alu_r61_n122), .A(dp_ex_stage_alu_r61_n124), .ZN(
        dp_ex_stage_alu_r61_n107) );
  AOI21_X1 dp_ex_stage_alu_r61_U161 ( .B1(dp_ex_stage_alu_r61_n107), .B2(
        dp_ex_stage_alu_r61_n108), .A(dp_ex_stage_alu_r61_n109), .ZN(
        dp_ex_stage_alu_r61_n102) );
  NAND2_X1 dp_ex_stage_alu_r61_U160 ( .A1(dp_ex_stage_alu_n30), .A2(
        dp_ex_stage_alu_r61_n176), .ZN(dp_ex_stage_alu_r61_n173) );
  INV_X1 dp_ex_stage_alu_r61_U159 ( .A(dp_ex_stage_alu_n23), .ZN(
        dp_ex_stage_alu_r61_n197) );
  NAND2_X1 dp_ex_stage_alu_r61_U158 ( .A1(dp_ex_stage_alu_n23), .A2(
        dp_ex_stage_alu_r61_n8), .ZN(dp_ex_stage_alu_r61_n194) );
  NAND2_X1 dp_ex_stage_alu_r61_U157 ( .A1(dp_ex_stage_alu_n50), .A2(
        dp_ex_stage_alu_r61_n9), .ZN(dp_ex_stage_alu_r61_n73) );
  INV_X1 dp_ex_stage_alu_r61_U156 ( .A(dp_ex_stage_muxA_out[6]), .ZN(
        dp_ex_stage_alu_r61_n209) );
  NAND2_X1 dp_ex_stage_alu_r61_U155 ( .A1(dp_ex_stage_muxA_out[6]), .A2(
        dp_ex_stage_alu_r61_n206), .ZN(dp_ex_stage_alu_r61_n193) );
  NAND2_X1 dp_ex_stage_alu_r61_U154 ( .A1(dp_ex_stage_muxB_out[30]), .A2(
        dp_ex_stage_alu_r61_n62), .ZN(dp_ex_stage_alu_r61_n100) );
  AND3_X1 dp_ex_stage_alu_r61_U153 ( .A1(dp_ex_stage_alu_r61_n99), .A2(
        dp_ex_stage_alu_r61_n100), .A3(dp_ex_stage_alu_r61_n54), .ZN(
        dp_ex_stage_alu_r61_n98) );
  INV_X1 dp_ex_stage_alu_r61_U152 ( .A(dp_ex_stage_muxB_out[5]), .ZN(
        dp_ex_stage_alu_r61_n196) );
  NAND2_X1 dp_ex_stage_alu_r61_U151 ( .A1(dp_ex_stage_muxA_out[5]), .A2(
        dp_ex_stage_alu_r61_n196), .ZN(dp_ex_stage_alu_r61_n195) );
  NAND2_X1 dp_ex_stage_alu_r61_U150 ( .A1(dp_ex_stage_alu_r61_n194), .A2(
        dp_ex_stage_alu_r61_n195), .ZN(dp_ex_stage_alu_r61_n191) );
  INV_X1 dp_ex_stage_alu_r61_U149 ( .A(dp_ex_stage_muxB_out[27]), .ZN(
        dp_ex_stage_alu_r61_n113) );
  NAND2_X1 dp_ex_stage_alu_r61_U148 ( .A1(dp_ex_stage_muxA_out[26]), .A2(
        dp_ex_stage_alu_r61_n112), .ZN(dp_ex_stage_alu_r61_n111) );
  NAND2_X1 dp_ex_stage_alu_r61_U147 ( .A1(dp_ex_stage_muxA_out[27]), .A2(
        dp_ex_stage_alu_r61_n113), .ZN(dp_ex_stage_alu_r61_n110) );
  NAND2_X1 dp_ex_stage_alu_r61_U146 ( .A1(dp_ex_stage_alu_r61_n110), .A2(
        dp_ex_stage_alu_r61_n111), .ZN(dp_ex_stage_alu_r61_n109) );
  INV_X1 dp_ex_stage_alu_r61_U145 ( .A(dp_ex_stage_muxB_out[10]), .ZN(
        dp_ex_stage_alu_r61_n176) );
  NOR2_X1 dp_ex_stage_alu_r61_U144 ( .A1(dp_ex_stage_muxB_out[30]), .A2(
        dp_ex_stage_alu_r61_n62), .ZN(dp_ex_stage_alu_r61_n222) );
  INV_X1 dp_ex_stage_alu_r61_U143 ( .A(dp_ex_stage_muxB_out[22]), .ZN(
        dp_ex_stage_alu_r61_n134) );
  INV_X1 dp_ex_stage_alu_r61_U142 ( .A(dp_ex_stage_muxB_out[26]), .ZN(
        dp_ex_stage_alu_r61_n112) );
  INV_X1 dp_ex_stage_alu_r61_U141 ( .A(dp_ex_stage_muxA_out[1]), .ZN(
        dp_ex_stage_alu_r61_n66) );
  NOR2_X1 dp_ex_stage_alu_r61_U140 ( .A1(dp_ex_stage_muxB_out[31]), .A2(
        dp_ex_stage_alu_r61_n32), .ZN(dp_ex_stage_alu_r61_n221) );
  NOR2_X1 dp_ex_stage_alu_r61_U139 ( .A1(dp_ex_stage_alu_r61_n221), .A2(
        dp_ex_stage_alu_r61_n1), .ZN(dp_ex_stage_alu_r61_n95) );
  NAND2_X1 dp_ex_stage_alu_r61_U138 ( .A1(dp_ex_stage_muxB_out[6]), .A2(
        dp_ex_stage_alu_r61_n209), .ZN(dp_ex_stage_alu_r61_n75) );
  NAND2_X1 dp_ex_stage_alu_r61_U137 ( .A1(dp_ex_stage_muxB_out[7]), .A2(
        dp_ex_stage_alu_r61_n11), .ZN(dp_ex_stage_alu_r61_n80) );
  NAND2_X1 dp_ex_stage_alu_r61_U136 ( .A1(dp_ex_stage_muxB_out[8]), .A2(
        dp_ex_stage_alu_r61_n12), .ZN(dp_ex_stage_alu_r61_n81) );
  INV_X1 dp_ex_stage_alu_r61_U135 ( .A(dp_ex_stage_muxB_out[17]), .ZN(
        dp_ex_stage_alu_r61_n150) );
  INV_X1 dp_ex_stage_alu_r61_U134 ( .A(dp_ex_stage_alu_n21), .ZN(
        dp_ex_stage_alu_r61_n65) );
  NOR2_X1 dp_ex_stage_alu_r61_U133 ( .A1(dp_ex_stage_alu_r61_n145), .A2(
        dp_ex_stage_alu_r61_n146), .ZN(dp_ex_stage_alu_r61_n144) );
  NAND4_X1 dp_ex_stage_alu_r61_U132 ( .A1(dp_ex_stage_muxA_out[14]), .A2(
        dp_ex_stage_alu_r61_n92), .A3(dp_ex_stage_alu_r61_n93), .A4(
        dp_ex_stage_alu_r61_n152), .ZN(dp_ex_stage_alu_r61_n143) );
  AOI21_X1 dp_ex_stage_alu_r61_U131 ( .B1(dp_ex_stage_alu_r61_n153), .B2(
        dp_ex_stage_alu_r61_n93), .A(dp_ex_stage_alu_r61_n154), .ZN(
        dp_ex_stage_alu_r61_n142) );
  AND2_X1 dp_ex_stage_alu_r61_U130 ( .A1(dp_ex_stage_alu_r61_n173), .A2(
        dp_ex_stage_alu_r61_n174), .ZN(dp_ex_stage_alu_r61_n6) );
  AND2_X1 dp_ex_stage_alu_r61_U129 ( .A1(dp_ex_stage_alu_r61_n6), .A2(
        dp_ex_stage_alu_r61_n162), .ZN(dp_ex_stage_alu_r61_n171) );
  INV_X1 dp_ex_stage_alu_r61_U128 ( .A(dp_ex_stage_muxB_out[14]), .ZN(
        dp_ex_stage_alu_r61_n152) );
  INV_X1 dp_ex_stage_alu_r61_U127 ( .A(dp_ex_stage_muxB_out[16]), .ZN(
        dp_ex_stage_alu_r61_n151) );
  NAND2_X1 dp_ex_stage_alu_r61_U126 ( .A1(dp_ex_stage_muxA_out[17]), .A2(
        dp_ex_stage_alu_r61_n150), .ZN(dp_ex_stage_alu_r61_n149) );
  NAND2_X1 dp_ex_stage_alu_r61_U125 ( .A1(dp_ex_stage_muxA_out[16]), .A2(
        dp_ex_stage_alu_r61_n151), .ZN(dp_ex_stage_alu_r61_n148) );
  NAND2_X1 dp_ex_stage_alu_r61_U124 ( .A1(dp_ex_stage_alu_r61_n148), .A2(
        dp_ex_stage_alu_r61_n149), .ZN(dp_ex_stage_alu_r61_n145) );
  INV_X1 dp_ex_stage_alu_r61_U123 ( .A(dp_ex_stage_muxB_out[6]), .ZN(
        dp_ex_stage_alu_r61_n206) );
  NAND2_X1 dp_ex_stage_alu_r61_U122 ( .A1(dp_ex_stage_muxB_out[26]), .A2(
        dp_ex_stage_alu_r61_n28), .ZN(dp_ex_stage_alu_r61_n48) );
  NAND2_X1 dp_ex_stage_alu_r61_U121 ( .A1(dp_ex_stage_muxB_out[25]), .A2(
        dp_ex_stage_alu_r61_n27), .ZN(dp_ex_stage_alu_r61_n57) );
  INV_X1 dp_ex_stage_alu_r61_U120 ( .A(dp_ex_stage_muxB_out[7]), .ZN(
        dp_ex_stage_alu_r61_n210) );
  NAND2_X1 dp_ex_stage_alu_r61_U119 ( .A1(dp_ex_stage_muxA_out[7]), .A2(
        dp_ex_stage_alu_r61_n210), .ZN(dp_ex_stage_alu_r61_n186) );
  NAND2_X1 dp_ex_stage_alu_r61_U118 ( .A1(dp_ex_stage_muxB_out[18]), .A2(
        dp_ex_stage_alu_r61_n22), .ZN(dp_ex_stage_alu_r61_n91) );
  NAND2_X1 dp_ex_stage_alu_r61_U117 ( .A1(dp_ex_stage_muxB_out[24]), .A2(
        dp_ex_stage_alu_r61_n26), .ZN(dp_ex_stage_alu_r61_n50) );
  NAND2_X1 dp_ex_stage_alu_r61_U116 ( .A1(dp_ex_stage_muxB_out[29]), .A2(
        dp_ex_stage_alu_r61_n101), .ZN(dp_ex_stage_alu_r61_n54) );
  NAND2_X1 dp_ex_stage_alu_r61_U115 ( .A1(dp_ex_stage_muxB_out[30]), .A2(
        dp_ex_stage_alu_r61_n62), .ZN(dp_ex_stage_alu_r61_n61) );
  INV_X1 dp_ex_stage_alu_r61_U114 ( .A(dp_ex_stage_muxA_out[5]), .ZN(
        dp_ex_stage_alu_r61_n205) );
  NAND2_X1 dp_ex_stage_alu_r61_U113 ( .A1(dp_ex_stage_muxB_out[5]), .A2(
        dp_ex_stage_alu_r61_n205), .ZN(dp_ex_stage_alu_r61_n82) );
  NAND2_X1 dp_ex_stage_alu_r61_U112 ( .A1(dp_ex_stage_muxB_out[11]), .A2(
        dp_ex_stage_alu_r61_n15), .ZN(dp_ex_stage_alu_r61_n86) );
  INV_X1 dp_ex_stage_alu_r61_U111 ( .A(dp_ex_stage_muxA_out[20]), .ZN(
        dp_ex_stage_alu_r61_n215) );
  NAND2_X1 dp_ex_stage_alu_r61_U110 ( .A1(dp_ex_stage_muxB_out[20]), .A2(
        dp_ex_stage_alu_r61_n215), .ZN(dp_ex_stage_alu_r61_n44) );
  NAND2_X1 dp_ex_stage_alu_r61_U109 ( .A1(dp_ex_stage_muxB_out[27]), .A2(
        dp_ex_stage_alu_r61_n29), .ZN(dp_ex_stage_alu_r61_n55) );
  NAND2_X1 dp_ex_stage_alu_r61_U108 ( .A1(dp_ex_stage_muxB_out[23]), .A2(
        dp_ex_stage_alu_r61_n25), .ZN(dp_ex_stage_alu_r61_n49) );
  INV_X1 dp_ex_stage_alu_r61_U107 ( .A(dp_ex_stage_muxB_out[8]), .ZN(
        dp_ex_stage_alu_r61_n177) );
  NAND4_X1 dp_ex_stage_alu_r61_U106 ( .A1(dp_ex_stage_muxA_out[8]), .A2(
        dp_ex_stage_alu_r61_n88), .A3(dp_ex_stage_alu_r61_n79), .A4(
        dp_ex_stage_alu_r61_n177), .ZN(dp_ex_stage_alu_r61_n170) );
  NAND2_X1 dp_ex_stage_alu_r61_U105 ( .A1(dp_ex_stage_muxB_out[14]), .A2(
        dp_ex_stage_alu_r61_n18), .ZN(dp_ex_stage_alu_r61_n85) );
  NOR2_X1 dp_ex_stage_alu_r61_U104 ( .A1(dp_ex_stage_muxB_out[15]), .A2(
        dp_ex_stage_alu_r61_n19), .ZN(dp_ex_stage_alu_r61_n153) );
  NAND2_X1 dp_ex_stage_alu_r61_U103 ( .A1(dp_ex_stage_muxB_out[13]), .A2(
        dp_ex_stage_alu_r61_n17), .ZN(dp_ex_stage_alu_r61_n94) );
  NOR2_X1 dp_ex_stage_alu_r61_U102 ( .A1(dp_ex_stage_muxB_out[28]), .A2(
        dp_ex_stage_alu_r61_n30), .ZN(dp_ex_stage_alu_r61_n105) );
  NAND2_X1 dp_ex_stage_alu_r61_U101 ( .A1(dp_ex_stage_muxB_out[28]), .A2(
        dp_ex_stage_alu_r61_n30), .ZN(dp_ex_stage_alu_r61_n56) );
  NOR2_X1 dp_ex_stage_alu_r61_U100 ( .A1(dp_ex_stage_muxB_out[21]), .A2(
        dp_ex_stage_alu_r61_n23), .ZN(dp_ex_stage_alu_r61_n136) );
  AOI21_X1 dp_ex_stage_alu_r61_U99 ( .B1(dp_ex_stage_alu_r61_n136), .B2(
        dp_ex_stage_alu_r61_n42), .A(dp_ex_stage_alu_r61_n137), .ZN(
        dp_ex_stage_alu_r61_n125) );
  NOR2_X1 dp_ex_stage_alu_r61_U98 ( .A1(dp_ex_stage_muxB_out[29]), .A2(
        dp_ex_stage_alu_r61_n101), .ZN(dp_ex_stage_alu_r61_n106) );
  NOR2_X1 dp_ex_stage_alu_r61_U97 ( .A1(dp_ex_stage_muxB_out[9]), .A2(
        dp_ex_stage_alu_r61_n13), .ZN(dp_ex_stage_alu_r61_n178) );
  AOI21_X1 dp_ex_stage_alu_r61_U96 ( .B1(dp_ex_stage_alu_r61_n178), .B2(
        dp_ex_stage_alu_r61_n79), .A(dp_ex_stage_alu_r61_n179), .ZN(
        dp_ex_stage_alu_r61_n169) );
  NAND2_X1 dp_ex_stage_alu_r61_U95 ( .A1(dp_ex_stage_muxB_out[21]), .A2(
        dp_ex_stage_alu_r61_n23), .ZN(dp_ex_stage_alu_r61_n51) );
  NAND2_X1 dp_ex_stage_alu_r61_U94 ( .A1(dp_ex_stage_alu_n45), .A2(
        dp_ex_stage_alu_r61_n65), .ZN(dp_ex_stage_alu_r61_n64) );
  NOR2_X1 dp_ex_stage_alu_r61_U93 ( .A1(dp_ex_stage_alu_n45), .A2(
        dp_ex_stage_alu_r61_n65), .ZN(dp_ex_stage_alu_r61_n198) );
  NAND2_X1 dp_ex_stage_alu_r61_U92 ( .A1(dp_ex_stage_muxB_out[9]), .A2(
        dp_ex_stage_alu_r61_n13), .ZN(dp_ex_stage_alu_r61_n88) );
  NAND2_X1 dp_ex_stage_alu_r61_U91 ( .A1(dp_ex_stage_muxB_out[15]), .A2(
        dp_ex_stage_alu_r61_n19), .ZN(dp_ex_stage_alu_r61_n92) );
  NAND2_X1 dp_ex_stage_alu_r61_U90 ( .A1(dp_ex_stage_muxB_out[22]), .A2(
        dp_ex_stage_alu_r61_n24), .ZN(dp_ex_stage_alu_r61_n42) );
  NAND2_X1 dp_ex_stage_alu_r61_U89 ( .A1(dp_ex_stage_muxA_out[2]), .A2(
        dp_ex_stage_alu_r61_n76), .ZN(dp_ex_stage_alu_r61_n184) );
  NAND2_X1 dp_ex_stage_alu_r61_U88 ( .A1(dp_ex_stage_alu_r61_n74), .A2(
        dp_ex_stage_alu_r61_n7), .ZN(dp_ex_stage_alu_r61_n183) );
  NAND2_X1 dp_ex_stage_alu_r61_U87 ( .A1(dp_ex_stage_alu_r61_n187), .A2(
        dp_ex_stage_alu_r61_n74), .ZN(dp_ex_stage_alu_r61_n185) );
  OAI211_X1 dp_ex_stage_alu_r61_U86 ( .C1(dp_ex_stage_alu_r61_n183), .C2(
        dp_ex_stage_alu_r61_n184), .A(dp_ex_stage_alu_r61_n185), .B(
        dp_ex_stage_alu_r61_n186), .ZN(dp_ex_stage_alu_r61_n182) );
  NAND2_X1 dp_ex_stage_alu_r61_U85 ( .A1(dp_ex_stage_alu_n22), .A2(
        dp_ex_stage_alu_r61_n197), .ZN(dp_ex_stage_alu_r61_n74) );
  INV_X1 dp_ex_stage_alu_r61_U84 ( .A(dp_ex_stage_muxB_out[13]), .ZN(
        dp_ex_stage_alu_r61_n180) );
  NAND2_X1 dp_ex_stage_alu_r61_U83 ( .A1(dp_ex_stage_alu_r61_n180), .A2(
        dp_ex_stage_muxA_out[13]), .ZN(dp_ex_stage_alu_r61_n161) );
  NAND2_X1 dp_ex_stage_alu_r61_U82 ( .A1(dp_ex_stage_muxB_out[16]), .A2(
        dp_ex_stage_alu_r61_n20), .ZN(dp_ex_stage_alu_r61_n93) );
  NAND2_X1 dp_ex_stage_alu_r61_U81 ( .A1(dp_ex_stage_muxB_out[10]), .A2(
        dp_ex_stage_alu_r61_n14), .ZN(dp_ex_stage_alu_r61_n79) );
  XNOR2_X1 dp_ex_stage_alu_r61_U80 ( .A(dp_ex_stage_muxB_out[31]), .B(
        dp_ex_stage_alu_r61_n31), .ZN(dp_ex_stage_alu_r61_n99) );
  NAND2_X1 dp_ex_stage_alu_r61_U79 ( .A1(dp_ex_stage_muxB_out[17]), .A2(
        dp_ex_stage_alu_r61_n21), .ZN(dp_ex_stage_alu_r61_n45) );
  NAND2_X1 dp_ex_stage_alu_r61_U78 ( .A1(dp_ex_stage_muxB_out[12]), .A2(
        dp_ex_stage_alu_r61_n16), .ZN(dp_ex_stage_alu_r61_n87) );
  INV_X1 dp_ex_stage_alu_r61_U77 ( .A(dp_ex_stage_muxB_out[23]), .ZN(
        dp_ex_stage_alu_r61_n133) );
  NAND2_X1 dp_ex_stage_alu_r61_U76 ( .A1(dp_ex_stage_muxA_out[23]), .A2(
        dp_ex_stage_alu_r61_n133), .ZN(dp_ex_stage_alu_r61_n132) );
  INV_X1 dp_ex_stage_alu_r61_U75 ( .A(dp_ex_stage_muxB_out[12]), .ZN(
        dp_ex_stage_alu_r61_n172) );
  NAND2_X1 dp_ex_stage_alu_r61_U74 ( .A1(dp_ex_stage_muxA_out[12]), .A2(
        dp_ex_stage_alu_r61_n172), .ZN(dp_ex_stage_alu_r61_n162) );
  INV_X1 dp_ex_stage_alu_r61_U73 ( .A(dp_ex_stage_muxA_out[19]), .ZN(
        dp_ex_stage_alu_r61_n214) );
  NAND2_X1 dp_ex_stage_alu_r61_U72 ( .A1(dp_ex_stage_muxB_out[19]), .A2(
        dp_ex_stage_alu_r61_n214), .ZN(dp_ex_stage_alu_r61_n43) );
  INV_X1 dp_ex_stage_alu_r61_U71 ( .A(dp_ex_stage_muxB_out[18]), .ZN(
        dp_ex_stage_alu_r61_n217) );
  NAND2_X1 dp_ex_stage_alu_r61_U70 ( .A1(dp_ex_stage_muxA_out[18]), .A2(
        dp_ex_stage_alu_r61_n217), .ZN(dp_ex_stage_alu_r61_n147) );
  INV_X1 dp_ex_stage_alu_r61_U69 ( .A(dp_ex_stage_muxB_out[24]), .ZN(
        dp_ex_stage_alu_r61_n130) );
  NAND2_X1 dp_ex_stage_alu_r61_U68 ( .A1(dp_ex_stage_muxA_out[24]), .A2(
        dp_ex_stage_alu_r61_n130), .ZN(dp_ex_stage_alu_r61_n118) );
  INV_X1 dp_ex_stage_alu_r61_U67 ( .A(dp_ex_stage_muxB_out[25]), .ZN(
        dp_ex_stage_alu_r61_n138) );
  NAND2_X1 dp_ex_stage_alu_r61_U66 ( .A1(dp_ex_stage_muxA_out[25]), .A2(
        dp_ex_stage_alu_r61_n138), .ZN(dp_ex_stage_alu_r61_n117) );
  INV_X1 dp_ex_stage_alu_r61_U65 ( .A(dp_ex_stage_muxB_out[11]), .ZN(
        dp_ex_stage_alu_r61_n175) );
  NAND2_X1 dp_ex_stage_alu_r61_U64 ( .A1(dp_ex_stage_muxA_out[11]), .A2(
        dp_ex_stage_alu_r61_n175), .ZN(dp_ex_stage_alu_r61_n174) );
  INV_X1 dp_ex_stage_alu_r61_U63 ( .A(dp_ex_stage_muxA_out[29]), .ZN(
        dp_ex_stage_alu_r61_n101) );
  INV_X1 dp_ex_stage_alu_r61_U62 ( .A(dp_ex_stage_muxA_out[30]), .ZN(
        dp_ex_stage_alu_r61_n62) );
  INV_X1 dp_ex_stage_alu_r61_U61 ( .A(dp_ex_stage_muxB_out[19]), .ZN(
        dp_ex_stage_alu_r61_n220) );
  NAND2_X1 dp_ex_stage_alu_r61_U60 ( .A1(dp_ex_stage_muxA_out[19]), .A2(
        dp_ex_stage_alu_r61_n220), .ZN(dp_ex_stage_alu_r61_n155) );
  INV_X1 dp_ex_stage_alu_r61_U59 ( .A(dp_ex_stage_muxB_out[20]), .ZN(
        dp_ex_stage_alu_r61_n135) );
  NAND4_X1 dp_ex_stage_alu_r61_U58 ( .A1(dp_ex_stage_muxA_out[20]), .A2(
        dp_ex_stage_alu_r61_n51), .A3(dp_ex_stage_alu_r61_n42), .A4(
        dp_ex_stage_alu_r61_n135), .ZN(dp_ex_stage_alu_r61_n126) );
  AOI21_X1 dp_ex_stage_alu_r61_U57 ( .B1(dp_ex_stage_alu_r61_n2), .B2(
        dp_ex_stage_alu_r61_n164), .A(dp_ex_stage_alu_r61_n165), .ZN(
        dp_ex_stage_alu_r61_n156) );
  NOR2_X1 dp_ex_stage_alu_r61_U56 ( .A1(dp_ex_stage_alu_r61_n159), .A2(
        dp_ex_stage_alu_r61_n160), .ZN(dp_ex_stage_alu_r61_n158) );
  AND3_X1 dp_ex_stage_alu_r61_U55 ( .A1(dp_ex_stage_alu_r61_n156), .A2(
        dp_ex_stage_alu_r61_n157), .A3(dp_ex_stage_alu_r61_n158), .ZN(
        dp_ex_stage_alu_r61_n140) );
  NOR2_X1 dp_ex_stage_alu_r61_U54 ( .A1(dp_ex_stage_alu_r61_n34), .A2(
        dp_ex_stage_alu_r61_n35), .ZN(dp_ex_stage_alu_r61_n33) );
  NAND2_X1 dp_ex_stage_alu_r61_U53 ( .A1(dp_ex_stage_alu_r61_n3), .A2(
        dp_ex_stage_alu_r61_n33), .ZN(dp_ex_stage_alu_N18) );
  NAND2_X1 dp_ex_stage_alu_r61_U52 ( .A1(dp_ex_stage_alu_r61_n56), .A2(
        dp_ex_stage_alu_r61_n57), .ZN(dp_ex_stage_alu_r61_n52) );
  NAND2_X1 dp_ex_stage_alu_r61_U51 ( .A1(dp_ex_stage_alu_r61_n44), .A2(
        dp_ex_stage_alu_r61_n45), .ZN(dp_ex_stage_alu_r61_n40) );
  NAND2_X1 dp_ex_stage_alu_r61_U50 ( .A1(dp_ex_stage_alu_r61_n54), .A2(
        dp_ex_stage_alu_r61_n55), .ZN(dp_ex_stage_alu_r61_n53) );
  NAND2_X1 dp_ex_stage_alu_r61_U49 ( .A1(dp_ex_stage_alu_r61_n48), .A2(
        dp_ex_stage_alu_r61_n49), .ZN(dp_ex_stage_alu_r61_n47) );
  AND2_X1 dp_ex_stage_alu_r61_U48 ( .A1(dp_ex_stage_alu_r61_n81), .A2(
        dp_ex_stage_alu_r61_n80), .ZN(dp_ex_stage_alu_r61_n5) );
  AND2_X1 dp_ex_stage_alu_r61_U47 ( .A1(dp_ex_stage_alu_r61_n5), .A2(
        dp_ex_stage_alu_r61_n79), .ZN(dp_ex_stage_alu_r61_n203) );
  NAND2_X1 dp_ex_stage_alu_r61_U46 ( .A1(dp_ex_stage_alu_r61_n85), .A2(
        dp_ex_stage_alu_r61_n94), .ZN(dp_ex_stage_alu_r61_n159) );
  NAND2_X1 dp_ex_stage_alu_r61_U45 ( .A1(dp_ex_stage_alu_r61_n50), .A2(
        dp_ex_stage_alu_r61_n51), .ZN(dp_ex_stage_alu_r61_n46) );
  NAND2_X1 dp_ex_stage_alu_r61_U44 ( .A1(dp_ex_stage_alu_r61_n42), .A2(
        dp_ex_stage_alu_r61_n43), .ZN(dp_ex_stage_alu_r61_n41) );
  NAND2_X1 dp_ex_stage_alu_r61_U43 ( .A1(dp_ex_stage_alu_r61_n73), .A2(
        dp_ex_stage_alu_r61_n74), .ZN(dp_ex_stage_alu_r61_n72) );
  NAND2_X1 dp_ex_stage_alu_r61_U42 ( .A1(dp_ex_stage_alu_r61_n75), .A2(
        dp_ex_stage_alu_r61_n76), .ZN(dp_ex_stage_alu_r61_n71) );
  NOR2_X1 dp_ex_stage_alu_r61_U41 ( .A1(dp_ex_stage_alu_r61_n71), .A2(
        dp_ex_stage_alu_r61_n72), .ZN(dp_ex_stage_alu_r61_n70) );
  NAND2_X1 dp_ex_stage_alu_r61_U40 ( .A1(dp_ex_stage_alu_r61_n93), .A2(
        dp_ex_stage_alu_r61_n94), .ZN(dp_ex_stage_alu_r61_n89) );
  NAND2_X1 dp_ex_stage_alu_r61_U39 ( .A1(dp_ex_stage_alu_r61_n91), .A2(
        dp_ex_stage_alu_r61_n92), .ZN(dp_ex_stage_alu_r61_n90) );
  NOR2_X1 dp_ex_stage_alu_r61_U38 ( .A1(dp_ex_stage_alu_r61_n89), .A2(
        dp_ex_stage_alu_r61_n90), .ZN(dp_ex_stage_alu_r61_n67) );
  NAND2_X1 dp_ex_stage_alu_r61_U37 ( .A1(dp_ex_stage_alu_r61_n87), .A2(
        dp_ex_stage_alu_r61_n88), .ZN(dp_ex_stage_alu_r61_n83) );
  NAND2_X1 dp_ex_stage_alu_r61_U36 ( .A1(dp_ex_stage_alu_r61_n85), .A2(
        dp_ex_stage_alu_r61_n86), .ZN(dp_ex_stage_alu_r61_n84) );
  NOR2_X1 dp_ex_stage_alu_r61_U35 ( .A1(dp_ex_stage_alu_r61_n83), .A2(
        dp_ex_stage_alu_r61_n84), .ZN(dp_ex_stage_alu_r61_n68) );
  AND2_X1 dp_ex_stage_alu_r61_U34 ( .A1(dp_ex_stage_alu_r61_n57), .A2(
        dp_ex_stage_alu_r61_n48), .ZN(dp_ex_stage_alu_r61_n120) );
  NAND2_X1 dp_ex_stage_alu_r61_U33 ( .A1(dp_ex_stage_alu_r61_n81), .A2(
        dp_ex_stage_alu_r61_n82), .ZN(dp_ex_stage_alu_r61_n77) );
  NAND2_X1 dp_ex_stage_alu_r61_U32 ( .A1(dp_ex_stage_alu_r61_n79), .A2(
        dp_ex_stage_alu_r61_n80), .ZN(dp_ex_stage_alu_r61_n78) );
  NOR2_X1 dp_ex_stage_alu_r61_U31 ( .A1(dp_ex_stage_alu_r61_n77), .A2(
        dp_ex_stage_alu_r61_n78), .ZN(dp_ex_stage_alu_r61_n69) );
  AND2_X1 dp_ex_stage_alu_r61_U30 ( .A1(dp_ex_stage_alu_r61_n44), .A2(
        dp_ex_stage_alu_r61_n43), .ZN(dp_ex_stage_alu_r61_n4) );
  AND2_X1 dp_ex_stage_alu_r61_U29 ( .A1(dp_ex_stage_alu_r61_n4), .A2(
        dp_ex_stage_alu_r61_n42), .ZN(dp_ex_stage_alu_r61_n213) );
  NAND2_X1 dp_ex_stage_alu_r61_U28 ( .A1(dp_ex_stage_muxA_out[22]), .A2(
        dp_ex_stage_alu_r61_n134), .ZN(dp_ex_stage_alu_r61_n131) );
  NAND2_X1 dp_ex_stage_alu_r61_U27 ( .A1(dp_ex_stage_alu_r61_n131), .A2(
        dp_ex_stage_alu_r61_n132), .ZN(dp_ex_stage_alu_r61_n128) );
  NOR2_X1 dp_ex_stage_alu_r61_U26 ( .A1(dp_ex_stage_alu_r61_n128), .A2(
        dp_ex_stage_alu_r61_n129), .ZN(dp_ex_stage_alu_r61_n127) );
  NAND2_X1 dp_ex_stage_alu_r61_U25 ( .A1(dp_ex_stage_alu_r61_n117), .A2(
        dp_ex_stage_alu_r61_n118), .ZN(dp_ex_stage_alu_r61_n116) );
  NOR2_X1 dp_ex_stage_alu_r61_U24 ( .A1(dp_ex_stage_alu_r61_n49), .A2(
        dp_ex_stage_alu_r61_n116), .ZN(dp_ex_stage_alu_r61_n115) );
  NOR2_X1 dp_ex_stage_alu_r61_U23 ( .A1(dp_ex_stage_alu_r61_n114), .A2(
        dp_ex_stage_alu_r61_n115), .ZN(dp_ex_stage_alu_r61_n108) );
  NAND2_X1 dp_ex_stage_alu_r61_U22 ( .A1(dp_ex_stage_alu_r61_n55), .A2(
        dp_ex_stage_alu_r61_n56), .ZN(dp_ex_stage_alu_r61_n103) );
  NOR2_X1 dp_ex_stage_alu_r61_U21 ( .A1(dp_ex_stage_alu_r61_n105), .A2(
        dp_ex_stage_alu_r61_n106), .ZN(dp_ex_stage_alu_r61_n104) );
  OAI21_X1 dp_ex_stage_alu_r61_U20 ( .B1(dp_ex_stage_alu_r61_n102), .B2(
        dp_ex_stage_alu_r61_n103), .A(dp_ex_stage_alu_r61_n104), .ZN(
        dp_ex_stage_alu_r61_n97) );
  NAND2_X1 dp_ex_stage_alu_r61_U19 ( .A1(dp_ex_stage_alu_r61_n63), .A2(
        dp_ex_stage_alu_r61_n64), .ZN(dp_ex_stage_alu_r61_n58) );
  NOR2_X1 dp_ex_stage_alu_r61_U18 ( .A1(dp_ex_stage_alu_r61_n58), .A2(
        dp_ex_stage_alu_r61_n59), .ZN(dp_ex_stage_alu_r61_n36) );
  AOI21_X1 dp_ex_stage_alu_r61_U17 ( .B1(dp_ex_stage_alu_r61_n186), .B2(
        dp_ex_stage_alu_r61_n207), .A(dp_ex_stage_alu_r61_n208), .ZN(
        dp_ex_stage_alu_r61_n201) );
  OAI211_X1 dp_ex_stage_alu_r61_U16 ( .C1(dp_ex_stage_alu_r61_n198), .C2(
        dp_ex_stage_alu_r61_n199), .A(dp_ex_stage_alu_r61_n200), .B(
        dp_ex_stage_alu_r61_n73), .ZN(dp_ex_stage_alu_r61_n188) );
  NOR2_X1 dp_ex_stage_alu_r61_U15 ( .A1(dp_ex_stage_alu_r61_n191), .A2(
        dp_ex_stage_alu_r61_n192), .ZN(dp_ex_stage_alu_r61_n190) );
  NAND2_X1 dp_ex_stage_alu_r61_U14 ( .A1(dp_ex_stage_alu_r61_n76), .A2(
        dp_ex_stage_alu_r61_n74), .ZN(dp_ex_stage_alu_r61_n189) );
  OAI21_X1 dp_ex_stage_alu_r61_U13 ( .B1(dp_ex_stage_alu_r61_n188), .B2(
        dp_ex_stage_alu_r61_n189), .A(dp_ex_stage_alu_r61_n190), .ZN(
        dp_ex_stage_alu_r61_n181) );
  AOI21_X1 dp_ex_stage_alu_r61_U12 ( .B1(dp_ex_stage_alu_r61_n155), .B2(
        dp_ex_stage_alu_r61_n218), .A(dp_ex_stage_alu_r61_n219), .ZN(
        dp_ex_stage_alu_r61_n211) );
  NOR2_X1 dp_ex_stage_alu_r61_U11 ( .A1(dp_ex_stage_alu_r61_n181), .A2(
        dp_ex_stage_alu_r61_n182), .ZN(dp_ex_stage_alu_r61_n167) );
  AND3_X1 dp_ex_stage_alu_r61_U10 ( .A1(dp_ex_stage_alu_r61_n169), .A2(
        dp_ex_stage_alu_r61_n170), .A3(dp_ex_stage_alu_r61_n171), .ZN(
        dp_ex_stage_alu_r61_n168) );
  AND3_X1 dp_ex_stage_alu_r61_U9 ( .A1(dp_ex_stage_alu_r61_n125), .A2(
        dp_ex_stage_alu_r61_n126), .A3(dp_ex_stage_alu_r61_n127), .ZN(
        dp_ex_stage_alu_r61_n124) );
  NOR2_X1 dp_ex_stage_alu_r61_U8 ( .A1(dp_ex_stage_alu_r61_n52), .A2(
        dp_ex_stage_alu_r61_n53), .ZN(dp_ex_stage_alu_r61_n37) );
  NOR2_X1 dp_ex_stage_alu_r61_U7 ( .A1(dp_ex_stage_alu_r61_n46), .A2(
        dp_ex_stage_alu_r61_n47), .ZN(dp_ex_stage_alu_r61_n38) );
  NOR2_X1 dp_ex_stage_alu_r61_U6 ( .A1(dp_ex_stage_alu_r61_n40), .A2(
        dp_ex_stage_alu_r61_n41), .ZN(dp_ex_stage_alu_r61_n39) );
  NAND4_X1 dp_ex_stage_alu_r61_U5 ( .A1(dp_ex_stage_alu_r61_n36), .A2(
        dp_ex_stage_alu_r61_n37), .A3(dp_ex_stage_alu_r61_n38), .A4(
        dp_ex_stage_alu_r61_n39), .ZN(dp_ex_stage_alu_r61_n35) );
  BUF_X1 dp_ex_stage_alu_r61_U4 ( .A(dp_ex_stage_alu_r61_n161), .Z(
        dp_ex_stage_alu_r61_n2) );
  INV_X1 dp_ex_stage_alu_r61_U3 ( .A(dp_ex_stage_alu_r61_n3), .ZN(
        dp_ex_stage_alu_N21) );
  AND2_X1 dp_ex_stage_alu_r61_U2 ( .A1(dp_ex_stage_alu_r61_n222), .A2(
        dp_ex_stage_alu_r61_n99), .ZN(dp_ex_stage_alu_r61_n1) );
  AND2_X1 dp_ex_stage_alu_r61_U1 ( .A1(dp_ex_stage_alu_r61_n95), .A2(
        dp_ex_stage_alu_r61_n96), .ZN(dp_ex_stage_alu_r61_n3) );
  INV_X1 dp_ex_stage_alu_r60_U318 ( .A(dp_ex_stage_alu_r60_n4), .ZN(
        dp_ex_stage_alu_r60_n306) );
  NOR2_X1 dp_ex_stage_alu_r60_U317 ( .A1(dp_ex_stage_alu_r60_n306), .A2(
        dp_ex_stage_alu_r60_n20), .ZN(dp_ex_stage_alu_r60_n305) );
  NAND3_X1 dp_ex_stage_alu_r60_U316 ( .A1(dp_ex_stage_alu_r60_n304), .A2(
        dp_ex_stage_alu_r60_n4), .A3(dp_ex_stage_alu_r60_n25), .ZN(
        dp_ex_stage_alu_r60_n301) );
  INV_X1 dp_ex_stage_alu_r60_U315 ( .A(dp_ex_stage_alu_r60_n121), .ZN(
        dp_ex_stage_alu_r60_n183) );
  INV_X1 dp_ex_stage_alu_r60_U314 ( .A(dp_ex_stage_alu_r60_n122), .ZN(
        dp_ex_stage_alu_r60_n303) );
  NOR2_X1 dp_ex_stage_alu_r60_U313 ( .A1(dp_ex_stage_alu_r60_n183), .A2(
        dp_ex_stage_alu_r60_n303), .ZN(dp_ex_stage_alu_r60_n302) );
  NAND2_X1 dp_ex_stage_alu_r60_U312 ( .A1(dp_ex_stage_alu_r60_n19), .A2(
        dp_ex_stage_alu_r60_n162), .ZN(dp_ex_stage_alu_r60_n296) );
  NAND3_X1 dp_ex_stage_alu_r60_U311 ( .A1(dp_ex_stage_alu_r60_n285), .A2(
        dp_ex_stage_alu_r60_n158), .A3(dp_ex_stage_alu_r60_n271), .ZN(
        dp_ex_stage_alu_r60_n284) );
  INV_X1 dp_ex_stage_alu_r60_U310 ( .A(dp_ex_stage_alu_r60_n151), .ZN(
        dp_ex_stage_alu_r60_n278) );
  NOR2_X1 dp_ex_stage_alu_r60_U309 ( .A1(dp_ex_stage_alu_r60_n13), .A2(
        dp_ex_stage_alu_r60_n278), .ZN(dp_ex_stage_alu_r60_n277) );
  INV_X1 dp_ex_stage_alu_r60_U308 ( .A(dp_ex_stage_alu_r60_n271), .ZN(
        dp_ex_stage_alu_r60_n272) );
  NOR2_X1 dp_ex_stage_alu_r60_U307 ( .A1(dp_ex_stage_alu_r60_n272), .A2(
        dp_ex_stage_alu_r60_n14), .ZN(dp_ex_stage_alu_r60_n270) );
  NAND3_X1 dp_ex_stage_alu_r60_U306 ( .A1(dp_ex_stage_alu_r60_n262), .A2(
        dp_ex_stage_alu_r60_n135), .A3(dp_ex_stage_alu_r60_n263), .ZN(
        dp_ex_stage_alu_r60_n261) );
  INV_X1 dp_ex_stage_alu_r60_U305 ( .A(dp_ex_stage_alu_r60_n252), .ZN(
        dp_ex_stage_alu_r60_n251) );
  NAND2_X1 dp_ex_stage_alu_r60_U304 ( .A1(dp_ex_stage_alu_r60_n251), .A2(
        dp_ex_stage_alu_r60_n121), .ZN(dp_ex_stage_alu_r60_n249) );
  NAND3_X1 dp_ex_stage_alu_r60_U303 ( .A1(dp_ex_stage_alu_r60_n245), .A2(
        dp_ex_stage_alu_r60_n109), .A3(dp_ex_stage_alu_r60_n232), .ZN(
        dp_ex_stage_alu_r60_n244) );
  INV_X1 dp_ex_stage_alu_r60_U302 ( .A(dp_ex_stage_alu_r60_n99), .ZN(
        dp_ex_stage_alu_r60_n93) );
  INV_X1 dp_ex_stage_alu_r60_U301 ( .A(dp_ex_stage_alu_r60_n226), .ZN(
        dp_ex_stage_alu_r60_n225) );
  NAND2_X1 dp_ex_stage_alu_r60_U300 ( .A1(dp_ex_stage_alu_r60_n225), .A2(
        dp_ex_stage_alu_r60_n99), .ZN(dp_ex_stage_alu_r60_n218) );
  INV_X1 dp_ex_stage_alu_r60_U299 ( .A(dp_ex_stage_alu_r60_n80), .ZN(
        dp_ex_stage_alu_r60_n220) );
  INV_X1 dp_ex_stage_alu_r60_U298 ( .A(dp_ex_stage_alu_r60_n222), .ZN(
        dp_ex_stage_alu_r60_n221) );
  OAI211_X1 dp_ex_stage_alu_r60_U297 ( .C1(dp_ex_stage_alu_r60_n12), .C2(
        dp_ex_stage_alu_r60_n218), .A(dp_ex_stage_alu_r60_n10), .B(
        dp_ex_stage_alu_r60_n219), .ZN(dp_ex_stage_alu_r60_n217) );
  NAND2_X1 dp_ex_stage_alu_r60_U296 ( .A1(dp_ex_stage_alu_r60_n21), .A2(
        dp_ex_stage_alu_r60_n84), .ZN(dp_ex_stage_alu_r60_n209) );
  INV_X1 dp_ex_stage_alu_r60_U295 ( .A(dp_ex_stage_alu_r60_n213), .ZN(
        dp_ex_stage_alu_r60_n211) );
  NAND2_X1 dp_ex_stage_alu_r60_U294 ( .A1(dp_ex_stage_alu_r60_n22), .A2(
        dp_ex_stage_alu_r60_n73), .ZN(dp_ex_stage_alu_r60_n196) );
  INV_X1 dp_ex_stage_alu_r60_U293 ( .A(dp_ex_stage_alu_r60_n201), .ZN(
        dp_ex_stage_alu_r60_n198) );
  INV_X1 dp_ex_stage_alu_r60_U292 ( .A(dp_ex_stage_alu_r60_n60), .ZN(
        dp_ex_stage_alu_r60_n199) );
  INV_X1 dp_ex_stage_alu_r60_U291 ( .A(dp_ex_stage_alu_r60_n187), .ZN(
        dp_ex_stage_alu_r60_n58) );
  NAND2_X1 dp_ex_stage_alu_r60_U290 ( .A1(dp_ex_stage_alu_r60_n67), .A2(
        dp_ex_stage_alu_r60_n61), .ZN(dp_ex_stage_alu_r60_n193) );
  NAND2_X1 dp_ex_stage_alu_r60_U289 ( .A1(dp_ex_stage_alu_r60_n191), .A2(
        dp_ex_stage_alu_r60_n192), .ZN(dp_ex_stage_alu_r60_n190) );
  INV_X1 dp_ex_stage_alu_r60_U288 ( .A(dp_ex_stage_alu_r60_n123), .ZN(
        dp_ex_stage_alu_r60_n182) );
  NOR2_X1 dp_ex_stage_alu_r60_U287 ( .A1(dp_ex_stage_alu_r60_n182), .A2(
        dp_ex_stage_alu_r60_n183), .ZN(dp_ex_stage_alu_r60_n180) );
  NAND3_X1 dp_ex_stage_alu_r60_U286 ( .A1(dp_ex_stage_alu_r60_n121), .A2(
        dp_ex_stage_alu_r60_n123), .A3(dp_ex_stage_alu_r60_n20), .ZN(
        dp_ex_stage_alu_r60_n177) );
  NAND4_X1 dp_ex_stage_alu_r60_U285 ( .A1(dp_ex_stage_alu_r60_n174), .A2(
        dp_ex_stage_alu_r60_n175), .A3(dp_ex_stage_alu_r60_n176), .A4(
        dp_ex_stage_alu_r60_n177), .ZN(dp_ex_stage_alu_r60_n100) );
  INV_X1 dp_ex_stage_alu_r60_U284 ( .A(dp_ex_stage_alu_r60_n155), .ZN(
        dp_ex_stage_alu_r60_n169) );
  NAND2_X1 dp_ex_stage_alu_r60_U283 ( .A1(dp_ex_stage_alu_r60_n169), .A2(
        dp_ex_stage_alu_r60_n170), .ZN(dp_ex_stage_alu_r60_n145) );
  INV_X1 dp_ex_stage_alu_r60_U282 ( .A(dp_ex_stage_alu_r60_n158), .ZN(
        dp_ex_stage_alu_r60_n156) );
  NAND3_X1 dp_ex_stage_alu_r60_U281 ( .A1(dp_ex_stage_alu_r60_n143), .A2(
        dp_ex_stage_alu_r60_n11), .A3(dp_ex_stage_alu_r60_n14), .ZN(
        dp_ex_stage_alu_r60_n142) );
  NAND2_X1 dp_ex_stage_alu_r60_U280 ( .A1(dp_ex_stage_alu_r60_n141), .A2(
        dp_ex_stage_alu_r60_n142), .ZN(dp_ex_stage_alu_r60_n130) );
  INV_X1 dp_ex_stage_alu_r60_U279 ( .A(dp_ex_stage_alu_r60_n11), .ZN(
        dp_ex_stage_alu_r60_n139) );
  NOR2_X1 dp_ex_stage_alu_r60_U278 ( .A1(dp_ex_stage_alu_r60_n139), .A2(
        dp_ex_stage_alu_r60_n13), .ZN(dp_ex_stage_alu_r60_n137) );
  INV_X1 dp_ex_stage_alu_r60_U277 ( .A(dp_ex_stage_alu_r60_n136), .ZN(
        dp_ex_stage_alu_r60_n134) );
  INV_X1 dp_ex_stage_alu_r60_U276 ( .A(dp_ex_stage_alu_r60_n135), .ZN(
        dp_ex_stage_alu_r60_n128) );
  NOR2_X1 dp_ex_stage_alu_r60_U275 ( .A1(dp_ex_stage_alu_r60_n134), .A2(
        dp_ex_stage_alu_r60_n128), .ZN(dp_ex_stage_alu_r60_n133) );
  INV_X1 dp_ex_stage_alu_r60_U274 ( .A(dp_ex_stage_alu_r60_n127), .ZN(
        dp_ex_stage_alu_r60_n125) );
  NAND2_X1 dp_ex_stage_alu_r60_U273 ( .A1(dp_ex_stage_alu_r60_n126), .A2(
        dp_ex_stage_alu_r60_n125), .ZN(dp_ex_stage_alu_r60_n116) );
  NAND2_X1 dp_ex_stage_alu_r60_U272 ( .A1(dp_ex_stage_alu_r60_n125), .A2(
        dp_ex_stage_alu_r60_n25), .ZN(dp_ex_stage_alu_r60_n117) );
  NAND3_X1 dp_ex_stage_alu_r60_U271 ( .A1(dp_ex_stage_alu_r60_n116), .A2(
        dp_ex_stage_alu_r60_n117), .A3(dp_ex_stage_alu_r60_n118), .ZN(
        dp_ex_stage_alu_r60_n115) );
  INV_X1 dp_ex_stage_alu_r60_U270 ( .A(dp_ex_stage_alu_r60_n110), .ZN(
        dp_ex_stage_alu_r60_n108) );
  NAND2_X1 dp_ex_stage_alu_r60_U269 ( .A1(dp_ex_stage_alu_r60_n108), .A2(
        dp_ex_stage_alu_r60_n109), .ZN(dp_ex_stage_alu_r60_n106) );
  INV_X1 dp_ex_stage_alu_r60_U268 ( .A(dp_ex_stage_alu_r60_n12), .ZN(
        dp_ex_stage_alu_r60_n97) );
  INV_X1 dp_ex_stage_alu_r60_U267 ( .A(dp_ex_stage_alu_r60_n94), .ZN(
        dp_ex_stage_alu_r60_n92) );
  NOR2_X1 dp_ex_stage_alu_r60_U266 ( .A1(dp_ex_stage_alu_r60_n92), .A2(
        dp_ex_stage_alu_r60_n93), .ZN(dp_ex_stage_alu_r60_n90) );
  NAND2_X1 dp_ex_stage_alu_r60_U265 ( .A1(dp_ex_stage_alu_r60_n21), .A2(
        dp_ex_stage_alu_r60_n80), .ZN(dp_ex_stage_alu_r60_n76) );
  INV_X1 dp_ex_stage_alu_r60_U264 ( .A(dp_ex_stage_alu_r60_n79), .ZN(
        dp_ex_stage_alu_r60_n78) );
  NAND2_X1 dp_ex_stage_alu_r60_U263 ( .A1(dp_ex_stage_alu_r60_n22), .A2(
        dp_ex_stage_alu_r60_n69), .ZN(dp_ex_stage_alu_r60_n63) );
  INV_X1 dp_ex_stage_alu_r60_U262 ( .A(dp_ex_stage_alu_r60_n68), .ZN(
        dp_ex_stage_alu_r60_n65) );
  INV_X1 dp_ex_stage_alu_r60_U261 ( .A(dp_ex_stage_alu_r60_n67), .ZN(
        dp_ex_stage_alu_r60_n66) );
  NAND2_X1 dp_ex_stage_alu_r60_U260 ( .A1(dp_ex_stage_alu_r60_n60), .A2(
        dp_ex_stage_alu_r60_n61), .ZN(dp_ex_stage_alu_r60_n59) );
  INV_X1 dp_ex_stage_alu_r60_U259 ( .A(dp_ex_stage_alu_N22), .ZN(
        dp_ex_stage_alu_N16) );
  INV_X1 dp_ex_stage_alu_r60_U258 ( .A(dp_ex_stage_muxA_out[31]), .ZN(
        dp_ex_stage_alu_r60_n53) );
  INV_X1 dp_ex_stage_alu_r60_U257 ( .A(dp_ex_stage_alu_n247), .ZN(
        dp_ex_stage_alu_r60_n52) );
  INV_X1 dp_ex_stage_alu_r60_U256 ( .A(dp_ex_stage_muxA_out[27]), .ZN(
        dp_ex_stage_alu_r60_n51) );
  INV_X1 dp_ex_stage_alu_r60_U255 ( .A(dp_ex_stage_muxA_out[26]), .ZN(
        dp_ex_stage_alu_r60_n50) );
  INV_X1 dp_ex_stage_alu_r60_U254 ( .A(dp_ex_stage_muxA_out[25]), .ZN(
        dp_ex_stage_alu_r60_n49) );
  INV_X1 dp_ex_stage_alu_r60_U253 ( .A(dp_ex_stage_muxA_out[24]), .ZN(
        dp_ex_stage_alu_r60_n48) );
  INV_X1 dp_ex_stage_alu_r60_U252 ( .A(dp_ex_stage_muxA_out[23]), .ZN(
        dp_ex_stage_alu_r60_n47) );
  INV_X1 dp_ex_stage_alu_r60_U251 ( .A(dp_ex_stage_muxA_out[22]), .ZN(
        dp_ex_stage_alu_r60_n46) );
  INV_X1 dp_ex_stage_alu_r60_U250 ( .A(dp_ex_stage_muxA_out[21]), .ZN(
        dp_ex_stage_alu_r60_n45) );
  INV_X1 dp_ex_stage_alu_r60_U249 ( .A(dp_ex_stage_muxA_out[18]), .ZN(
        dp_ex_stage_alu_r60_n44) );
  INV_X1 dp_ex_stage_alu_r60_U248 ( .A(dp_ex_stage_muxA_out[17]), .ZN(
        dp_ex_stage_alu_r60_n43) );
  INV_X1 dp_ex_stage_alu_r60_U247 ( .A(dp_ex_stage_muxA_out[16]), .ZN(
        dp_ex_stage_alu_r60_n42) );
  INV_X1 dp_ex_stage_alu_r60_U246 ( .A(dp_ex_stage_muxA_out[15]), .ZN(
        dp_ex_stage_alu_r60_n41) );
  INV_X1 dp_ex_stage_alu_r60_U245 ( .A(dp_ex_stage_muxA_out[14]), .ZN(
        dp_ex_stage_alu_r60_n40) );
  INV_X1 dp_ex_stage_alu_r60_U244 ( .A(dp_ex_stage_muxA_out[13]), .ZN(
        dp_ex_stage_alu_r60_n39) );
  INV_X1 dp_ex_stage_alu_r60_U243 ( .A(dp_ex_stage_muxA_out[12]), .ZN(
        dp_ex_stage_alu_r60_n38) );
  INV_X1 dp_ex_stage_alu_r60_U242 ( .A(dp_ex_stage_muxA_out[11]), .ZN(
        dp_ex_stage_alu_r60_n37) );
  INV_X1 dp_ex_stage_alu_r60_U241 ( .A(dp_ex_stage_muxA_out[10]), .ZN(
        dp_ex_stage_alu_r60_n36) );
  INV_X1 dp_ex_stage_alu_r60_U240 ( .A(dp_ex_stage_muxA_out[9]), .ZN(
        dp_ex_stage_alu_r60_n35) );
  INV_X1 dp_ex_stage_alu_r60_U239 ( .A(dp_ex_stage_muxA_out[8]), .ZN(
        dp_ex_stage_alu_r60_n34) );
  INV_X1 dp_ex_stage_alu_r60_U238 ( .A(dp_ex_stage_muxA_out[7]), .ZN(
        dp_ex_stage_alu_r60_n33) );
  INV_X1 dp_ex_stage_alu_r60_U237 ( .A(dp_ex_stage_muxA_out[3]), .ZN(
        dp_ex_stage_alu_r60_n32) );
  INV_X1 dp_ex_stage_alu_r60_U236 ( .A(dp_ex_stage_muxA_out[2]), .ZN(
        dp_ex_stage_alu_r60_n31) );
  INV_X1 dp_ex_stage_alu_r60_U235 ( .A(dp_ex_stage_muxB_out[4]), .ZN(
        dp_ex_stage_alu_r60_n30) );
  INV_X1 dp_ex_stage_alu_r60_U234 ( .A(dp_ex_stage_alu_n77), .ZN(
        dp_ex_stage_alu_r60_n29) );
  INV_X1 dp_ex_stage_alu_r60_U233 ( .A(dp_ex_stage_alu_n73), .ZN(
        dp_ex_stage_alu_r60_n28) );
  INV_X1 dp_ex_stage_alu_r60_U232 ( .A(dp_ex_stage_alu_n46), .ZN(
        dp_ex_stage_alu_r60_n27) );
  INV_X1 dp_ex_stage_alu_r60_U231 ( .A(dp_ex_stage_alu_n45), .ZN(
        dp_ex_stage_alu_r60_n26) );
  NAND2_X1 dp_ex_stage_alu_r60_U230 ( .A1(dp_ex_stage_alu_r60_n32), .A2(
        dp_ex_stage_alu_n77), .ZN(dp_ex_stage_alu_r60_n162) );
  NOR2_X1 dp_ex_stage_alu_r60_U229 ( .A1(dp_ex_stage_alu_r60_n266), .A2(
        dp_ex_stage_alu_r60_n267), .ZN(dp_ex_stage_alu_r60_n254) );
  NAND2_X1 dp_ex_stage_alu_r60_U228 ( .A1(dp_ex_stage_alu_r60_n256), .A2(
        dp_ex_stage_alu_r60_n257), .ZN(dp_ex_stage_alu_r60_n255) );
  AOI21_X1 dp_ex_stage_alu_r60_U227 ( .B1(dp_ex_stage_alu_r60_n253), .B2(
        dp_ex_stage_alu_r60_n254), .A(dp_ex_stage_alu_r60_n255), .ZN(
        dp_ex_stage_alu_r60_n240) );
  OAI21_X1 dp_ex_stage_alu_r60_U226 ( .B1(dp_ex_stage_alu_r60_n240), .B2(
        dp_ex_stage_alu_r60_n239), .A(dp_ex_stage_alu_r60_n241), .ZN(
        dp_ex_stage_alu_r60_n215) );
  AOI21_X1 dp_ex_stage_alu_r60_U225 ( .B1(dp_ex_stage_alu_r60_n215), .B2(
        dp_ex_stage_alu_r60_n216), .A(dp_ex_stage_alu_r60_n217), .ZN(
        dp_ex_stage_alu_r60_n208) );
  NAND2_X1 dp_ex_stage_alu_r60_U224 ( .A1(dp_ex_stage_alu_n46), .A2(
        dp_ex_stage_alu_r60_n291), .ZN(dp_ex_stage_alu_r60_n290) );
  OAI21_X1 dp_ex_stage_alu_r60_U223 ( .B1(dp_ex_stage_alu_r60_n208), .B2(
        dp_ex_stage_alu_r60_n209), .A(dp_ex_stage_alu_r60_n210), .ZN(
        dp_ex_stage_alu_r60_n204) );
  OAI21_X1 dp_ex_stage_alu_r60_U222 ( .B1(dp_ex_stage_alu_r60_n195), .B2(
        dp_ex_stage_alu_r60_n196), .A(dp_ex_stage_alu_r60_n197), .ZN(
        dp_ex_stage_alu_r60_n191) );
  INV_X1 dp_ex_stage_alu_r60_U221 ( .A(dp_ex_stage_muxA_out[4]), .ZN(
        dp_ex_stage_alu_r60_n298) );
  NAND2_X1 dp_ex_stage_alu_r60_U220 ( .A1(dp_ex_stage_muxA_out[4]), .A2(
        dp_ex_stage_alu_r60_n30), .ZN(dp_ex_stage_alu_r60_n285) );
  NAND2_X1 dp_ex_stage_alu_r60_U219 ( .A1(dp_ex_stage_alu_r60_n7), .A2(
        dp_ex_stage_alu_r60_n31), .ZN(dp_ex_stage_alu_r60_n163) );
  NAND2_X1 dp_ex_stage_alu_r60_U218 ( .A1(dp_ex_stage_muxA_out[6]), .A2(
        dp_ex_stage_alu_r60_n286), .ZN(dp_ex_stage_alu_r60_n271) );
  NAND2_X1 dp_ex_stage_alu_r60_U217 ( .A1(dp_ex_stage_muxA_out[10]), .A2(
        dp_ex_stage_alu_r60_n274), .ZN(dp_ex_stage_alu_r60_n262) );
  NOR3_X1 dp_ex_stage_alu_r60_U216 ( .A1(dp_ex_stage_alu_r60_n144), .A2(
        dp_ex_stage_alu_r60_n13), .A3(dp_ex_stage_alu_r60_n259), .ZN(
        dp_ex_stage_alu_r60_n258) );
  NOR2_X1 dp_ex_stage_alu_r60_U215 ( .A1(dp_ex_stage_alu_r60_n258), .A2(
        dp_ex_stage_alu_r60_n20), .ZN(dp_ex_stage_alu_r60_n257) );
  AOI21_X1 dp_ex_stage_alu_r60_U214 ( .B1(dp_ex_stage_alu_r60_n204), .B2(
        dp_ex_stage_alu_r60_n203), .A(dp_ex_stage_alu_r60_n205), .ZN(
        dp_ex_stage_alu_r60_n195) );
  INV_X1 dp_ex_stage_alu_r60_U213 ( .A(dp_ex_stage_muxB_out[31]), .ZN(
        dp_ex_stage_alu_r60_n315) );
  NOR2_X1 dp_ex_stage_alu_r60_U212 ( .A1(dp_ex_stage_muxB_out[31]), .A2(
        dp_ex_stage_alu_r60_n53), .ZN(dp_ex_stage_alu_r60_n185) );
  NAND2_X1 dp_ex_stage_alu_r60_U211 ( .A1(dp_ex_stage_alu_r60_n56), .A2(
        dp_ex_stage_alu_r60_n57), .ZN(dp_ex_stage_alu_r60_n55) );
  NOR2_X1 dp_ex_stage_alu_r60_U210 ( .A1(dp_ex_stage_alu_r60_n185), .A2(
        dp_ex_stage_alu_r60_n3), .ZN(dp_ex_stage_alu_r60_n54) );
  NAND2_X1 dp_ex_stage_alu_r60_U209 ( .A1(dp_ex_stage_alu_r60_n54), .A2(
        dp_ex_stage_alu_r60_n55), .ZN(dp_ex_stage_alu_N22) );
  INV_X1 dp_ex_stage_alu_r60_U208 ( .A(dp_ex_stage_muxA_out[1]), .ZN(
        dp_ex_stage_alu_r60_n291) );
  INV_X1 dp_ex_stage_alu_r60_U207 ( .A(dp_ex_stage_muxB_out[10]), .ZN(
        dp_ex_stage_alu_r60_n274) );
  INV_X1 dp_ex_stage_alu_r60_U206 ( .A(dp_ex_stage_muxA_out[30]), .ZN(
        dp_ex_stage_alu_r60_n314) );
  NOR2_X1 dp_ex_stage_alu_r60_U205 ( .A1(dp_ex_stage_muxB_out[30]), .A2(
        dp_ex_stage_alu_r60_n314), .ZN(dp_ex_stage_alu_r60_n313) );
  INV_X1 dp_ex_stage_alu_r60_U204 ( .A(dp_ex_stage_muxB_out[30]), .ZN(
        dp_ex_stage_alu_r60_n188) );
  NOR2_X1 dp_ex_stage_alu_r60_U203 ( .A1(dp_ex_stage_muxA_out[30]), .A2(
        dp_ex_stage_alu_r60_n188), .ZN(dp_ex_stage_alu_r60_n186) );
  NAND2_X1 dp_ex_stage_alu_r60_U202 ( .A1(dp_ex_stage_muxB_out[10]), .A2(
        dp_ex_stage_alu_r60_n36), .ZN(dp_ex_stage_alu_r60_n129) );
  NAND2_X1 dp_ex_stage_alu_r60_U201 ( .A1(dp_ex_stage_alu_r60_n1), .A2(
        dp_ex_stage_alu_r60_n298), .ZN(dp_ex_stage_alu_r60_n157) );
  NAND2_X1 dp_ex_stage_alu_r60_U200 ( .A1(dp_ex_stage_alu_r60_n28), .A2(
        dp_ex_stage_muxA_out[2]), .ZN(dp_ex_stage_alu_r60_n293) );
  NAND2_X1 dp_ex_stage_alu_r60_U199 ( .A1(dp_ex_stage_muxB_out[8]), .A2(
        dp_ex_stage_alu_r60_n34), .ZN(dp_ex_stage_alu_r60_n140) );
  AND2_X1 dp_ex_stage_alu_r60_U198 ( .A1(dp_ex_stage_muxB_out[11]), .A2(
        dp_ex_stage_alu_r60_n37), .ZN(dp_ex_stage_alu_r60_n25) );
  NAND2_X1 dp_ex_stage_alu_r60_U197 ( .A1(dp_ex_stage_alu_r60_n15), .A2(
        dp_ex_stage_alu_r60_n27), .ZN(dp_ex_stage_alu_r60_n168) );
  INV_X1 dp_ex_stage_alu_r60_U196 ( .A(dp_ex_stage_muxB_out[9]), .ZN(
        dp_ex_stage_alu_r60_n265) );
  NAND2_X1 dp_ex_stage_alu_r60_U195 ( .A1(dp_ex_stage_muxA_out[9]), .A2(
        dp_ex_stage_alu_r60_n265), .ZN(dp_ex_stage_alu_r60_n136) );
  INV_X1 dp_ex_stage_alu_r60_U194 ( .A(dp_ex_stage_muxB_out[8]), .ZN(
        dp_ex_stage_alu_r60_n275) );
  NAND2_X1 dp_ex_stage_alu_r60_U193 ( .A1(dp_ex_stage_muxA_out[8]), .A2(
        dp_ex_stage_alu_r60_n275), .ZN(dp_ex_stage_alu_r60_n259) );
  NAND2_X1 dp_ex_stage_alu_r60_U192 ( .A1(dp_ex_stage_alu_r60_n29), .A2(
        dp_ex_stage_muxA_out[3]), .ZN(dp_ex_stage_alu_r60_n173) );
  INV_X1 dp_ex_stage_alu_r60_U191 ( .A(dp_ex_stage_muxA_out[29]), .ZN(
        dp_ex_stage_alu_r60_n194) );
  NAND2_X1 dp_ex_stage_alu_r60_U190 ( .A1(dp_ex_stage_muxB_out[29]), .A2(
        dp_ex_stage_alu_r60_n194), .ZN(dp_ex_stage_alu_r60_n67) );
  NOR2_X1 dp_ex_stage_alu_r60_U189 ( .A1(dp_ex_stage_muxA_out[0]), .A2(
        dp_ex_stage_alu_r60_n26), .ZN(dp_ex_stage_alu_r60_n166) );
  INV_X1 dp_ex_stage_alu_r60_U188 ( .A(dp_ex_stage_muxB_out[5]), .ZN(
        dp_ex_stage_alu_r60_n287) );
  NAND2_X1 dp_ex_stage_alu_r60_U187 ( .A1(dp_ex_stage_muxA_out[5]), .A2(
        dp_ex_stage_alu_r60_n287), .ZN(dp_ex_stage_alu_r60_n158) );
  NAND2_X1 dp_ex_stage_alu_r60_U186 ( .A1(dp_ex_stage_muxB_out[23]), .A2(
        dp_ex_stage_alu_r60_n47), .ZN(dp_ex_stage_alu_r60_n84) );
  NOR2_X1 dp_ex_stage_alu_r60_U185 ( .A1(dp_ex_stage_alu_r60_n15), .A2(
        dp_ex_stage_alu_r60_n27), .ZN(dp_ex_stage_alu_r60_n167) );
  INV_X1 dp_ex_stage_alu_r60_U184 ( .A(dp_ex_stage_muxB_out[7]), .ZN(
        dp_ex_stage_alu_r60_n297) );
  NAND2_X1 dp_ex_stage_alu_r60_U183 ( .A1(dp_ex_stage_muxA_out[7]), .A2(
        dp_ex_stage_alu_r60_n297), .ZN(dp_ex_stage_alu_r60_n273) );
  NAND2_X1 dp_ex_stage_alu_r60_U182 ( .A1(dp_ex_stage_muxB_out[13]), .A2(
        dp_ex_stage_alu_r60_n39), .ZN(dp_ex_stage_alu_r60_n122) );
  NAND2_X1 dp_ex_stage_alu_r60_U181 ( .A1(dp_ex_stage_muxB_out[7]), .A2(
        dp_ex_stage_alu_r60_n33), .ZN(dp_ex_stage_alu_r60_n151) );
  NAND2_X1 dp_ex_stage_alu_r60_U180 ( .A1(dp_ex_stage_muxB_out[24]), .A2(
        dp_ex_stage_alu_r60_n48), .ZN(dp_ex_stage_alu_r60_n79) );
  NAND2_X1 dp_ex_stage_alu_r60_U179 ( .A1(dp_ex_stage_muxB_out[16]), .A2(
        dp_ex_stage_alu_r60_n42), .ZN(dp_ex_stage_alu_r60_n110) );
  NAND2_X1 dp_ex_stage_alu_r60_U178 ( .A1(dp_ex_stage_muxB_out[28]), .A2(
        dp_ex_stage_alu_r60_n52), .ZN(dp_ex_stage_alu_r60_n68) );
  NAND2_X1 dp_ex_stage_alu_r60_U177 ( .A1(dp_ex_stage_muxB_out[26]), .A2(
        dp_ex_stage_alu_r60_n50), .ZN(dp_ex_stage_alu_r60_n74) );
  NAND2_X1 dp_ex_stage_alu_r60_U176 ( .A1(dp_ex_stage_muxB_out[22]), .A2(
        dp_ex_stage_alu_r60_n46), .ZN(dp_ex_stage_alu_r60_n85) );
  NAND2_X1 dp_ex_stage_alu_r60_U175 ( .A1(dp_ex_stage_muxB_out[17]), .A2(
        dp_ex_stage_alu_r60_n43), .ZN(dp_ex_stage_alu_r60_n107) );
  INV_X1 dp_ex_stage_alu_r60_U174 ( .A(dp_ex_stage_muxA_out[5]), .ZN(
        dp_ex_stage_alu_r60_n279) );
  NAND2_X1 dp_ex_stage_alu_r60_U173 ( .A1(dp_ex_stage_muxB_out[5]), .A2(
        dp_ex_stage_alu_r60_n279), .ZN(dp_ex_stage_alu_r60_n159) );
  NAND2_X1 dp_ex_stage_alu_r60_U172 ( .A1(dp_ex_stage_muxB_out[12]), .A2(
        dp_ex_stage_alu_r60_n38), .ZN(dp_ex_stage_alu_r60_n124) );
  NAND2_X1 dp_ex_stage_alu_r60_U171 ( .A1(dp_ex_stage_alu_r60_n44), .A2(
        dp_ex_stage_muxB_out[18]), .ZN(dp_ex_stage_alu_r60_n112) );
  AND2_X1 dp_ex_stage_alu_r60_U170 ( .A1(dp_ex_stage_muxB_out[25]), .A2(
        dp_ex_stage_alu_r60_n49), .ZN(dp_ex_stage_alu_r60_n24) );
  INV_X1 dp_ex_stage_alu_r60_U169 ( .A(dp_ex_stage_muxB_out[13]), .ZN(
        dp_ex_stage_alu_r60_n307) );
  AND2_X1 dp_ex_stage_alu_r60_U168 ( .A1(dp_ex_stage_muxA_out[25]), .A2(
        dp_ex_stage_alu_r60_n212), .ZN(dp_ex_stage_alu_r60_n23) );
  NAND2_X1 dp_ex_stage_alu_r60_U167 ( .A1(dp_ex_stage_muxB_out[15]), .A2(
        dp_ex_stage_alu_r60_n41), .ZN(dp_ex_stage_alu_r60_n121) );
  INV_X1 dp_ex_stage_alu_r60_U166 ( .A(dp_ex_stage_muxB_out[22]), .ZN(
        dp_ex_stage_alu_r60_n233) );
  NAND2_X1 dp_ex_stage_alu_r60_U165 ( .A1(dp_ex_stage_muxA_out[22]), .A2(
        dp_ex_stage_alu_r60_n233), .ZN(dp_ex_stage_alu_r60_n222) );
  NAND2_X1 dp_ex_stage_alu_r60_U164 ( .A1(dp_ex_stage_muxB_out[21]), .A2(
        dp_ex_stage_alu_r60_n45), .ZN(dp_ex_stage_alu_r60_n99) );
  INV_X1 dp_ex_stage_alu_r60_U163 ( .A(dp_ex_stage_muxA_out[0]), .ZN(
        dp_ex_stage_alu_r60_n292) );
  NAND2_X1 dp_ex_stage_alu_r60_U162 ( .A1(dp_ex_stage_muxB_out[14]), .A2(
        dp_ex_stage_alu_r60_n40), .ZN(dp_ex_stage_alu_r60_n123) );
  INV_X1 dp_ex_stage_alu_r60_U161 ( .A(dp_ex_stage_muxA_out[20]), .ZN(
        dp_ex_stage_alu_r60_n234) );
  NAND2_X1 dp_ex_stage_alu_r60_U160 ( .A1(dp_ex_stage_muxB_out[20]), .A2(
        dp_ex_stage_alu_r60_n234), .ZN(dp_ex_stage_alu_r60_n94) );
  NAND2_X1 dp_ex_stage_alu_r60_U159 ( .A1(dp_ex_stage_muxB_out[27]), .A2(
        dp_ex_stage_alu_r60_n51), .ZN(dp_ex_stage_alu_r60_n73) );
  INV_X1 dp_ex_stage_alu_r60_U158 ( .A(dp_ex_stage_muxB_out[23]), .ZN(
        dp_ex_stage_alu_r60_n223) );
  NAND2_X1 dp_ex_stage_alu_r60_U157 ( .A1(dp_ex_stage_muxA_out[23]), .A2(
        dp_ex_stage_alu_r60_n223), .ZN(dp_ex_stage_alu_r60_n80) );
  INV_X1 dp_ex_stage_alu_r60_U156 ( .A(dp_ex_stage_muxB_out[28]), .ZN(
        dp_ex_stage_alu_r60_n202) );
  NAND2_X1 dp_ex_stage_alu_r60_U155 ( .A1(dp_ex_stage_alu_n247), .A2(
        dp_ex_stage_alu_r60_n202), .ZN(dp_ex_stage_alu_r60_n201) );
  INV_X1 dp_ex_stage_alu_r60_U154 ( .A(dp_ex_stage_muxB_out[27]), .ZN(
        dp_ex_stage_alu_r60_n207) );
  NAND2_X1 dp_ex_stage_alu_r60_U153 ( .A1(dp_ex_stage_muxA_out[27]), .A2(
        dp_ex_stage_alu_r60_n207), .ZN(dp_ex_stage_alu_r60_n69) );
  XNOR2_X1 dp_ex_stage_alu_r60_U152 ( .A(dp_ex_stage_muxA_out[31]), .B(
        dp_ex_stage_muxB_out[31]), .ZN(dp_ex_stage_alu_r60_n187) );
  INV_X1 dp_ex_stage_alu_r60_U151 ( .A(dp_ex_stage_muxB_out[24]), .ZN(
        dp_ex_stage_alu_r60_n214) );
  NAND2_X1 dp_ex_stage_alu_r60_U150 ( .A1(dp_ex_stage_muxA_out[24]), .A2(
        dp_ex_stage_alu_r60_n214), .ZN(dp_ex_stage_alu_r60_n213) );
  INV_X1 dp_ex_stage_alu_r60_U149 ( .A(dp_ex_stage_muxA_out[19]), .ZN(
        dp_ex_stage_alu_r60_n238) );
  NAND2_X1 dp_ex_stage_alu_r60_U148 ( .A1(dp_ex_stage_muxB_out[19]), .A2(
        dp_ex_stage_alu_r60_n238), .ZN(dp_ex_stage_alu_r60_n111) );
  INV_X1 dp_ex_stage_alu_r60_U147 ( .A(dp_ex_stage_muxB_out[17]), .ZN(
        dp_ex_stage_alu_r60_n247) );
  NAND2_X1 dp_ex_stage_alu_r60_U146 ( .A1(dp_ex_stage_muxA_out[17]), .A2(
        dp_ex_stage_alu_r60_n247), .ZN(dp_ex_stage_alu_r60_n109) );
  INV_X1 dp_ex_stage_alu_r60_U145 ( .A(dp_ex_stage_muxB_out[26]), .ZN(
        dp_ex_stage_alu_r60_n311) );
  NAND2_X1 dp_ex_stage_alu_r60_U144 ( .A1(dp_ex_stage_muxA_out[26]), .A2(
        dp_ex_stage_alu_r60_n311), .ZN(dp_ex_stage_alu_r60_n206) );
  INV_X1 dp_ex_stage_alu_r60_U143 ( .A(dp_ex_stage_muxB_out[21]), .ZN(
        dp_ex_stage_alu_r60_n224) );
  NAND2_X1 dp_ex_stage_alu_r60_U142 ( .A1(dp_ex_stage_muxA_out[21]), .A2(
        dp_ex_stage_alu_r60_n224), .ZN(dp_ex_stage_alu_r60_n89) );
  INV_X1 dp_ex_stage_alu_r60_U141 ( .A(dp_ex_stage_muxB_out[15]), .ZN(
        dp_ex_stage_alu_r60_n248) );
  NAND2_X1 dp_ex_stage_alu_r60_U140 ( .A1(dp_ex_stage_muxA_out[15]), .A2(
        dp_ex_stage_alu_r60_n248), .ZN(dp_ex_stage_alu_r60_n179) );
  INV_X1 dp_ex_stage_alu_r60_U139 ( .A(dp_ex_stage_muxB_out[11]), .ZN(
        dp_ex_stage_alu_r60_n264) );
  NAND2_X1 dp_ex_stage_alu_r60_U138 ( .A1(dp_ex_stage_muxA_out[11]), .A2(
        dp_ex_stage_alu_r60_n264), .ZN(dp_ex_stage_alu_r60_n135) );
  INV_X1 dp_ex_stage_alu_r60_U137 ( .A(dp_ex_stage_muxB_out[16]), .ZN(
        dp_ex_stage_alu_r60_n309) );
  NAND2_X1 dp_ex_stage_alu_r60_U136 ( .A1(dp_ex_stage_muxA_out[16]), .A2(
        dp_ex_stage_alu_r60_n309), .ZN(dp_ex_stage_alu_r60_n245) );
  INV_X1 dp_ex_stage_alu_r60_U135 ( .A(dp_ex_stage_muxB_out[14]), .ZN(
        dp_ex_stage_alu_r60_n310) );
  NAND2_X1 dp_ex_stage_alu_r60_U134 ( .A1(dp_ex_stage_muxA_out[14]), .A2(
        dp_ex_stage_alu_r60_n310), .ZN(dp_ex_stage_alu_r60_n252) );
  INV_X1 dp_ex_stage_alu_r60_U133 ( .A(dp_ex_stage_muxB_out[12]), .ZN(
        dp_ex_stage_alu_r60_n308) );
  NAND2_X1 dp_ex_stage_alu_r60_U132 ( .A1(dp_ex_stage_muxA_out[12]), .A2(
        dp_ex_stage_alu_r60_n308), .ZN(dp_ex_stage_alu_r60_n263) );
  INV_X1 dp_ex_stage_alu_r60_U131 ( .A(dp_ex_stage_muxB_out[29]), .ZN(
        dp_ex_stage_alu_r60_n200) );
  NAND2_X1 dp_ex_stage_alu_r60_U130 ( .A1(dp_ex_stage_muxA_out[29]), .A2(
        dp_ex_stage_alu_r60_n200), .ZN(dp_ex_stage_alu_r60_n60) );
  INV_X1 dp_ex_stage_alu_r60_U129 ( .A(dp_ex_stage_muxB_out[6]), .ZN(
        dp_ex_stage_alu_r60_n286) );
  INV_X1 dp_ex_stage_alu_r60_U128 ( .A(dp_ex_stage_muxB_out[20]), .ZN(
        dp_ex_stage_alu_r60_n235) );
  NAND2_X1 dp_ex_stage_alu_r60_U127 ( .A1(dp_ex_stage_muxA_out[20]), .A2(
        dp_ex_stage_alu_r60_n235), .ZN(dp_ex_stage_alu_r60_n226) );
  XNOR2_X1 dp_ex_stage_alu_r60_U126 ( .A(dp_ex_stage_muxA_out[30]), .B(
        dp_ex_stage_muxB_out[30]), .ZN(dp_ex_stage_alu_r60_n61) );
  INV_X1 dp_ex_stage_alu_r60_U125 ( .A(dp_ex_stage_muxB_out[18]), .ZN(
        dp_ex_stage_alu_r60_n246) );
  NAND2_X1 dp_ex_stage_alu_r60_U124 ( .A1(dp_ex_stage_muxA_out[18]), .A2(
        dp_ex_stage_alu_r60_n246), .ZN(dp_ex_stage_alu_r60_n232) );
  INV_X1 dp_ex_stage_alu_r60_U123 ( .A(dp_ex_stage_muxB_out[19]), .ZN(
        dp_ex_stage_alu_r60_n250) );
  NAND2_X1 dp_ex_stage_alu_r60_U122 ( .A1(dp_ex_stage_muxA_out[19]), .A2(
        dp_ex_stage_alu_r60_n250), .ZN(dp_ex_stage_alu_r60_n95) );
  NOR2_X1 dp_ex_stage_alu_r60_U121 ( .A1(dp_ex_stage_alu_r60_n220), .A2(
        dp_ex_stage_alu_r60_n221), .ZN(dp_ex_stage_alu_r60_n219) );
  NAND2_X1 dp_ex_stage_alu_r60_U120 ( .A1(dp_ex_stage_alu_r60_n180), .A2(
        dp_ex_stage_alu_r60_n181), .ZN(dp_ex_stage_alu_r60_n174) );
  NAND2_X1 dp_ex_stage_alu_r60_U119 ( .A1(dp_ex_stage_alu_r60_n137), .A2(
        dp_ex_stage_alu_r60_n138), .ZN(dp_ex_stage_alu_r60_n132) );
  NOR2_X1 dp_ex_stage_alu_r60_U118 ( .A1(dp_ex_stage_muxA_out[31]), .A2(
        dp_ex_stage_alu_r60_n315), .ZN(dp_ex_stage_alu_r60_n312) );
  NOR2_X1 dp_ex_stage_alu_r60_U117 ( .A1(dp_ex_stage_alu_r60_n312), .A2(
        dp_ex_stage_alu_r60_n2), .ZN(dp_ex_stage_alu_r60_n189) );
  NAND2_X1 dp_ex_stage_alu_r60_U116 ( .A1(dp_ex_stage_alu_r60_n190), .A2(
        dp_ex_stage_alu_r60_n189), .ZN(dp_ex_stage_alu_N20) );
  NAND2_X1 dp_ex_stage_alu_r60_U115 ( .A1(dp_ex_stage_alu_r60_n90), .A2(
        dp_ex_stage_alu_r60_n91), .ZN(dp_ex_stage_alu_r60_n88) );
  NOR2_X1 dp_ex_stage_alu_r60_U114 ( .A1(dp_ex_stage_alu_r60_n260), .A2(
        dp_ex_stage_alu_r60_n261), .ZN(dp_ex_stage_alu_r60_n256) );
  NAND2_X1 dp_ex_stage_alu_r60_U113 ( .A1(dp_ex_stage_alu_r60_n305), .A2(
        dp_ex_stage_alu_r60_n127), .ZN(dp_ex_stage_alu_r60_n300) );
  NAND2_X1 dp_ex_stage_alu_r60_U112 ( .A1(dp_ex_stage_alu_r60_n143), .A2(
        dp_ex_stage_alu_r60_n151), .ZN(dp_ex_stage_alu_r60_n150) );
  NAND2_X1 dp_ex_stage_alu_r60_U111 ( .A1(dp_ex_stage_alu_r60_n73), .A2(
        dp_ex_stage_alu_r60_n74), .ZN(dp_ex_stage_alu_r60_n72) );
  NAND2_X1 dp_ex_stage_alu_r60_U110 ( .A1(dp_ex_stage_alu_r60_n84), .A2(
        dp_ex_stage_alu_r60_n85), .ZN(dp_ex_stage_alu_r60_n83) );
  NAND2_X1 dp_ex_stage_alu_r60_U109 ( .A1(dp_ex_stage_alu_r60_n121), .A2(
        dp_ex_stage_alu_r60_n122), .ZN(dp_ex_stage_alu_r60_n120) );
  AND2_X1 dp_ex_stage_alu_r60_U108 ( .A1(dp_ex_stage_alu_r60_n232), .A2(
        dp_ex_stage_alu_r60_n95), .ZN(dp_ex_stage_alu_r60_n231) );
  NAND2_X1 dp_ex_stage_alu_r60_U107 ( .A1(dp_ex_stage_alu_r60_n11), .A2(
        dp_ex_stage_alu_r60_n152), .ZN(dp_ex_stage_alu_r60_n149) );
  NAND2_X1 dp_ex_stage_alu_r60_U106 ( .A1(dp_ex_stage_alu_r60_n123), .A2(
        dp_ex_stage_alu_r60_n124), .ZN(dp_ex_stage_alu_r60_n119) );
  NAND2_X1 dp_ex_stage_alu_r60_U105 ( .A1(dp_ex_stage_alu_r60_n270), .A2(
        dp_ex_stage_alu_r60_n155), .ZN(dp_ex_stage_alu_r60_n269) );
  NAND2_X1 dp_ex_stage_alu_r60_U104 ( .A1(dp_ex_stage_alu_r60_n69), .A2(
        dp_ex_stage_alu_r60_n206), .ZN(dp_ex_stage_alu_r60_n205) );
  AND2_X1 dp_ex_stage_alu_r60_U103 ( .A1(dp_ex_stage_alu_r60_n201), .A2(
        dp_ex_stage_alu_r60_n68), .ZN(dp_ex_stage_alu_r60_n22) );
  AND2_X1 dp_ex_stage_alu_r60_U102 ( .A1(dp_ex_stage_alu_r60_n213), .A2(
        dp_ex_stage_alu_r60_n79), .ZN(dp_ex_stage_alu_r60_n21) );
  NOR2_X1 dp_ex_stage_alu_r60_U101 ( .A1(dp_ex_stage_alu_r60_n128), .A2(
        dp_ex_stage_alu_r60_n129), .ZN(dp_ex_stage_alu_r60_n126) );
  NOR2_X1 dp_ex_stage_alu_r60_U100 ( .A1(dp_ex_stage_alu_r60_n24), .A2(
        dp_ex_stage_alu_r60_n184), .ZN(dp_ex_stage_alu_r60_n203) );
  NAND2_X1 dp_ex_stage_alu_r60_U99 ( .A1(dp_ex_stage_alu_r60_n95), .A2(
        dp_ex_stage_alu_r60_n232), .ZN(dp_ex_stage_alu_r60_n236) );
  NAND2_X1 dp_ex_stage_alu_r60_U98 ( .A1(dp_ex_stage_alu_r60_n229), .A2(
        dp_ex_stage_alu_r60_n230), .ZN(dp_ex_stage_alu_r60_n228) );
  OAI21_X1 dp_ex_stage_alu_r60_U97 ( .B1(dp_ex_stage_alu_r60_n107), .B2(
        dp_ex_stage_alu_r60_n236), .A(dp_ex_stage_alu_r60_n237), .ZN(
        dp_ex_stage_alu_r60_n227) );
  NOR2_X1 dp_ex_stage_alu_r60_U96 ( .A1(dp_ex_stage_alu_r60_n227), .A2(
        dp_ex_stage_alu_r60_n228), .ZN(dp_ex_stage_alu_r60_n216) );
  NOR2_X1 dp_ex_stage_alu_r60_U95 ( .A1(dp_ex_stage_alu_r60_n58), .A2(
        dp_ex_stage_alu_r60_n193), .ZN(dp_ex_stage_alu_r60_n192) );
  NAND2_X1 dp_ex_stage_alu_r60_U94 ( .A1(dp_ex_stage_alu_r60_n158), .A2(
        dp_ex_stage_alu_r60_n173), .ZN(dp_ex_stage_alu_r60_n172) );
  NOR2_X1 dp_ex_stage_alu_r60_U93 ( .A1(dp_ex_stage_alu_r60_n171), .A2(
        dp_ex_stage_alu_r60_n172), .ZN(dp_ex_stage_alu_r60_n170) );
  NAND2_X1 dp_ex_stage_alu_r60_U92 ( .A1(dp_ex_stage_alu_r60_n259), .A2(
        dp_ex_stage_alu_r60_n140), .ZN(dp_ex_stage_alu_r60_n138) );
  NOR2_X1 dp_ex_stage_alu_r60_U91 ( .A1(dp_ex_stage_alu_r60_n295), .A2(
        dp_ex_stage_alu_r60_n294), .ZN(dp_ex_stage_alu_r60_n280) );
  AOI21_X1 dp_ex_stage_alu_r60_U90 ( .B1(dp_ex_stage_alu_r60_n282), .B2(
        dp_ex_stage_alu_r60_n283), .A(dp_ex_stage_alu_r60_n284), .ZN(
        dp_ex_stage_alu_r60_n281) );
  NAND2_X1 dp_ex_stage_alu_r60_U89 ( .A1(dp_ex_stage_alu_r60_n281), .A2(
        dp_ex_stage_alu_r60_n280), .ZN(dp_ex_stage_alu_r60_n253) );
  NOR2_X1 dp_ex_stage_alu_r60_U88 ( .A1(dp_ex_stage_alu_r60_n119), .A2(
        dp_ex_stage_alu_r60_n120), .ZN(dp_ex_stage_alu_r60_n118) );
  NOR2_X1 dp_ex_stage_alu_r60_U87 ( .A1(dp_ex_stage_alu_r60_n23), .A2(
        dp_ex_stage_alu_r60_n184), .ZN(dp_ex_stage_alu_r60_n70) );
  NAND2_X1 dp_ex_stage_alu_r60_U86 ( .A1(dp_ex_stage_alu_r60_n293), .A2(
        dp_ex_stage_alu_r60_n163), .ZN(dp_ex_stage_alu_r60_n164) );
  NAND2_X1 dp_ex_stage_alu_r60_U85 ( .A1(dp_ex_stage_alu_r60_n206), .A2(
        dp_ex_stage_alu_r60_n74), .ZN(dp_ex_stage_alu_r60_n184) );
  OAI21_X1 dp_ex_stage_alu_r60_U84 ( .B1(dp_ex_stage_alu_r60_n166), .B2(
        dp_ex_stage_alu_r60_n167), .A(dp_ex_stage_alu_r60_n168), .ZN(
        dp_ex_stage_alu_r60_n165) );
  NOR2_X1 dp_ex_stage_alu_r60_U83 ( .A1(dp_ex_stage_alu_r60_n6), .A2(
        dp_ex_stage_alu_r60_n165), .ZN(dp_ex_stage_alu_r60_n160) );
  NAND2_X1 dp_ex_stage_alu_r60_U82 ( .A1(dp_ex_stage_alu_r60_n162), .A2(
        dp_ex_stage_alu_r60_n163), .ZN(dp_ex_stage_alu_r60_n161) );
  NOR2_X1 dp_ex_stage_alu_r60_U81 ( .A1(dp_ex_stage_alu_r60_n160), .A2(
        dp_ex_stage_alu_r60_n161), .ZN(dp_ex_stage_alu_r60_n146) );
  NOR2_X1 dp_ex_stage_alu_r60_U80 ( .A1(dp_ex_stage_alu_r60_n5), .A2(
        dp_ex_stage_alu_r60_n136), .ZN(dp_ex_stage_alu_r60_n260) );
  NOR2_X1 dp_ex_stage_alu_r60_U79 ( .A1(dp_ex_stage_alu_r60_n171), .A2(
        dp_ex_stage_alu_r60_n173), .ZN(dp_ex_stage_alu_r60_n294) );
  NOR2_X1 dp_ex_stage_alu_r60_U78 ( .A1(dp_ex_stage_alu_r60_n159), .A2(
        dp_ex_stage_alu_r60_n9), .ZN(dp_ex_stage_alu_r60_n153) );
  NOR2_X1 dp_ex_stage_alu_r60_U77 ( .A1(dp_ex_stage_alu_r60_n58), .A2(
        dp_ex_stage_alu_r60_n59), .ZN(dp_ex_stage_alu_r60_n57) );
  NAND2_X1 dp_ex_stage_alu_r60_U76 ( .A1(dp_ex_stage_alu_r60_n290), .A2(
        dp_ex_stage_alu_r60_n162), .ZN(dp_ex_stage_alu_r60_n289) );
  NOR2_X1 dp_ex_stage_alu_r60_U75 ( .A1(dp_ex_stage_alu_r60_n288), .A2(
        dp_ex_stage_alu_r60_n289), .ZN(dp_ex_stage_alu_r60_n283) );
  AND2_X1 dp_ex_stage_alu_r60_U74 ( .A1(dp_ex_stage_alu_r60_n179), .A2(
        dp_ex_stage_alu_r60_n109), .ZN(dp_ex_stage_alu_r60_n175) );
  NAND2_X1 dp_ex_stage_alu_r60_U73 ( .A1(dp_ex_stage_alu_r60_n99), .A2(
        dp_ex_stage_alu_r60_n94), .ZN(dp_ex_stage_alu_r60_n96) );
  NAND2_X1 dp_ex_stage_alu_r60_U72 ( .A1(dp_ex_stage_alu_r60_n88), .A2(
        dp_ex_stage_alu_r60_n89), .ZN(dp_ex_stage_alu_r60_n87) );
  OAI21_X1 dp_ex_stage_alu_r60_U71 ( .B1(dp_ex_stage_alu_r60_n95), .B2(
        dp_ex_stage_alu_r60_n96), .A(dp_ex_stage_alu_r60_n97), .ZN(
        dp_ex_stage_alu_r60_n86) );
  NOR2_X1 dp_ex_stage_alu_r60_U70 ( .A1(dp_ex_stage_alu_r60_n86), .A2(
        dp_ex_stage_alu_r60_n87), .ZN(dp_ex_stage_alu_r60_n82) );
  NAND2_X1 dp_ex_stage_alu_r60_U69 ( .A1(dp_ex_stage_alu_r60_n252), .A2(
        dp_ex_stage_alu_r60_n123), .ZN(dp_ex_stage_alu_r60_n181) );
  NAND2_X1 dp_ex_stage_alu_r60_U68 ( .A1(dp_ex_stage_alu_r60_n273), .A2(
        dp_ex_stage_alu_r60_n8), .ZN(dp_ex_stage_alu_r60_n276) );
  NAND2_X1 dp_ex_stage_alu_r60_U67 ( .A1(dp_ex_stage_alu_r60_n269), .A2(
        dp_ex_stage_alu_r60_n268), .ZN(dp_ex_stage_alu_r60_n267) );
  OAI21_X1 dp_ex_stage_alu_r60_U66 ( .B1(dp_ex_stage_alu_r60_n159), .B2(
        dp_ex_stage_alu_r60_n276), .A(dp_ex_stage_alu_r60_n277), .ZN(
        dp_ex_stage_alu_r60_n266) );
  NAND2_X1 dp_ex_stage_alu_r60_U65 ( .A1(dp_ex_stage_alu_r60_n226), .A2(
        dp_ex_stage_alu_r60_n94), .ZN(dp_ex_stage_alu_r60_n91) );
  NAND4_X1 dp_ex_stage_alu_r60_U64 ( .A1(dp_ex_stage_alu_r60_n99), .A2(
        dp_ex_stage_alu_r60_n111), .A3(dp_ex_stage_alu_r60_n94), .A4(
        dp_ex_stage_alu_r60_n112), .ZN(dp_ex_stage_alu_r60_n103) );
  NOR2_X1 dp_ex_stage_alu_r60_U63 ( .A1(dp_ex_stage_alu_r60_n178), .A2(
        dp_ex_stage_alu_r60_n179), .ZN(dp_ex_stage_alu_r60_n243) );
  AOI21_X1 dp_ex_stage_alu_r60_U62 ( .B1(dp_ex_stage_alu_r60_n70), .B2(
        dp_ex_stage_alu_r60_n71), .A(dp_ex_stage_alu_r60_n72), .ZN(
        dp_ex_stage_alu_r60_n62) );
  NOR2_X1 dp_ex_stage_alu_r60_U61 ( .A1(dp_ex_stage_alu_r60_n65), .A2(
        dp_ex_stage_alu_r60_n66), .ZN(dp_ex_stage_alu_r60_n64) );
  OAI21_X1 dp_ex_stage_alu_r60_U60 ( .B1(dp_ex_stage_alu_r60_n62), .B2(
        dp_ex_stage_alu_r60_n63), .A(dp_ex_stage_alu_r60_n64), .ZN(
        dp_ex_stage_alu_r60_n56) );
  NAND2_X1 dp_ex_stage_alu_r60_U59 ( .A1(dp_ex_stage_alu_r60_n4), .A2(
        dp_ex_stage_alu_r60_n124), .ZN(dp_ex_stage_alu_r60_n127) );
  NAND2_X1 dp_ex_stage_alu_r60_U58 ( .A1(dp_ex_stage_alu_r60_n222), .A2(
        dp_ex_stage_alu_r60_n85), .ZN(dp_ex_stage_alu_r60_n98) );
  OAI21_X1 dp_ex_stage_alu_r60_U57 ( .B1(dp_ex_stage_alu_r60_n296), .B2(
        dp_ex_stage_alu_r60_n171), .A(dp_ex_stage_alu_r60_n273), .ZN(
        dp_ex_stage_alu_r60_n295) );
  AOI21_X1 dp_ex_stage_alu_r60_U56 ( .B1(dp_ex_stage_alu_r60_n81), .B2(
        dp_ex_stage_alu_r60_n82), .A(dp_ex_stage_alu_r60_n83), .ZN(
        dp_ex_stage_alu_r60_n75) );
  NOR2_X1 dp_ex_stage_alu_r60_U55 ( .A1(dp_ex_stage_alu_r60_n78), .A2(
        dp_ex_stage_alu_r60_n24), .ZN(dp_ex_stage_alu_r60_n77) );
  OAI21_X1 dp_ex_stage_alu_r60_U54 ( .B1(dp_ex_stage_alu_r60_n75), .B2(
        dp_ex_stage_alu_r60_n76), .A(dp_ex_stage_alu_r60_n77), .ZN(
        dp_ex_stage_alu_r60_n71) );
  NOR2_X1 dp_ex_stage_alu_r60_U53 ( .A1(dp_ex_stage_alu_r60_n198), .A2(
        dp_ex_stage_alu_r60_n199), .ZN(dp_ex_stage_alu_r60_n197) );
  OAI21_X1 dp_ex_stage_alu_r60_U52 ( .B1(dp_ex_stage_alu_r60_n178), .B2(
        dp_ex_stage_alu_r60_n249), .A(dp_ex_stage_alu_r60_n95), .ZN(
        dp_ex_stage_alu_r60_n242) );
  NOR2_X1 dp_ex_stage_alu_r60_U51 ( .A1(dp_ex_stage_alu_r60_n211), .A2(
        dp_ex_stage_alu_r60_n23), .ZN(dp_ex_stage_alu_r60_n210) );
  NAND2_X1 dp_ex_stage_alu_r60_U50 ( .A1(dp_ex_stage_alu_r60_n262), .A2(
        dp_ex_stage_alu_r60_n129), .ZN(dp_ex_stage_alu_r60_n144) );
  NAND2_X1 dp_ex_stage_alu_r60_U49 ( .A1(dp_ex_stage_alu_r60_n271), .A2(
        dp_ex_stage_alu_r60_n152), .ZN(dp_ex_stage_alu_r60_n155) );
  NAND2_X1 dp_ex_stage_alu_r60_U48 ( .A1(dp_ex_stage_alu_r60_n285), .A2(
        dp_ex_stage_alu_r60_n157), .ZN(dp_ex_stage_alu_r60_n171) );
  NAND2_X1 dp_ex_stage_alu_r60_U47 ( .A1(dp_ex_stage_alu_r60_n245), .A2(
        dp_ex_stage_alu_r60_n110), .ZN(dp_ex_stage_alu_r60_n178) );
  NAND2_X1 dp_ex_stage_alu_r60_U46 ( .A1(dp_ex_stage_alu_r60_n112), .A2(
        dp_ex_stage_alu_r60_n232), .ZN(dp_ex_stage_alu_r60_n105) );
  NOR3_X1 dp_ex_stage_alu_r60_U45 ( .A1(dp_ex_stage_alu_r60_n156), .A2(
        dp_ex_stage_alu_r60_n155), .A3(dp_ex_stage_alu_r60_n157), .ZN(
        dp_ex_stage_alu_r60_n154) );
  OAI22_X1 dp_ex_stage_alu_r60_U44 ( .A1(dp_ex_stage_alu_r60_n105), .A2(
        dp_ex_stage_alu_r60_n106), .B1(dp_ex_stage_alu_r60_n107), .B2(
        dp_ex_stage_alu_r60_n105), .ZN(dp_ex_stage_alu_r60_n104) );
  NOR2_X1 dp_ex_stage_alu_r60_U43 ( .A1(dp_ex_stage_alu_r60_n127), .A2(
        dp_ex_stage_alu_r60_n5), .ZN(dp_ex_stage_alu_r60_n141) );
  NOR2_X1 dp_ex_stage_alu_r60_U42 ( .A1(dp_ex_stage_alu_r60_n105), .A2(
        dp_ex_stage_alu_r60_n178), .ZN(dp_ex_stage_alu_r60_n176) );
  NOR2_X1 dp_ex_stage_alu_r60_U41 ( .A1(dp_ex_stage_alu_r60_n181), .A2(
        dp_ex_stage_alu_r60_n178), .ZN(dp_ex_stage_alu_r60_n299) );
  NOR2_X1 dp_ex_stage_alu_r60_U40 ( .A1(dp_ex_stage_alu_r60_n138), .A2(
        dp_ex_stage_alu_r60_n144), .ZN(dp_ex_stage_alu_r60_n268) );
  NOR2_X1 dp_ex_stage_alu_r60_U39 ( .A1(dp_ex_stage_alu_r60_n91), .A2(
        dp_ex_stage_alu_r60_n98), .ZN(dp_ex_stage_alu_r60_n229) );
  NOR2_X1 dp_ex_stage_alu_r60_U38 ( .A1(dp_ex_stage_alu_r60_n164), .A2(
        dp_ex_stage_alu_r60_n171), .ZN(dp_ex_stage_alu_r60_n282) );
  NAND2_X1 dp_ex_stage_alu_r60_U37 ( .A1(dp_ex_stage_alu_r60_n132), .A2(
        dp_ex_stage_alu_r60_n133), .ZN(dp_ex_stage_alu_r60_n131) );
  NOR2_X1 dp_ex_stage_alu_r60_U36 ( .A1(dp_ex_stage_alu_r60_n130), .A2(
        dp_ex_stage_alu_r60_n131), .ZN(dp_ex_stage_alu_r60_n114) );
  AOI21_X1 dp_ex_stage_alu_r60_U35 ( .B1(dp_ex_stage_alu_r60_n113), .B2(
        dp_ex_stage_alu_r60_n114), .A(dp_ex_stage_alu_r60_n115), .ZN(
        dp_ex_stage_alu_r60_n101) );
  NOR2_X1 dp_ex_stage_alu_r60_U34 ( .A1(dp_ex_stage_alu_r60_n103), .A2(
        dp_ex_stage_alu_r60_n104), .ZN(dp_ex_stage_alu_r60_n102) );
  OAI21_X1 dp_ex_stage_alu_r60_U33 ( .B1(dp_ex_stage_alu_r60_n100), .B2(
        dp_ex_stage_alu_r60_n101), .A(dp_ex_stage_alu_r60_n102), .ZN(
        dp_ex_stage_alu_r60_n81) );
  NAND4_X1 dp_ex_stage_alu_r60_U32 ( .A1(dp_ex_stage_alu_r60_n299), .A2(
        dp_ex_stage_alu_r60_n300), .A3(dp_ex_stage_alu_r60_n301), .A4(
        dp_ex_stage_alu_r60_n302), .ZN(dp_ex_stage_alu_r60_n239) );
  NOR3_X1 dp_ex_stage_alu_r60_U31 ( .A1(dp_ex_stage_alu_r60_n242), .A2(
        dp_ex_stage_alu_r60_n243), .A3(dp_ex_stage_alu_r60_n244), .ZN(
        dp_ex_stage_alu_r60_n241) );
  NOR2_X1 dp_ex_stage_alu_r60_U30 ( .A1(dp_ex_stage_alu_r60_n153), .A2(
        dp_ex_stage_alu_r60_n154), .ZN(dp_ex_stage_alu_r60_n147) );
  NOR2_X1 dp_ex_stage_alu_r60_U29 ( .A1(dp_ex_stage_alu_r60_n149), .A2(
        dp_ex_stage_alu_r60_n150), .ZN(dp_ex_stage_alu_r60_n148) );
  OAI211_X1 dp_ex_stage_alu_r60_U28 ( .C1(dp_ex_stage_alu_r60_n145), .C2(
        dp_ex_stage_alu_r60_n146), .A(dp_ex_stage_alu_r60_n147), .B(
        dp_ex_stage_alu_r60_n148), .ZN(dp_ex_stage_alu_r60_n113) );
  AND2_X1 dp_ex_stage_alu_r60_U27 ( .A1(dp_ex_stage_muxA_out[13]), .A2(
        dp_ex_stage_alu_r60_n307), .ZN(dp_ex_stage_alu_r60_n20) );
  AND2_X1 dp_ex_stage_alu_r60_U26 ( .A1(dp_ex_stage_muxA_out[2]), .A2(
        dp_ex_stage_alu_r60_n28), .ZN(dp_ex_stage_alu_r60_n19) );
  AND2_X1 dp_ex_stage_alu_r60_U25 ( .A1(dp_ex_stage_alu_r60_n190), .A2(
        dp_ex_stage_alu_r60_n189), .ZN(dp_ex_stage_alu_N17) );
  OR2_X1 dp_ex_stage_alu_r60_U24 ( .A1(dp_ex_stage_alu_n46), .A2(
        dp_ex_stage_alu_r60_n291), .ZN(dp_ex_stage_alu_r60_n17) );
  OR2_X1 dp_ex_stage_alu_r60_U23 ( .A1(dp_ex_stage_alu_n45), .A2(
        dp_ex_stage_alu_r60_n292), .ZN(dp_ex_stage_alu_r60_n16) );
  AND2_X1 dp_ex_stage_alu_r60_U22 ( .A1(dp_ex_stage_alu_r60_n16), .A2(
        dp_ex_stage_alu_r60_n17), .ZN(dp_ex_stage_alu_r60_n288) );
  CLKBUF_X1 dp_ex_stage_alu_r60_U21 ( .A(dp_ex_stage_muxA_out[1]), .Z(
        dp_ex_stage_alu_r60_n15) );
  AND2_X1 dp_ex_stage_alu_r60_U20 ( .A1(dp_ex_stage_muxA_out[7]), .A2(
        dp_ex_stage_alu_r60_n297), .ZN(dp_ex_stage_alu_r60_n14) );
  AND2_X2 dp_ex_stage_alu_r60_U19 ( .A1(dp_ex_stage_muxB_out[9]), .A2(
        dp_ex_stage_alu_r60_n35), .ZN(dp_ex_stage_alu_r60_n13) );
  OR2_X1 dp_ex_stage_alu_r60_U18 ( .A1(dp_ex_stage_alu_r60_n286), .A2(
        dp_ex_stage_muxA_out[6]), .ZN(dp_ex_stage_alu_r60_n152) );
  CLKBUF_X1 dp_ex_stage_alu_r60_U17 ( .A(dp_ex_stage_alu_r60_n98), .Z(
        dp_ex_stage_alu_r60_n12) );
  CLKBUF_X1 dp_ex_stage_alu_r60_U16 ( .A(dp_ex_stage_alu_r60_n140), .Z(
        dp_ex_stage_alu_r60_n11) );
  OR2_X1 dp_ex_stage_alu_r60_U15 ( .A1(dp_ex_stage_alu_r60_n98), .A2(
        dp_ex_stage_alu_r60_n89), .ZN(dp_ex_stage_alu_r60_n10) );
  AND2_X1 dp_ex_stage_alu_r60_U14 ( .A1(dp_ex_stage_alu_r60_n99), .A2(
        dp_ex_stage_alu_r60_n111), .ZN(dp_ex_stage_alu_r60_n237) );
  INV_X1 dp_ex_stage_alu_r60_U13 ( .A(dp_ex_stage_alu_r60_n169), .ZN(
        dp_ex_stage_alu_r60_n9) );
  BUF_X1 dp_ex_stage_alu_r60_U12 ( .A(dp_ex_stage_alu_r60_n271), .Z(
        dp_ex_stage_alu_r60_n8) );
  CLKBUF_X1 dp_ex_stage_alu_r60_U11 ( .A(dp_ex_stage_alu_r60_n164), .Z(
        dp_ex_stage_alu_r60_n6) );
  NAND2_X1 dp_ex_stage_alu_r60_U10 ( .A1(dp_ex_stage_alu_r60_n262), .A2(
        dp_ex_stage_alu_r60_n129), .ZN(dp_ex_stage_alu_r60_n5) );
  NAND2_X1 dp_ex_stage_alu_r60_U9 ( .A1(dp_ex_stage_muxA_out[12]), .A2(
        dp_ex_stage_alu_r60_n308), .ZN(dp_ex_stage_alu_r60_n4) );
  CLKBUF_X1 dp_ex_stage_alu_r60_U8 ( .A(dp_ex_stage_alu_n73), .Z(
        dp_ex_stage_alu_r60_n7) );
  AND2_X1 dp_ex_stage_alu_r60_U7 ( .A1(dp_ex_stage_alu_r60_n186), .A2(
        dp_ex_stage_alu_r60_n187), .ZN(dp_ex_stage_alu_r60_n3) );
  AND2_X1 dp_ex_stage_alu_r60_U6 ( .A1(dp_ex_stage_alu_r60_n313), .A2(
        dp_ex_stage_alu_r60_n187), .ZN(dp_ex_stage_alu_r60_n2) );
  INV_X1 dp_ex_stage_alu_r60_U5 ( .A(dp_ex_stage_muxB_out[25]), .ZN(
        dp_ex_stage_alu_r60_n212) );
  NAND2_X1 dp_ex_stage_alu_r60_U4 ( .A1(dp_ex_stage_alu_r60_n231), .A2(
        dp_ex_stage_alu_r60_n105), .ZN(dp_ex_stage_alu_r60_n230) );
  INV_X1 dp_ex_stage_alu_r60_U3 ( .A(dp_ex_stage_alu_r60_n13), .ZN(
        dp_ex_stage_alu_r60_n143) );
  INV_X1 dp_ex_stage_alu_r60_U2 ( .A(dp_ex_stage_alu_r60_n20), .ZN(
        dp_ex_stage_alu_r60_n304) );
  CLKBUF_X1 dp_ex_stage_alu_r60_U1 ( .A(dp_ex_stage_muxB_out[4]), .Z(
        dp_ex_stage_alu_r60_n1) );
endmodule

