
module DLX ( CLK, RST, IRAM_ADDRESS, IRAM_ISSUE, IRAM_READY, IRAM_DATA, 
        DRAM_ADDRESS, DRAM_ISSUE, DRAM_READNOTWRITE, DRAM_READY, DRAM_DATA );
  output [31:0] IRAM_ADDRESS;
  input [31:0] IRAM_DATA;
  output [31:0] DRAM_ADDRESS;
  inout [31:0] DRAM_DATA;
  input CLK, RST, IRAM_READY, DRAM_READY;
  output IRAM_ISSUE, DRAM_ISSUE, DRAM_READNOTWRITE;
  wire   pipe_if_id_en_i, pipe_clear_n_i, rf_spill_i, rf_fill_i, rf_rs1_en_i,
         rf_rs2_en_i, imm_isoff_i, imm_uns_i, reg31_sel_i, regrd_sel_i,
         muxA_sel_i, muxB_sel_i, is_zero_i, mem_in_en_i, npc_wb_en_i,
         jump_en_i, pc_latch_en_i, wb_mux_sel_i, rf_we_i, \CU_I/n272 ,
         \CU_I/n271 , \CU_I/n270 , \CU_I/n269 , \CU_I/n268 , \CU_I/n267 ,
         \CU_I/n266 , \CU_I/n265 , \CU_I/n264 , \CU_I/n263 , \CU_I/n262 ,
         \CU_I/n261 , \CU_I/n260 , \CU_I/n259 , \CU_I/n258 , \CU_I/n257 ,
         \CU_I/n256 , \CU_I/n255 , \CU_I/n76 , \CU_I/n75 , \CU_I/n74 ,
         \CU_I/n73 , \CU_I/n72 , \CU_I/n71 , \CU_I/n70 , \CU_I/n69 ,
         \CU_I/n68 , \CU_I/n67 , \CU_I/n66 , \CU_I/n65 , \CU_I/n64 ,
         \CU_I/n63 , \CU_I/n62 , \CU_I/n61 , \CU_I/n60 , \CU_I/n59 ,
         \CU_I/n58 , \CU_I/n57 , \CU_I/n56 , \CU_I/n54 , \CU_I/n53 ,
         \CU_I/n52 , \CU_I/n51 , \CU_I/n50 , \CU_I/n49 , \CU_I/n48 ,
         \CU_I/n46 , \CU_I/n45 , \CU_I/n44 , \CU_I/n43 , \CU_I/n42 ,
         \CU_I/n41 , \CU_I/n40 , \CU_I/n29 , \CU_I/n28 , \CU_I/n26 ,
         \CU_I/n25 , \CU_I/n24 , \CU_I/n20 , \CU_I/n18 , \CU_I/n14 , \CU_I/n1 ,
         \CU_I/n254 , \CU_I/n253 , \CU_I/n252 , \CU_I/n251 , \CU_I/n250 ,
         \CU_I/n249 , \CU_I/n248 , \CU_I/n247 , \CU_I/n246 , \CU_I/n245 ,
         \CU_I/n244 , \CU_I/n243 , \CU_I/n242 , \CU_I/n241 , \CU_I/n240 ,
         \CU_I/n239 , \CU_I/n238 , \CU_I/n237 , \CU_I/n236 , \CU_I/n235 ,
         \CU_I/n234 , \CU_I/n233 , \CU_I/n232 , \CU_I/n231 , \CU_I/n230 ,
         \CU_I/n229 , \CU_I/n228 , \CU_I/n227 , \CU_I/n226 , \CU_I/n225 ,
         \CU_I/n224 , \CU_I/n223 , \CU_I/n222 , \CU_I/n221 , \CU_I/n220 ,
         \CU_I/n219 , \CU_I/n218 , \CU_I/n217 , \CU_I/n216 , \CU_I/n215 ,
         \CU_I/n214 , \CU_I/n213 , \CU_I/n212 , \CU_I/n211 , \CU_I/n210 ,
         \CU_I/n209 , \CU_I/n208 , \CU_I/n207 , \CU_I/n206 , \CU_I/n205 ,
         \CU_I/n204 , \CU_I/n203 , \CU_I/n202 , \CU_I/n201 , \CU_I/n200 ,
         \CU_I/n199 , \CU_I/n198 , \CU_I/n197 , \CU_I/n196 , \CU_I/n195 ,
         \CU_I/n194 , \CU_I/n193 , \CU_I/n192 , \CU_I/n191 , \CU_I/n190 ,
         \CU_I/n189 , \CU_I/n188 , \CU_I/n187 , \CU_I/n186 , \CU_I/n185 ,
         \CU_I/n184 , \CU_I/n183 , \CU_I/n182 , \CU_I/n181 , \CU_I/n180 ,
         \CU_I/n179 , \CU_I/n178 , \CU_I/n177 , \CU_I/n176 , \CU_I/n175 ,
         \CU_I/n174 , \CU_I/n173 , \CU_I/n172 , \CU_I/n171 , \CU_I/n170 ,
         \CU_I/n169 , \CU_I/n168 , \CU_I/n167 , \CU_I/n166 , \CU_I/n165 ,
         \CU_I/n164 , \CU_I/n163 , \CU_I/n162 , \CU_I/n161 , \CU_I/n160 ,
         \CU_I/n159 , \CU_I/n158 , \CU_I/n157 , \CU_I/n156 , \CU_I/n155 ,
         \CU_I/n154 , \CU_I/n153 , \CU_I/n152 , \CU_I/n151 , \CU_I/n150 ,
         \CU_I/n149 , \CU_I/n148 , \CU_I/n147 , \CU_I/n146 , \CU_I/n145 ,
         \CU_I/n144 , \CU_I/n143 , \CU_I/n142 , \CU_I/n141 , \CU_I/n140 ,
         \CU_I/n139 , \CU_I/n138 , \CU_I/n137 , \CU_I/n136 , \CU_I/n135 ,
         \CU_I/n134 , \CU_I/n133 , \CU_I/n132 , \CU_I/n131 , \CU_I/n130 ,
         \CU_I/n129 , \CU_I/n128 , \CU_I/n127 , \CU_I/n126 , \CU_I/n125 ,
         \CU_I/n124 , \CU_I/n123 , \CU_I/n122 , \CU_I/n121 , \CU_I/n120 ,
         \CU_I/n119 , \CU_I/n118 , \CU_I/n117 , \CU_I/n116 , \CU_I/n115 ,
         \CU_I/n114 , \CU_I/n113 , \CU_I/n112 , \CU_I/n111 , \CU_I/n110 ,
         \CU_I/n109 , \CU_I/n108 , \CU_I/n107 , \CU_I/n106 , \CU_I/n105 ,
         \CU_I/n104 , \CU_I/n103 , \CU_I/n102 , \CU_I/n101 , \CU_I/n100 ,
         \CU_I/n99 , \CU_I/n98 , \CU_I/n97 , \CU_I/n96 , \CU_I/n95 ,
         \CU_I/n94 , \CU_I/n93 , \CU_I/n92 , \CU_I/n91 , \CU_I/n90 ,
         \CU_I/n89 , \CU_I/n88 , \CU_I/n87 , \CU_I/n86 , \CU_I/n85 ,
         \CU_I/n84 , \CU_I/n83 , \CU_I/n82 , \CU_I/n81 , \CU_I/n80 ,
         \CU_I/n79 , \CU_I/n78 , \CU_I/n77 , \CU_I/n37 , \CU_I/n36 ,
         \CU_I/n35 , \CU_I/n34 , \CU_I/n33 , \CU_I/n32 , \CU_I/n31 ,
         \CU_I/n30 , \CU_I/n27 , \CU_I/n23 , \CU_I/n22 , \CU_I/n21 ,
         \CU_I/n19 , \CU_I/n17 , \CU_I/n16 , \CU_I/n15 , \CU_I/n13 ,
         \CU_I/n12 , \CU_I/n11 , \CU_I/n10 , \CU_I/n9 , \CU_I/n8 , \CU_I/n7 ,
         \CU_I/n6 , \CU_I/n5 , \CU_I/n4 , \CU_I/n3 , \CU_I/n2 , \CU_I/cw3[4] ,
         \CU_I/cw3[5] , \CU_I/cw1[1] , \CU_I/n273 , \dp/n1027 , \dp/n1026 ,
         \dp/n1025 , \dp/n1024 , \dp/n1023 , \dp/n1022 , \dp/n1021 ,
         \dp/n1020 , \dp/n1019 , \dp/n1018 , \dp/n1017 , \dp/n1016 , \dp/n648 ,
         \dp/n647 , \dp/n646 , \dp/n645 , \dp/n644 , \dp/n643 , \dp/n642 ,
         \dp/n641 , \dp/n640 , \dp/n639 , \dp/n638 , \dp/n637 , \dp/n636 ,
         \dp/n635 , \dp/n634 , \dp/n633 , \dp/n632 , \dp/n631 , \dp/n630 ,
         \dp/n629 , \dp/n628 , \dp/n627 , \dp/n626 , \dp/n625 , \dp/n624 ,
         \dp/n623 , \dp/n622 , \dp/n621 , \dp/n620 , \dp/n619 , \dp/n618 ,
         \dp/n617 , \dp/n616 , \dp/n615 , \dp/n614 , \dp/n613 , \dp/n612 ,
         \dp/n611 , \dp/n610 , \dp/n609 , \dp/n608 , \dp/n607 , \dp/n606 ,
         \dp/n605 , \dp/n604 , \dp/n603 , \dp/n602 , \dp/n601 , \dp/n600 ,
         \dp/n599 , \dp/n598 , \dp/n597 , \dp/n596 , \dp/n595 , \dp/n594 ,
         \dp/n593 , \dp/n592 , \dp/n591 , \dp/n590 , \dp/n589 , \dp/n588 ,
         \dp/n587 , \dp/n586 , \dp/n585 , \dp/n584 , \dp/n525 , \dp/n523 ,
         \dp/n521 , \dp/n519 , \dp/n517 , \dp/n413 , \dp/n412 , \dp/n411 ,
         \dp/n410 , \dp/n409 , \dp/n408 , \dp/n407 , \dp/n406 , \dp/n405 ,
         \dp/n404 , \dp/n403 , \dp/n402 , \dp/n334 , \dp/n333 , \dp/n332 ,
         \dp/n331 , \dp/n330 , \dp/n329 , \dp/n328 , \dp/n327 , \dp/n326 ,
         \dp/n325 , \dp/n324 , \dp/n323 , \dp/n322 , \dp/n321 , \dp/n320 ,
         \dp/n319 , \dp/n318 , \dp/n317 , \dp/n316 , \dp/n315 , \dp/n314 ,
         \dp/n313 , \dp/n312 , \dp/n311 , \dp/n310 , \dp/n309 , \dp/n308 ,
         \dp/n307 , \dp/n306 , \dp/n305 , \dp/n304 , \dp/n303 , \dp/n300 ,
         \dp/n299 , \dp/n297 , \dp/n296 , \dp/n295 , \dp/n294 , \dp/n293 ,
         \dp/n292 , \dp/n291 , \dp/n290 , \dp/n289 , \dp/n288 , \dp/n287 ,
         \dp/n286 , \dp/n285 , \dp/n284 , \dp/n283 , \dp/n282 , \dp/n281 ,
         \dp/n280 , \dp/n279 , \dp/n278 , \dp/n277 , \dp/n276 , \dp/n275 ,
         \dp/n274 , \dp/n273 , \dp/n272 , \dp/n271 , \dp/n270 , \dp/n269 ,
         \dp/n268 , \dp/n267 , \dp/n266 , \dp/n265 , \dp/n264 , \dp/n263 ,
         \dp/n262 , \dp/n261 , \dp/n260 , \dp/n259 , \dp/n258 , \dp/n257 ,
         \dp/n256 , \dp/n255 , \dp/n254 , \dp/n253 , \dp/n252 , \dp/n251 ,
         \dp/n250 , \dp/n249 , \dp/n248 , \dp/n247 , \dp/n246 , \dp/n245 ,
         \dp/n244 , \dp/n243 , \dp/n242 , \dp/n241 , \dp/n240 , \dp/n239 ,
         \dp/n238 , \dp/n237 , \dp/n236 , \dp/n235 , \dp/n234 , \dp/n233 ,
         \dp/n232 , \dp/n231 , \dp/n230 , \dp/n229 , \dp/n228 , \dp/n227 ,
         \dp/n226 , \dp/n225 , \dp/n224 , \dp/n223 , \dp/n222 , \dp/n221 ,
         \dp/n220 , \dp/n219 , \dp/n218 , \dp/n217 , \dp/n216 , \dp/n215 ,
         \dp/n214 , \dp/n213 , \dp/n212 , \dp/n211 , \dp/n210 , \dp/n209 ,
         \dp/n208 , \dp/n207 , \dp/n206 , \dp/n205 , \dp/n204 , \dp/n203 ,
         \dp/n202 , \dp/n201 , \dp/n200 , \dp/n199 , \dp/n198 , \dp/n197 ,
         \dp/n196 , \dp/n195 , \dp/n194 , \dp/n193 , \dp/n192 , \dp/n191 ,
         \dp/n190 , \dp/n189 , \dp/n188 , \dp/n187 , \dp/n186 , \dp/n185 ,
         \dp/n184 , \dp/n183 , \dp/n182 , \dp/n181 , \dp/n180 , \dp/n179 ,
         \dp/n178 , \dp/n177 , \dp/n176 , \dp/n175 , \dp/n174 , \dp/n173 ,
         \dp/n172 , \dp/n171 , \dp/n170 , \dp/n169 , \dp/n168 , \dp/n167 ,
         \dp/n166 , \dp/n165 , \dp/n164 , \dp/n163 , \dp/n162 , \dp/n161 ,
         \dp/n160 , \dp/n159 , \dp/n158 , \dp/n157 , \dp/n156 , \dp/n155 ,
         \dp/n154 , \dp/n153 , \dp/n152 , \dp/n151 , \dp/n150 , \dp/n149 ,
         \dp/n148 , \dp/n147 , \dp/n146 , \dp/n145 , \dp/n144 , \dp/n143 ,
         \dp/n142 , \dp/n141 , \dp/n140 , \dp/n139 , \dp/n138 , \dp/n137 ,
         \dp/n136 , \dp/n135 , \dp/n134 , \dp/n133 , \dp/n130 , \dp/n129 ,
         \dp/n128 , \dp/n127 , \dp/n126 , \dp/n125 , \dp/n124 , \dp/n123 ,
         \dp/n122 , \dp/n121 , \dp/n120 , \dp/n119 , \dp/n118 , \dp/n117 ,
         \dp/n116 , \dp/n115 , \dp/n114 , \dp/n113 , \dp/n112 , \dp/n111 ,
         \dp/n110 , \dp/n109 , \dp/n108 , \dp/n107 , \dp/n106 , \dp/n105 ,
         \dp/n104 , \dp/n103 , \dp/n102 , \dp/n101 , \dp/n100 , \dp/n99 ,
         \dp/n98 , \dp/n97 , \dp/n96 , \dp/n95 , \dp/n94 , \dp/n93 , \dp/n92 ,
         \dp/n91 , \dp/n90 , \dp/n89 , \dp/n88 , \dp/n87 , \dp/n86 , \dp/n85 ,
         \dp/n84 , \dp/n83 , \dp/n82 , \dp/n81 , \dp/n80 , \dp/n79 , \dp/n78 ,
         \dp/n77 , \dp/n76 , \dp/n75 , \dp/n74 , \dp/n73 , \dp/n72 , \dp/n71 ,
         \dp/n70 , \dp/n67 , \dp/n66 , \dp/n65 , \dp/n64 , \dp/n63 , \dp/n62 ,
         \dp/n61 , \dp/n60 , \dp/n59 , \dp/n58 , \dp/n57 , \dp/n56 , \dp/n55 ,
         \dp/n54 , \dp/n53 , \dp/n52 , \dp/n51 , \dp/n50 , \dp/n49 , \dp/n48 ,
         \dp/n47 , \dp/n46 , \dp/n45 , \dp/n44 , \dp/n43 , \dp/n42 , \dp/n41 ,
         \dp/n40 , \dp/n39 , \dp/n38 , \dp/n37 , \dp/n36 , \dp/n35 , \dp/n34 ,
         \dp/n33 , \dp/n32 , \dp/n31 , \dp/n30 , \dp/n29 , \dp/n28 , \dp/n27 ,
         \dp/n26 , \dp/n25 , \dp/n24 , \dp/n23 , \dp/n22 , \dp/n21 , \dp/n20 ,
         \dp/n19 , \dp/n18 , \dp/n17 , \dp/n16 , \dp/n15 , \dp/n14 , \dp/n13 ,
         \dp/n12 , \dp/n11 , \dp/n10 , \dp/n9 , \dp/n8 , \dp/n7 , \dp/n6 ,
         \dp/n5 , \dp/n4 , \dp/n3 , \dp/n1015 , \dp/n1014 , \dp/n1013 ,
         \dp/n1012 , \dp/n1011 , \dp/n1010 , \dp/n1009 , \dp/n1008 ,
         \dp/n1007 , \dp/n1006 , \dp/n1005 , \dp/n1004 , \dp/n1003 ,
         \dp/n1002 , \dp/n1001 , \dp/n1000 , \dp/n999 , \dp/n998 , \dp/n997 ,
         \dp/n996 , \dp/n995 , \dp/n994 , \dp/n993 , \dp/n992 , \dp/n991 ,
         \dp/n990 , \dp/n989 , \dp/n988 , \dp/n987 , \dp/n986 , \dp/n985 ,
         \dp/n984 , \dp/n983 , \dp/n982 , \dp/n981 , \dp/n980 , \dp/n979 ,
         \dp/n978 , \dp/n977 , \dp/n976 , \dp/n975 , \dp/n974 , \dp/n973 ,
         \dp/n972 , \dp/n971 , \dp/n970 , \dp/n969 , \dp/n968 , \dp/n967 ,
         \dp/n966 , \dp/n965 , \dp/n964 , \dp/n963 , \dp/n962 , \dp/n961 ,
         \dp/n960 , \dp/n959 , \dp/n958 , \dp/n957 , \dp/n956 , \dp/n955 ,
         \dp/n954 , \dp/n953 , \dp/n952 , \dp/n951 , \dp/n950 , \dp/n949 ,
         \dp/n948 , \dp/n947 , \dp/n946 , \dp/n945 , \dp/n944 , \dp/n943 ,
         \dp/n942 , \dp/n941 , \dp/n940 , \dp/n939 , \dp/n938 , \dp/n937 ,
         \dp/n936 , \dp/n935 , \dp/n934 , \dp/n933 , \dp/n932 , \dp/n931 ,
         \dp/n930 , \dp/n929 , \dp/n928 , \dp/n927 , \dp/n926 , \dp/n925 ,
         \dp/n924 , \dp/n923 , \dp/n922 , \dp/n921 , \dp/n920 , \dp/n919 ,
         \dp/n918 , \dp/n917 , \dp/n916 , \dp/n915 , \dp/n914 , \dp/n913 ,
         \dp/n912 , \dp/n911 , \dp/n910 , \dp/n909 , \dp/n908 , \dp/n907 ,
         \dp/n906 , \dp/n905 , \dp/n904 , \dp/n903 , \dp/n902 , \dp/n901 ,
         \dp/n900 , \dp/n899 , \dp/n898 , \dp/n897 , \dp/n896 , \dp/n895 ,
         \dp/n894 , \dp/n893 , \dp/n892 , \dp/n891 , \dp/n890 , \dp/n889 ,
         \dp/n888 , \dp/n887 , \dp/n886 , \dp/n885 , \dp/n884 , \dp/n883 ,
         \dp/n882 , \dp/n881 , \dp/n880 , \dp/n879 , \dp/n878 , \dp/n877 ,
         \dp/n876 , \dp/n875 , \dp/n874 , \dp/n873 , \dp/n872 , \dp/n871 ,
         \dp/n870 , \dp/n869 , \dp/n868 , \dp/n867 , \dp/n866 , \dp/n865 ,
         \dp/n864 , \dp/n863 , \dp/n862 , \dp/n861 , \dp/n860 , \dp/n859 ,
         \dp/n858 , \dp/n857 , \dp/n856 , \dp/n855 , \dp/n854 , \dp/n853 ,
         \dp/n852 , \dp/n851 , \dp/n850 , \dp/n849 , \dp/n848 , \dp/n847 ,
         \dp/n846 , \dp/n845 , \dp/n844 , \dp/n843 , \dp/n842 , \dp/n841 ,
         \dp/n840 , \dp/n839 , \dp/n838 , \dp/n837 , \dp/n836 , \dp/n835 ,
         \dp/n834 , \dp/n833 , \dp/n832 , \dp/n831 , \dp/n830 , \dp/n829 ,
         \dp/n828 , \dp/n827 , \dp/n826 , \dp/n825 , \dp/n824 , \dp/n823 ,
         \dp/n822 , \dp/n821 , \dp/n820 , \dp/n819 , \dp/n818 , \dp/n817 ,
         \dp/n816 , \dp/n815 , \dp/n814 , \dp/n813 , \dp/n812 , \dp/n811 ,
         \dp/n810 , \dp/n809 , \dp/n808 , \dp/n807 , \dp/n806 , \dp/n805 ,
         \dp/n804 , \dp/n803 , \dp/n802 , \dp/n801 , \dp/n800 , \dp/n799 ,
         \dp/n798 , \dp/n797 , \dp/n796 , \dp/n795 , \dp/n794 , \dp/n793 ,
         \dp/n792 , \dp/n791 , \dp/n790 , \dp/n789 , \dp/n788 , \dp/n787 ,
         \dp/n786 , \dp/n785 , \dp/n784 , \dp/n783 , \dp/n782 , \dp/n781 ,
         \dp/n780 , \dp/n779 , \dp/n778 , \dp/n777 , \dp/n776 , \dp/n775 ,
         \dp/n774 , \dp/n773 , \dp/n772 , \dp/n771 , \dp/n770 , \dp/n769 ,
         \dp/n768 , \dp/n767 , \dp/n766 , \dp/n765 , \dp/n764 , \dp/n763 ,
         \dp/n762 , \dp/n761 , \dp/n760 , \dp/n759 , \dp/n758 , \dp/n757 ,
         \dp/n756 , \dp/n755 , \dp/n754 , \dp/n753 , \dp/n752 , \dp/n751 ,
         \dp/n750 , \dp/n749 , \dp/n748 , \dp/n747 , \dp/n746 , \dp/n745 ,
         \dp/n744 , \dp/n743 , \dp/n742 , \dp/n741 , \dp/n740 , \dp/n739 ,
         \dp/n738 , \dp/n737 , \dp/n736 , \dp/n735 , \dp/n734 , \dp/n733 ,
         \dp/n732 , \dp/n731 , \dp/n730 , \dp/n729 , \dp/n728 , \dp/n727 ,
         \dp/n726 , \dp/n725 , \dp/n724 , \dp/n723 , \dp/n722 , \dp/n721 ,
         \dp/n720 , \dp/n719 , \dp/n718 , \dp/n717 , \dp/n716 , \dp/n715 ,
         \dp/n714 , \dp/n713 , \dp/n712 , \dp/n706 , \dp/n705 , \dp/n704 ,
         \dp/n703 , \dp/n702 , \dp/n701 , \dp/n700 , \dp/n699 , \dp/n698 ,
         \dp/n697 , \dp/n696 , \dp/n695 , \dp/n694 , \dp/n693 , \dp/n692 ,
         \dp/n691 , \dp/n690 , \dp/n689 , \dp/n688 , \dp/n687 , \dp/n686 ,
         \dp/n685 , \dp/n684 , \dp/n683 , \dp/n682 , \dp/n681 , \dp/n680 ,
         \dp/n679 , \dp/n678 , \dp/n677 , \dp/n676 , \dp/n675 , \dp/n674 ,
         \dp/n673 , \dp/n672 , \dp/n671 , \dp/n670 , \dp/n669 , \dp/n668 ,
         \dp/n667 , \dp/n666 , \dp/n665 , \dp/n664 , \dp/n663 , \dp/n662 ,
         \dp/n661 , \dp/n660 , \dp/n659 , \dp/n658 , \dp/n657 , \dp/n656 ,
         \dp/n655 , \dp/n654 , \dp/n653 , \dp/n652 , \dp/n651 , \dp/n650 ,
         \dp/n649 , \dp/n583 , \dp/n582 , \dp/n581 , \dp/n580 , \dp/n579 ,
         \dp/n578 , \dp/n577 , \dp/n576 , \dp/n575 , \dp/n574 , \dp/n573 ,
         \dp/n572 , \dp/n571 , \dp/n570 , \dp/n569 , \dp/n568 , \dp/n567 ,
         \dp/n566 , \dp/n565 , \dp/n564 , \dp/n563 , \dp/n562 , \dp/n561 ,
         \dp/n560 , \dp/n559 , \dp/n558 , \dp/n557 , \dp/n556 , \dp/n555 ,
         \dp/n554 , \dp/n553 , \dp/n552 , \dp/n551 , \dp/n550 , \dp/n549 ,
         \dp/n548 , \dp/n547 , \dp/n546 , \dp/n545 , \dp/n544 , \dp/n543 ,
         \dp/n542 , \dp/n541 , \dp/n540 , \dp/n539 , \dp/n538 , \dp/n537 ,
         \dp/n536 , \dp/n535 , \dp/n534 , \dp/n533 , \dp/n532 , \dp/n531 ,
         \dp/n530 , \dp/n529 , \dp/n528 , \dp/n527 , \dp/n526 , \dp/n524 ,
         \dp/n522 , \dp/n520 , \dp/n518 , \dp/n516 , \dp/n515 , \dp/n514 ,
         \dp/n513 , \dp/n512 , \dp/n511 , \dp/n510 , \dp/n509 , \dp/n508 ,
         \dp/n507 , \dp/n506 , \dp/n505 , \dp/n504 , \dp/n503 , \dp/n502 ,
         \dp/n501 , \dp/n500 , \dp/n499 , \dp/n498 , \dp/n497 , \dp/n496 ,
         \dp/n495 , \dp/n494 , \dp/n493 , \dp/n492 , \dp/n491 , \dp/n490 ,
         \dp/n489 , \dp/n488 , \dp/n487 , \dp/n486 , \dp/n485 , \dp/n484 ,
         \dp/n483 , \dp/n482 , \dp/n481 , \dp/n480 , \dp/n479 , \dp/n478 ,
         \dp/n477 , \dp/n476 , \dp/n475 , \dp/n474 , \dp/n473 , \dp/n472 ,
         \dp/n471 , \dp/n470 , \dp/n469 , \dp/n468 , \dp/n467 , \dp/n466 ,
         \dp/n465 , \dp/n464 , \dp/n463 , \dp/n462 , \dp/n461 , \dp/n460 ,
         \dp/n459 , \dp/n458 , \dp/n457 , \dp/n456 , \dp/n455 , \dp/n454 ,
         \dp/n453 , \dp/n452 , \dp/n451 , \dp/n450 , \dp/n449 , \dp/n448 ,
         \dp/n447 , \dp/n446 , \dp/n445 , \dp/n444 , \dp/n443 , \dp/n442 ,
         \dp/n441 , \dp/n440 , \dp/n439 , \dp/n438 , \dp/n437 , \dp/n436 ,
         \dp/n435 , \dp/n434 , \dp/n433 , \dp/n432 , \dp/n431 , \dp/n430 ,
         \dp/n429 , \dp/n428 , \dp/n427 , \dp/n426 , \dp/n425 , \dp/n424 ,
         \dp/n423 , \dp/n422 , \dp/n421 , \dp/n420 , \dp/n419 , \dp/n418 ,
         \dp/n417 , \dp/n416 , \dp/n415 , \dp/n414 , \dp/n401 , \dp/n400 ,
         \dp/n399 , \dp/n398 , \dp/n397 , \dp/n396 , \dp/n395 , \dp/n394 ,
         \dp/n393 , \dp/n392 , \dp/n391 , \dp/n390 , \dp/n389 , \dp/n388 ,
         \dp/n387 , \dp/n386 , \dp/n385 , \dp/n384 , \dp/n383 , \dp/n382 ,
         \dp/n381 , \dp/n380 , \dp/n379 , \dp/n378 , \dp/n377 , \dp/n376 ,
         \dp/n375 , \dp/n374 , \dp/n373 , \dp/n372 , \dp/n371 , \dp/n370 ,
         \dp/n369 , \dp/n368 , \dp/n367 , \dp/n366 , \dp/n365 , \dp/n364 ,
         \dp/n363 , \dp/n362 , \dp/n361 , \dp/n360 , \dp/n359 , \dp/n358 ,
         \dp/n357 , \dp/n356 , \dp/n355 , \dp/n354 , \dp/n353 , \dp/n352 ,
         \dp/n351 , \dp/n350 , \dp/n349 , \dp/n348 , \dp/n347 , \dp/n346 ,
         \dp/n345 , \dp/n344 , \dp/n343 , \dp/n342 , \dp/n341 , \dp/n340 ,
         \dp/n339 , \dp/n338 , \dp/n337 , \dp/n336 , \dp/n335 , \dp/n302 ,
         \dp/n301 , \dp/n298 , \dp/n132 , \dp/n131 , \dp/n69 , \dp/n68 ,
         \dp/branch_t_ex_o , \dp/ir[0] , \dp/ir[1] , \dp/ir[2] , \dp/ir[3] ,
         \dp/ir[4] , \dp/ir[5] , \dp/ir[6] , \dp/ir[7] , \dp/ir[8] ,
         \dp/ir[9] , \dp/ir[10] , \dp/ir[11] , \dp/ir[12] , \dp/ir[13] ,
         \dp/ir[14] , \dp/ir[15] , \dp/ir[16] , \dp/ir[17] , \dp/ir[18] ,
         \dp/ir[19] , \dp/ir[20] , \dp/ir[21] , \dp/ir[22] , \dp/ir[23] ,
         \dp/ir[24] , \dp/ir[25] , \dp/if_stage/n104 , \dp/if_stage/n103 ,
         \dp/if_stage/n102 , \dp/if_stage/n101 , \dp/if_stage/n100 ,
         \dp/if_stage/n99 , \dp/if_stage/n96 , \dp/if_stage/n97 ,
         \dp/if_stage/n95 , \dp/if_stage/n94 , \dp/if_stage/n93 ,
         \dp/if_stage/n92 , \dp/if_stage/n91 , \dp/if_stage/n90 ,
         \dp/if_stage/n89 , \dp/if_stage/n88 , \dp/if_stage/n87 ,
         \dp/if_stage/n86 , \dp/if_stage/n85 , \dp/if_stage/n84 ,
         \dp/if_stage/n83 , \dp/if_stage/n82 , \dp/if_stage/n81 ,
         \dp/if_stage/n80 , \dp/if_stage/n79 , \dp/if_stage/n78 ,
         \dp/if_stage/n77 , \dp/if_stage/n76 , \dp/if_stage/n75 ,
         \dp/if_stage/n74 , \dp/if_stage/n73 , \dp/if_stage/n72 ,
         \dp/if_stage/n71 , \dp/if_stage/n70 , \dp/if_stage/n69 ,
         \dp/if_stage/n68 , \dp/if_stage/n67 , \dp/if_stage/n66 ,
         \dp/if_stage/n65 , \dp/if_stage/n64 , \dp/if_stage/n63 ,
         \dp/if_stage/n62 , \dp/if_stage/n61 , \dp/if_stage/n60 ,
         \dp/if_stage/n59 , \dp/if_stage/n58 , \dp/if_stage/n57 ,
         \dp/if_stage/n56 , \dp/if_stage/n55 , \dp/if_stage/n54 ,
         \dp/if_stage/n53 , \dp/if_stage/n52 , \dp/if_stage/n51 ,
         \dp/if_stage/n50 , \dp/if_stage/n49 , \dp/if_stage/n48 ,
         \dp/if_stage/n47 , \dp/if_stage/n46 , \dp/if_stage/n45 ,
         \dp/if_stage/n44 , \dp/if_stage/n43 , \dp/if_stage/n42 ,
         \dp/if_stage/n41 , \dp/if_stage/n40 , \dp/if_stage/n39 ,
         \dp/if_stage/n38 , \dp/if_stage/n37 , \dp/if_stage/n36 ,
         \dp/if_stage/n35 , \dp/if_stage/n34 , \dp/if_stage/n33 ,
         \dp/if_stage/n32 , \dp/if_stage/n31 , \dp/if_stage/n30 ,
         \dp/if_stage/n29 , \dp/if_stage/n28 , \dp/if_stage/n27 ,
         \dp/if_stage/n26 , \dp/if_stage/n25 , \dp/if_stage/n24 ,
         \dp/if_stage/n23 , \dp/if_stage/n22 , \dp/if_stage/n21 ,
         \dp/if_stage/n20 , \dp/if_stage/n19 , \dp/if_stage/n18 ,
         \dp/if_stage/n17 , \dp/if_stage/n16 , \dp/if_stage/n15 ,
         \dp/if_stage/n14 , \dp/if_stage/n13 , \dp/if_stage/n12 ,
         \dp/if_stage/n11 , \dp/if_stage/n10 , \dp/if_stage/n9 ,
         \dp/if_stage/n8 , \dp/if_stage/n7 , \dp/if_stage/n6 ,
         \dp/if_stage/n5 , \dp/if_stage/n4 , \dp/if_stage/n3 ,
         \dp/if_stage/n2 , \dp/if_stage/n1 , \dp/if_stage/mux/n14 ,
         \dp/if_stage/mux/n13 , \dp/if_stage/mux/n12 , \dp/if_stage/mux/n11 ,
         \dp/if_stage/mux/n10 , \dp/if_stage/mux/n9 , \dp/if_stage/mux/n8 ,
         \dp/if_stage/mux/n7 , \dp/if_stage/mux/n6 , \dp/if_stage/mux/n5 ,
         \dp/if_stage/mux/n4 , \dp/if_stage/mux/n3 , \dp/if_stage/mux/n2 ,
         \dp/if_stage/mux/n1 , \dp/if_stage/mux/n65 , \dp/if_stage/mux/n64 ,
         \dp/if_stage/mux/n63 , \dp/if_stage/mux/n62 , \dp/if_stage/mux/n61 ,
         \dp/if_stage/mux/n60 , \dp/if_stage/mux/n59 , \dp/if_stage/mux/n58 ,
         \dp/if_stage/mux/n57 , \dp/if_stage/mux/n56 , \dp/if_stage/mux/n55 ,
         \dp/if_stage/mux/n54 , \dp/if_stage/mux/n53 , \dp/if_stage/mux/n52 ,
         \dp/if_stage/mux/n51 , \dp/if_stage/mux/n50 , \dp/if_stage/mux/n49 ,
         \dp/if_stage/mux/n48 , \dp/if_stage/mux/n47 , \dp/if_stage/mux/n46 ,
         \dp/if_stage/mux/n45 , \dp/if_stage/mux/n44 , \dp/if_stage/mux/n43 ,
         \dp/if_stage/mux/n42 , \dp/if_stage/mux/n41 , \dp/if_stage/mux/n40 ,
         \dp/if_stage/mux/n39 , \dp/if_stage/mux/n38 , \dp/if_stage/mux/n37 ,
         \dp/if_stage/mux/n36 , \dp/if_stage/mux/n35 , \dp/if_stage/mux/n34 ,
         \dp/if_stage/add_77/n57 , \dp/if_stage/add_77/n56 ,
         \dp/if_stage/add_77/n55 , \dp/if_stage/add_77/n54 ,
         \dp/if_stage/add_77/n53 , \dp/if_stage/add_77/n52 ,
         \dp/if_stage/add_77/n51 , \dp/if_stage/add_77/n50 ,
         \dp/if_stage/add_77/n49 , \dp/if_stage/add_77/n48 ,
         \dp/if_stage/add_77/n47 , \dp/if_stage/add_77/n46 ,
         \dp/if_stage/add_77/n45 , \dp/if_stage/add_77/n44 ,
         \dp/if_stage/add_77/n43 , \dp/if_stage/add_77/n42 ,
         \dp/if_stage/add_77/n41 , \dp/if_stage/add_77/n40 ,
         \dp/if_stage/add_77/n39 , \dp/if_stage/add_77/n38 ,
         \dp/if_stage/add_77/n37 , \dp/if_stage/add_77/n36 ,
         \dp/if_stage/add_77/n35 , \dp/if_stage/add_77/n34 ,
         \dp/if_stage/add_77/n33 , \dp/if_stage/add_77/n32 ,
         \dp/if_stage/add_77/n31 , \dp/if_stage/add_77/n30 , \dp/id_stage/n40 ,
         \dp/id_stage/n39 , \dp/id_stage/n38 , \dp/id_stage/n37 ,
         \dp/id_stage/n36 , \dp/id_stage/n35 , \dp/id_stage/n34 ,
         \dp/id_stage/n33 , \dp/id_stage/n32 , \dp/id_stage/n31 ,
         \dp/id_stage/n30 , \dp/id_stage/n29 , \dp/id_stage/n28 ,
         \dp/id_stage/n27 , \dp/id_stage/n26 , \dp/id_stage/n25 ,
         \dp/id_stage/n24 , \dp/id_stage/n16 , \dp/id_stage/n15 ,
         \dp/id_stage/n14 , \dp/id_stage/n13 , \dp/id_stage/n12 ,
         \dp/id_stage/n11 , \dp/id_stage/n10 , \dp/id_stage/n9 ,
         \dp/id_stage/n8 , \dp/id_stage/n7 , \dp/id_stage/n6 ,
         \dp/id_stage/n5 , \dp/id_stage/n4 , \dp/id_stage/n3 ,
         \dp/id_stage/n2 , \dp/id_stage/n1 , \dp/id_stage/n23 ,
         \dp/id_stage/n22 , \dp/id_stage/n21 , \dp/id_stage/n20 ,
         \dp/id_stage/n19 , \dp/id_stage/n18 , \dp/id_stage/n17 ,
         \dp/id_stage/regfile/cpu_work , \dp/id_stage/regfile/sel_wp ,
         \dp/id_stage/regfile/end_sf , \dp/id_stage/regfile/canrestore ,
         \dp/id_stage/regfile/cansave , \dp/id_stage/regfile/up_dwn_rest ,
         \dp/id_stage/regfile/up_dwn_save , \dp/id_stage/regfile/up_dwn_cwp ,
         \dp/id_stage/regfile/up_dwn_swp ,
         \dp/id_stage/regfile/rst_spill_fill , \dp/id_stage/regfile/rst_swp ,
         \dp/id_stage/regfile/cnt_save , \dp/id_stage/regfile/cnt_cwp ,
         \dp/id_stage/regfile/cnt_swp , \dp/id_stage/regfile/rst_rf ,
         \dp/id_stage/regfile/rf_enable , \dp/id_stage/regfile/wr_cu ,
         \dp/id_stage/regfile/rd_cu , \dp/id_stage/regfile/ControlUnit/n15 ,
         \dp/id_stage/regfile/ControlUnit/n11 ,
         \dp/id_stage/regfile/ControlUnit/n9 ,
         \dp/id_stage/regfile/ControlUnit/n8 ,
         \dp/id_stage/regfile/ControlUnit/n5 ,
         \dp/id_stage/regfile/ControlUnit/n4 ,
         \dp/id_stage/regfile/ControlUnit/n3 ,
         \dp/id_stage/regfile/ControlUnit/n2 ,
         \dp/id_stage/regfile/ControlUnit/n40 ,
         \dp/id_stage/regfile/ControlUnit/n39 ,
         \dp/id_stage/regfile/ControlUnit/n38 ,
         \dp/id_stage/regfile/ControlUnit/n37 ,
         \dp/id_stage/regfile/ControlUnit/n36 ,
         \dp/id_stage/regfile/ControlUnit/n35 ,
         \dp/id_stage/regfile/ControlUnit/n34 ,
         \dp/id_stage/regfile/ControlUnit/n33 ,
         \dp/id_stage/regfile/ControlUnit/n32 ,
         \dp/id_stage/regfile/ControlUnit/n31 ,
         \dp/id_stage/regfile/ControlUnit/n30 ,
         \dp/id_stage/regfile/ControlUnit/n29 ,
         \dp/id_stage/regfile/ControlUnit/n28 ,
         \dp/id_stage/regfile/ControlUnit/n27 ,
         \dp/id_stage/regfile/ControlUnit/n26 ,
         \dp/id_stage/regfile/ControlUnit/n25 ,
         \dp/id_stage/regfile/ControlUnit/n24 ,
         \dp/id_stage/regfile/ControlUnit/n23 ,
         \dp/id_stage/regfile/ControlUnit/n22 ,
         \dp/id_stage/regfile/ControlUnit/n21 ,
         \dp/id_stage/regfile/ControlUnit/n20 ,
         \dp/id_stage/regfile/ControlUnit/n19 ,
         \dp/id_stage/regfile/ControlUnit/n18 ,
         \dp/id_stage/regfile/ControlUnit/n17 ,
         \dp/id_stage/regfile/ControlUnit/n16 ,
         \dp/id_stage/regfile/ControlUnit/n14 ,
         \dp/id_stage/regfile/ControlUnit/n13 ,
         \dp/id_stage/regfile/ControlUnit/n12 ,
         \dp/id_stage/regfile/ControlUnit/current_state[0] ,
         \dp/id_stage/regfile/ControlUnit/current_state[1] ,
         \dp/id_stage/regfile/ControlUnit/current_state[2] ,
         \dp/id_stage/regfile/ControlUnit/current_state[3] ,
         \dp/id_stage/regfile/DataPath/mux_en_control_out ,
         \dp/id_stage/regfile/DataPath/mux_wr_control_out ,
         \dp/id_stage/regfile/DataPath/mux_rd2_control_out ,
         \dp/id_stage/regfile/DataPath/mux_rd1_control_out ,
         \dp/id_stage/regfile/DataPath/cwp_1[0] ,
         \dp/id_stage/regfile/DataPath/spill_fill_addr[0] ,
         \dp/id_stage/regfile/DataPath/spill_fill_addr[1] ,
         \dp/id_stage/regfile/DataPath/spill_fill_addr[2] ,
         \dp/id_stage/regfile/DataPath/spill_fill_addr[3] ,
         \dp/id_stage/regfile/DataPath/spill_fill_addr[4] ,
         \dp/id_stage/regfile/DataPath/spill_fill_addr[5] ,
         \dp/id_stage/regfile/DataPath/sf_wp[0] ,
         \dp/id_stage/regfile/DataPath/addr_sf_in[0] ,
         \dp/id_stage/regfile/DataPath/addr_sf_in[1] ,
         \dp/id_stage/regfile/DataPath/addr_sf_in[2] ,
         \dp/id_stage/regfile/DataPath/CWP[0] ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n4 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n3 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n2 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n1 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n22 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n21 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n20 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n19 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/n18 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/N5 ,
         \dp/id_stage/regfile/DataPath/Conv_RD1/N1 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n13 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n12 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n11 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n10 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n9 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n4 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n3 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n2 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/n1 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/N5 ,
         \dp/id_stage/regfile/DataPath/Conv_RD2/N1 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n13 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n12 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n11 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n10 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n9 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n8 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n4 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n3 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n2 ,
         \dp/id_stage/regfile/DataPath/Conv_W/n1 ,
         \dp/id_stage/regfile/DataPath/Conv_W/N5 ,
         \dp/id_stage/regfile/DataPath/Conv_W/N1 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n10 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n9 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n8 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n7 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n6 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n5 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n4 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n3 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n2 ,
         \dp/id_stage/regfile/DataPath/SF_converter/n1 ,
         \dp/id_stage/regfile/DataPath/SF_converter/N5 ,
         \dp/id_stage/regfile/DataPath/SF_converter/N1 ,
         \dp/id_stage/regfile/DataPath/Cwp_counter/n4 ,
         \dp/id_stage/regfile/DataPath/Cwp_counter/n2 ,
         \dp/id_stage/regfile/DataPath/Cwp_counter/n5 ,
         \dp/id_stage/regfile/DataPath/Cwp_counter/n3 ,
         \dp/id_stage/regfile/DataPath/Cwp_counter/n1 ,
         \dp/id_stage/regfile/DataPath/Swp_counter/n8 ,
         \dp/id_stage/regfile/DataPath/Swp_counter/n7 ,
         \dp/id_stage/regfile/DataPath/Swp_counter/n6 ,
         \dp/id_stage/regfile/DataPath/Swp_counter/n4 ,
         \dp/id_stage/regfile/DataPath/Swp_counter/n2 ,
         \dp/id_stage/regfile/DataPath/Swp_counter/Q[0] ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n16 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n12 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n4 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n3 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n2 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n1 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n21 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n20 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n19 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n18 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n17 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n15 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n14 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n13 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n11 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n10 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n9 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n8 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n7 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n6 ,
         \dp/id_stage/regfile/DataPath/Spill_fill_counter/n5 ,
         \dp/id_stage/regfile/DataPath/CANSAVE_counter/n8 ,
         \dp/id_stage/regfile/DataPath/CANSAVE_counter/n7 ,
         \dp/id_stage/regfile/DataPath/CANSAVE_counter/n6 ,
         \dp/id_stage/regfile/DataPath/CANSAVE_counter/n4 ,
         \dp/id_stage/regfile/DataPath/CANSAVE_counter/n2 ,
         \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n8 ,
         \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n7 ,
         \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n6 ,
         \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n4 ,
         \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n2 ,
         \dp/id_stage/regfile/DataPath/Mux_rd/n1 ,
         \dp/id_stage/regfile/DataPath/Mux_rd/n13 ,
         \dp/id_stage/regfile/DataPath/Mux_rd/n12 ,
         \dp/id_stage/regfile/DataPath/Mux_rd/n11 ,
         \dp/id_stage/regfile/DataPath/Mux_rd/n10 ,
         \dp/id_stage/regfile/DataPath/Mux_rd/n9 ,
         \dp/id_stage/regfile/DataPath/Mux_rd/n8 ,
         \dp/id_stage/regfile/DataPath/Mux_wr/n7 ,
         \dp/id_stage/regfile/DataPath/Mux_wr/n6 ,
         \dp/id_stage/regfile/DataPath/Mux_wr/n5 ,
         \dp/id_stage/regfile/DataPath/Mux_wr/n4 ,
         \dp/id_stage/regfile/DataPath/Mux_wr/n3 ,
         \dp/id_stage/regfile/DataPath/Mux_wr/n2 ,
         \dp/id_stage/regfile/DataPath/Mux_wr/n1 ,
         \dp/id_stage/regfile/DataPath/Mux_sf/n1 ,
         \dp/id_stage/regfile/DataPath/Mux_sf/n3 ,
         \dp/id_stage/regfile/DataPath/Mux_rd1_control/n2 ,
         \dp/id_stage/regfile/DataPath/Mux_rd1_control/n3 ,
         \dp/id_stage/regfile/DataPath/Mux_rd2_control/n4 ,
         \dp/id_stage/regfile/DataPath/Mux_rd2_control/n2 ,
         \dp/id_stage/regfile/DataPath/Mux_wr_control/n4 ,
         \dp/id_stage/regfile/DataPath/Mux_wr_control/n2 ,
         \dp/id_stage/regfile/DataPath/Mux_en_control/n4 ,
         \dp/id_stage/regfile/DataPath/Mux_en_control/n2 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4276 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4242 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4241 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4240 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4239 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4235 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4231 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4230 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4229 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4228 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4227 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4226 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4225 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4222 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4221 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4220 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4219 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4218 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4217 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4216 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4213 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4212 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4211 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4210 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4209 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4208 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4207 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4204 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4203 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4202 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4201 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4200 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4199 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4198 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4195 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4194 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4193 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4192 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4191 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4190 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4189 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4186 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4185 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4184 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4183 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4182 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4181 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4180 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4177 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4176 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4175 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4174 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4173 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4172 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4171 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4168 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4167 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4166 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4165 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4164 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4163 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4162 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4159 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4158 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4157 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4156 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4155 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4154 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4153 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4150 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4149 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4148 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4147 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4146 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4145 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4144 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4141 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4140 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4139 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4138 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4137 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4136 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4135 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4132 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4131 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4130 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4129 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4128 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4127 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4126 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4123 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4122 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4121 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4120 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4119 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4118 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4117 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4114 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4113 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4112 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4111 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4110 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4109 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4108 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4105 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4104 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4103 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4102 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4101 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4100 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4099 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4096 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4095 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4094 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4093 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4092 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4091 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4090 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4087 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4086 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4085 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4084 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4083 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4082 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4081 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4078 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4077 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4076 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4075 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4074 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4073 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4072 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4069 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4068 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4067 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4066 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4065 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4064 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4063 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4060 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4059 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4058 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4057 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4056 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4055 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4054 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4051 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4050 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4049 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4048 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4047 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4046 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4045 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4042 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4041 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4040 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4039 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4038 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4037 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4036 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4033 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4032 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4031 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4030 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4029 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4028 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4027 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4024 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4023 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4022 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4021 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4020 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4019 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4018 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4015 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4014 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4013 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4012 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4011 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4010 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4009 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4006 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4005 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4004 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4003 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4002 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4001 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4000 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3997 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3996 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3995 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3994 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3993 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3992 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3991 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3988 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3987 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3986 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3985 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3984 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3983 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3982 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3979 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3978 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3977 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3976 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3975 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3974 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3973 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3970 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3969 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3968 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3967 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3966 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3965 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3964 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3961 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3960 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3959 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3958 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3957 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3956 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3955 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3952 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3951 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3950 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3949 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3948 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3947 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3946 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3943 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3942 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3941 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3940 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3939 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3938 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3937 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3934 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3933 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3932 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3931 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3930 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3929 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3928 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3925 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3924 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3923 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3922 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3921 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3920 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3919 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3916 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3915 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3914 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3913 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3912 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3911 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3910 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1925 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1858 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1857 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1756 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1755 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1688 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1687 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1586 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1585 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1518 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1516 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1348 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1346 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1226 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1220 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1213 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1207 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1189 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1177 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1176 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1175 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1174 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1173 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1172 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1171 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1170 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1169 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3692 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3691 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3690 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3689 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3688 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3687 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3686 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3685 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3684 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3683 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3682 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3681 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3680 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3679 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3678 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3677 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3676 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3675 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3674 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3673 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3672 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3671 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3670 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3669 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3668 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3667 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3666 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3665 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3664 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3663 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3662 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3661 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3660 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3659 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3658 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3657 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3656 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3655 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3654 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3653 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3652 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3651 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3650 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3649 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3648 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3647 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3646 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3645 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3644 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3643 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3642 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3641 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3640 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3639 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3638 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3637 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3636 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3635 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3634 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3633 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3632 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3631 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3630 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3629 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3628 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3627 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3626 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3625 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3624 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3623 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3622 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3621 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3620 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3619 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3618 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3617 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3616 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3615 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3614 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3613 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3612 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3611 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3610 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3609 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3608 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3607 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3606 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3605 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3604 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3603 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3602 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3601 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3600 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3599 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3598 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3597 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3596 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3595 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3594 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3593 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3592 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3591 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3590 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3589 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3588 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3587 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3586 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3585 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3584 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3583 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3582 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3581 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3580 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3579 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3578 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3577 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3576 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3575 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3574 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3573 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3572 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3571 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3570 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3569 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3568 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3567 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3566 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3565 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3564 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3563 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3562 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3561 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3560 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3559 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3558 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3557 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3556 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3555 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3554 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3553 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3552 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3551 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3550 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3549 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3548 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3547 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3546 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3545 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3544 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3543 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3542 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3541 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3540 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3539 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3538 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3537 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3536 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3535 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3534 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3533 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3532 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3531 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3530 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3529 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3528 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3527 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3526 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3525 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3524 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3523 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3522 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3521 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3520 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3519 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3518 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3517 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3516 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3515 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3514 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3513 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3512 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3511 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3510 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3509 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3508 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3507 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3506 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3505 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3504 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3503 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3502 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3501 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3500 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3499 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3498 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3497 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3496 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3495 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3494 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3493 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3492 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3491 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3490 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3489 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3488 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3487 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3486 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3485 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3484 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3483 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3482 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3481 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3480 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3479 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3478 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3477 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3476 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3475 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3474 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3473 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3472 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3471 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3470 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3469 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3468 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3467 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3466 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3465 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3464 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3463 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3462 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3461 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3460 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3459 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3458 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3457 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3456 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3455 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3454 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3453 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3452 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3451 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3450 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3449 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3448 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3447 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3446 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3445 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3444 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3443 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3442 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3441 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3440 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3439 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3438 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3437 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3436 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3435 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3434 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3433 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3432 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3431 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3430 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3429 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3428 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3427 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3426 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3425 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3424 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3423 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3422 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3421 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3420 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3419 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3418 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3417 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3416 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3415 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3414 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3413 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3412 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3411 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3410 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3409 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3408 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3407 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3406 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3405 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3404 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3403 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3402 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3401 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3400 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3399 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3398 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3397 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3396 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3395 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3394 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3393 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3392 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3391 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3390 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3389 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3388 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3387 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3386 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3385 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3384 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3383 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3382 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3381 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3380 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3379 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3378 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3377 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3376 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3375 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3374 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3373 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3372 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3371 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3370 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3369 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3368 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3367 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3366 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3365 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3364 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3363 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3362 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3361 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3360 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3359 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3358 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3357 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3356 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3355 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3354 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3353 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3352 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3351 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3350 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3349 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3348 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3347 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3346 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3345 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3344 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3343 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3342 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3341 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3340 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3339 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3338 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3337 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3336 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3335 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3334 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3333 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3332 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3331 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3330 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3329 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3328 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3327 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3326 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3325 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3324 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3323 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3322 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3321 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3320 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3319 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3318 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3317 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3316 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3315 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3314 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3313 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3312 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3311 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3310 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3309 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3308 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3307 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3306 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3305 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3304 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3303 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3302 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3301 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3300 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3299 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3298 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3297 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3296 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3295 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3294 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3293 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3292 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3291 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3290 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3289 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3288 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3287 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3286 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3285 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3284 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3283 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3282 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3281 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3280 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3279 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3278 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3277 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3276 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3275 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3274 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3273 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3272 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3271 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3270 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3269 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3268 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3267 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3266 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3265 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3264 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3263 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3262 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3261 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3260 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3259 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3258 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3257 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3256 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3255 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3254 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3253 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3252 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3251 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3250 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3249 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3248 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3247 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3246 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3245 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3244 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3243 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3242 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3241 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3240 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3239 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3238 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3237 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3236 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3235 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3234 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3233 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3232 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3231 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3230 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3229 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3228 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3227 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3226 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3225 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3224 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3223 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3222 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3221 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3220 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3219 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3218 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3217 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3216 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3215 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3214 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3213 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3212 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3211 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3210 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3209 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3208 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3207 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3206 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3205 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3204 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3203 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3202 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3201 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3200 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3199 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3198 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3197 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3196 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3195 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3194 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3193 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3192 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3191 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3190 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3189 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3188 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3187 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3186 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3185 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3184 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3183 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3182 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3181 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3180 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3179 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3178 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3177 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3176 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3175 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3174 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3173 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3172 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3171 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3170 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3169 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3168 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3167 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3166 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3165 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3164 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3163 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3162 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3161 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3158 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3155 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3154 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3153 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3152 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3151 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3150 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3149 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3148 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3147 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3146 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3145 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3144 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3143 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3142 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3141 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3140 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3139 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3138 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3137 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3136 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3135 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3134 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3133 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3132 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3131 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3130 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3129 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3128 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3127 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3126 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3125 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3124 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3123 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3122 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3121 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3120 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3119 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3118 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3117 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3116 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3115 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3114 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3113 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3112 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3111 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3110 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3109 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3108 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3107 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3106 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3105 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3104 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3103 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3102 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3101 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3100 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3099 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3098 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3097 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3096 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3095 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3094 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3093 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3092 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3091 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3090 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3089 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3088 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3087 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3086 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3085 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3084 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3083 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3082 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3081 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3080 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3079 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3078 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3077 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3076 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3075 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3074 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3073 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3072 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3071 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3070 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3069 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3068 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3067 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3066 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3065 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3064 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3063 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3062 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3061 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3060 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3059 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3058 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3057 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3056 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3055 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3054 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3053 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3052 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3051 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3050 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3049 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3048 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3047 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3046 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3045 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3044 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3043 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3042 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3041 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3040 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3039 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3038 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3037 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3036 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3035 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3034 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3033 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3032 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3031 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3030 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3029 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3028 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3027 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3026 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3025 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3024 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3023 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3022 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3021 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3020 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3019 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3018 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3017 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3016 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3015 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3014 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3013 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3012 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3011 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3010 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3009 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3008 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3007 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3006 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3005 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3004 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3003 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3002 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3001 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3000 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2999 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2998 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2997 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2996 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2995 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2994 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2993 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2992 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2991 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2990 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2989 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2988 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2987 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2986 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2985 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2984 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2983 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2982 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2981 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2980 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2979 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2978 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2977 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2976 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2975 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2974 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2973 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2972 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2971 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2970 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2969 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2968 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2967 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2966 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2965 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2964 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2963 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2962 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2961 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2960 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2959 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2958 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2957 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2956 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2955 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2954 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2953 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2952 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2951 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2950 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2949 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2948 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2947 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2946 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2945 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2944 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2943 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2942 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2941 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2940 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2939 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2938 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2937 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2936 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2935 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2934 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2933 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2932 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2931 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2930 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2929 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2928 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2927 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2926 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2925 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2924 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2923 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2922 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2921 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2920 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2919 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2918 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2917 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2916 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2915 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2914 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2913 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2912 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2911 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2910 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2909 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2908 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2907 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2906 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2905 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2904 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2903 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2902 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2901 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2900 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2899 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2898 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2897 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2896 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2895 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2894 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2893 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2892 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2891 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2890 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2889 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2888 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2887 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2886 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2885 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2884 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2883 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2882 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2881 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2880 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2879 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2878 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2877 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2876 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2875 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2874 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2873 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2872 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2871 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2870 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2869 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2868 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2867 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2866 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2865 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2864 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2863 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2862 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2861 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2860 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2859 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2858 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2857 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2856 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2855 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2854 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2853 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2852 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2851 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2850 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2849 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2848 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2847 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2846 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2845 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2844 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2843 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2842 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2841 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2840 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2839 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2838 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2837 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2836 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2835 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2834 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2833 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2832 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2831 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2830 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2829 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2828 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2827 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2826 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2825 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2824 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2823 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2822 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2821 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2820 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2819 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2818 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2817 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2816 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2815 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2814 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2813 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2812 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2811 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2810 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2809 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2808 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2807 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2806 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2805 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2804 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2803 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2802 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2801 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2800 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2799 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2798 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2797 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2796 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2795 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2794 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2793 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2792 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2791 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2790 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2789 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2788 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2787 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2786 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2785 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2784 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2783 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2782 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2781 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2780 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2779 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2778 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2777 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2776 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2775 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2774 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2773 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2772 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2771 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2770 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2769 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2768 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2767 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2766 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2765 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2764 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2763 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2762 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2761 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2760 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2759 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2758 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2757 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2756 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2755 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2754 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2753 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2752 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2751 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2750 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2749 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2748 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2747 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2746 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2745 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2744 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2743 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2742 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2741 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2740 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2739 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2738 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2737 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2736 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2735 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2734 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2733 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2732 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2731 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2730 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2729 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2728 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2727 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2726 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2725 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2724 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2723 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2722 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2721 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2720 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2719 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2718 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2717 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2716 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2715 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2714 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2713 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2712 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2711 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2710 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2709 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2708 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2707 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2706 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2705 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2704 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2703 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2702 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2701 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2700 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2699 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2698 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2697 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2696 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2695 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2694 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2693 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2692 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2691 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2690 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2689 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2688 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2687 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2686 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2685 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2684 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2683 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2682 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2681 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2680 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2679 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2678 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2677 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2676 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2675 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2674 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2673 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2672 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2671 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2670 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2669 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2668 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2667 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2666 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2665 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2664 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2663 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2662 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2661 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2660 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2659 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2658 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2657 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2656 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2655 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2654 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2653 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2652 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2651 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2650 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2649 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2648 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2647 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2646 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2645 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2644 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2643 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2642 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2641 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2640 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2639 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2638 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2637 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2636 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2635 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2634 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2633 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2632 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2631 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2630 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2629 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2628 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2627 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2626 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2625 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2624 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2623 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2622 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2621 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2620 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2619 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2618 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2617 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2616 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2615 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2614 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2613 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2612 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2611 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2610 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2609 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2608 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2607 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2606 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2605 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2604 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2603 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2602 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2601 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2600 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2599 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2598 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2597 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2596 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2595 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2594 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2593 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2592 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2591 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2590 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2589 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2588 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2587 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2586 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2585 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2584 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2583 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2582 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2581 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2580 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2579 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2578 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2577 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2576 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2575 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2574 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2573 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2572 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2571 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2570 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2569 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2568 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2567 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2566 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2565 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2564 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2563 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2562 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2561 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2560 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2559 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2558 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2557 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2556 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2555 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2554 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2553 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2552 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2551 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2550 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2549 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2548 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2547 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2546 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2545 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2544 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2543 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2542 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2541 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2540 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2539 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2538 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2537 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2536 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2535 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2534 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2531 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2528 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2527 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2526 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2525 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2524 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2523 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2522 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2521 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2520 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2519 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2518 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2517 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2516 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2515 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2514 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2513 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2512 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2511 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2510 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2509 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2508 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2507 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2506 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2505 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2504 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2503 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2502 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2501 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2500 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2499 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2498 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2497 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2496 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2495 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2494 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2493 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2492 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2491 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2490 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2489 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2488 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2487 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2486 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2485 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2484 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2483 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2482 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2481 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2480 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2479 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2478 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2477 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2476 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2475 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2474 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2473 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2472 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2471 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2470 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2469 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2468 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2467 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2466 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2465 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2464 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2463 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2462 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2461 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2460 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2459 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2458 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2457 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2456 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2455 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2454 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2453 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2452 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2451 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2450 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2449 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2448 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2447 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2446 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2445 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2444 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2443 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2442 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2441 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2440 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2439 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2438 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2437 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2436 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2435 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2434 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2433 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2432 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2431 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2430 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2429 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2428 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2427 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2426 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2425 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2424 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2423 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2422 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2421 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2420 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2419 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2418 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2417 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2416 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2415 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2414 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2413 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2412 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2411 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2410 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2409 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2408 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2407 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2406 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2405 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2404 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2403 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2402 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2401 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2400 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2399 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2398 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2397 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2396 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2395 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2394 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2393 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2392 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2391 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2390 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2389 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2388 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2387 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2386 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2385 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2384 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2383 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2382 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2381 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2380 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2379 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2378 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2377 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2376 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2375 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2374 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2373 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2372 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2371 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2370 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2369 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2368 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2367 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2366 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2365 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2364 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2363 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2362 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2361 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2360 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2359 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2358 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2357 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2356 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2355 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2354 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2353 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2352 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2351 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2350 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2349 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2348 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2347 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2346 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2345 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2344 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2343 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2342 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2341 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2340 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2339 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2338 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2337 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2336 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2335 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2334 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2333 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2332 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2331 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2330 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2329 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2328 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2327 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2326 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2325 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2324 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2323 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2322 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2321 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2320 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2319 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2318 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2317 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2316 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2315 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2314 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2313 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2312 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2311 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2310 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2309 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2308 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2307 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2306 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2305 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2304 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2303 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2302 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2301 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2300 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2299 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2298 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2297 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2296 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2295 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2294 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2293 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2292 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2291 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2290 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2289 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2288 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2287 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2286 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2285 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2284 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2283 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2282 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2281 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2280 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2279 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2278 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2277 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2276 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2275 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2274 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2273 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2272 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2271 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2270 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2269 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2268 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2267 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2266 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2265 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2264 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2263 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2262 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2261 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2260 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2259 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2258 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2257 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2256 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2255 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2254 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2253 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2252 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2251 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2250 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2249 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2248 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2247 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2246 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2245 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2244 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2243 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2242 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2241 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2240 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2239 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2238 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2237 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2236 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2235 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2234 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2233 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2232 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2231 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2230 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2229 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2228 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2227 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2226 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2225 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2224 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2223 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2222 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2221 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2220 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2219 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2218 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2217 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2216 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2215 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2214 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2213 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2212 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2211 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2210 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2209 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2208 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2207 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2206 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2205 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2204 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2203 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2202 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2201 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2200 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2199 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2198 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2197 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2196 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2195 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2194 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2193 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2192 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2191 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2190 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2189 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2188 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2187 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2186 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2185 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2184 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2183 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2182 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2181 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2180 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2179 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2178 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2177 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2176 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2175 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2174 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2173 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2172 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2171 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2170 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2169 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2168 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2167 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2166 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2165 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2164 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2163 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2162 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2161 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2160 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2159 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2158 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2157 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2156 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2155 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2154 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2153 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2152 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2151 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2150 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2149 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2148 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2147 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2146 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2145 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2144 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2143 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2142 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2141 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2140 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2139 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2138 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2137 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2136 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2135 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2134 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2133 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2132 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2131 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2130 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2129 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2128 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2127 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2126 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2125 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2124 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2123 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2122 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2121 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2120 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2119 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2118 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2117 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2116 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2115 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2114 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2113 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2112 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2111 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2110 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2109 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2108 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2107 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2106 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2105 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2104 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2103 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2102 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2101 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2100 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2099 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2098 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2097 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2096 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2095 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2094 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2093 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2092 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2091 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2090 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2089 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2088 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2087 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2086 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2085 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2084 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2083 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2082 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2081 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2080 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2079 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2078 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2077 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2076 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2075 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2074 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2073 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2072 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2071 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2070 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2069 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2068 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2067 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2066 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2065 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2064 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2063 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2062 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2061 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2060 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2059 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2058 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2057 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2056 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2055 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2054 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2053 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2052 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2051 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2050 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2049 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2048 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2047 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2046 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2045 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2044 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2043 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2042 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2041 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2040 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2039 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2038 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2037 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2036 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2035 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2034 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2033 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2032 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2031 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2030 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2029 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2028 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2027 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2026 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2025 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2024 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2023 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2022 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2021 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2020 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2019 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2018 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2017 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2016 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2015 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2014 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2013 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2012 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2011 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2010 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2009 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2008 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2007 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2006 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2005 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2004 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2003 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2002 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2001 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2000 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1999 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1998 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1997 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1996 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1995 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1994 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1993 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1992 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1991 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1990 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1989 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1988 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1987 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1986 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1985 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1984 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1983 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1982 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1981 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1980 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1979 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1978 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1977 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1976 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1975 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1974 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1973 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1972 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1971 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1970 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1969 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1968 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1967 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1966 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1965 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1964 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1963 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1962 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1961 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1960 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1959 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1958 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1957 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1956 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1955 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1954 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1953 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1952 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1951 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1950 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1949 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1948 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1947 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1946 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1945 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1944 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1943 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1942 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1941 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1940 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1939 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1938 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1937 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1936 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1935 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1934 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1933 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1932 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1931 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1930 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1929 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1928 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1927 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1924 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1923 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1922 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1921 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1920 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1919 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1918 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1917 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1916 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1915 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1914 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1913 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1912 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1911 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1910 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1909 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1908 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1907 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1906 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1905 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1904 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1903 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1902 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1901 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1900 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1899 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1898 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1897 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1896 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1895 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1894 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1892 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1891 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1890 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1889 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1888 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1887 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1886 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1885 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1884 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1883 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1882 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1881 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1880 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1879 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1878 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1877 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1876 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1875 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1874 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1873 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1872 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1871 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1870 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1869 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1868 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1867 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1866 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1865 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1864 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1863 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1862 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1861 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1859 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1856 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1855 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1854 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1853 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1852 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1851 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1850 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1849 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1848 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1847 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1846 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1845 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1844 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1843 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1842 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1841 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1840 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1839 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1838 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1837 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1836 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1835 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1834 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1833 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1832 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1831 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1830 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1829 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1828 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1827 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1826 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1824 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1822 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1821 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1820 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1819 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1818 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1817 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1816 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1815 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1814 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1813 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1812 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1811 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1810 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1809 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1808 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1807 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1806 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1805 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1804 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1803 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1802 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1801 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1800 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1799 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1798 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1797 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1796 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1795 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1794 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1793 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1792 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1790 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1789 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1788 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1787 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1786 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1785 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1784 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1783 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1782 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1781 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1780 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1779 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1778 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1777 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1776 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1775 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1774 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1773 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1772 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1771 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1770 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1769 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1768 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1767 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1766 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1765 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1764 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1763 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1762 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1761 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1760 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1759 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1757 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1754 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1753 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1752 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1751 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1750 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1749 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1748 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1747 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1746 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1745 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1744 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1743 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1742 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1741 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1740 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1739 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1738 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1737 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1736 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1735 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1734 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1733 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1732 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1731 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1730 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1729 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1728 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1727 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1726 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1725 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1724 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1722 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1721 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1720 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1719 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1718 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1717 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1716 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1715 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1714 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1713 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1712 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1711 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1710 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1709 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1708 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1707 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1706 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1705 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1704 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1703 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1702 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1701 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1700 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1699 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1698 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1697 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1696 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1695 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1694 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1693 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1692 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1691 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1689 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1685 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1684 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1683 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1682 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1681 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1680 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1679 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1678 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1677 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1676 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1675 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1674 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1673 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1672 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1671 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1670 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1669 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1668 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1667 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1666 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1665 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1664 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1663 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1662 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1661 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1660 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1659 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1658 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1657 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1656 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1655 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1653 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1652 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1651 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1650 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1649 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1648 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1647 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1646 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1645 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1644 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1643 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1642 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1641 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1640 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1639 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1638 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1637 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1636 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1635 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1634 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1633 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1632 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1631 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1630 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1629 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1628 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1627 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1626 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1625 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1624 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1623 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1622 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1620 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1619 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1618 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1617 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1616 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1615 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1614 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1613 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1612 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1611 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1610 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1609 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1608 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1607 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1606 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1605 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1604 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1603 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1602 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1601 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1600 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1599 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1598 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1597 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1596 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1595 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1594 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1593 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1592 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1591 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1590 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1589 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1587 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1584 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1583 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1582 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1581 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1580 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1579 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1578 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1577 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1576 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1575 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1574 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1573 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1572 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1571 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1570 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1569 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1568 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1567 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1566 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1565 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1564 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1563 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1562 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1561 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1560 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1559 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1558 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1557 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1556 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1555 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1554 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1552 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1551 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1550 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1549 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1548 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1547 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1546 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1545 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1544 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1543 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1542 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1541 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1540 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1539 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1538 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1537 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1536 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1535 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1534 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1533 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1532 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1531 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1530 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1529 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1528 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1527 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1526 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1525 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1524 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1523 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1522 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1521 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1519 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1515 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1514 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1513 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1512 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1511 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1510 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1509 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1508 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1507 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1506 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1505 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1504 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1503 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1502 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1501 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1500 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1499 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1498 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1497 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1496 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1495 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1494 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1493 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1492 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1491 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1490 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1489 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1488 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1487 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1486 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1485 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1483 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1482 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1481 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1480 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1479 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1478 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1477 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1476 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1475 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1474 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1473 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1472 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1471 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1470 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1469 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1468 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1467 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1466 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1465 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1464 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1463 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1462 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1461 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1460 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1459 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1458 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1457 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1456 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1455 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1454 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1453 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1452 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1450 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1449 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1448 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1447 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1446 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1445 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1444 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1443 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1442 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1441 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1440 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1439 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1438 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1437 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1436 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1435 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1434 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1433 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1432 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1431 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1430 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1429 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1428 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1427 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1426 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1425 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1424 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1423 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1422 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1421 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1420 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1419 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1417 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1416 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1415 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1414 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1413 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1412 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1411 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1410 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1409 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1408 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1407 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1406 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1405 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1404 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1403 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1402 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1401 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1400 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1399 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1398 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1397 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1396 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1395 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1394 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1393 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1392 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1391 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1390 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1389 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1388 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1387 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1386 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1384 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1383 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1382 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1381 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1380 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1379 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1378 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1377 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1376 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1375 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1374 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1373 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1372 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1371 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1370 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1369 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1368 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1367 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1366 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1365 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1364 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1363 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1362 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1361 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1360 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1359 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1358 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1357 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1356 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1355 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1354 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1353 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1352 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1350 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1349 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1347 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1344 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1342 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1341 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1339 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1338 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1337 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1336 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1335 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1334 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1333 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1332 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1331 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1330 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1329 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1328 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1327 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1326 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1325 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1324 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1323 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1322 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1321 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1320 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1319 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1318 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1317 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1316 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1315 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1314 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1313 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1312 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1311 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1310 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1309 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1308 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1306 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1305 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1304 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1303 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1302 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1301 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1300 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1299 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1298 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1297 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1296 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1295 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1294 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1293 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1292 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1291 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1290 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1289 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1288 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1287 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1286 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1285 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1284 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1283 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1282 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1281 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1280 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1279 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1278 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1277 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1276 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1275 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1274 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1272 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1271 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1270 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1269 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1268 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1267 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1266 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1265 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1264 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1263 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1262 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1261 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1260 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1259 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1258 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1257 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1256 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1255 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1254 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1253 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1252 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1251 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1250 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1249 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1248 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1247 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1246 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1245 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1244 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1243 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1242 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1241 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1240 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1239 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1237 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1201 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1199 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1198 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1197 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1196 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1195 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1194 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1193 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1192 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1191 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1190 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1153 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1152 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1151 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1150 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1149 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1148 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1147 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1146 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1145 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1144 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1143 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1142 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1141 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1140 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1139 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1138 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1137 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1136 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1135 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1134 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1133 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1132 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1131 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1130 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1129 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1128 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1127 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1126 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1125 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1124 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1123 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1122 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1121 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1120 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1119 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1118 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1117 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1116 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1115 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1114 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1113 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1112 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1111 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1110 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1109 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1108 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1107 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1106 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1105 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1104 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1103 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1102 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1101 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1100 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1099 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1098 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1097 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1096 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1095 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1094 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1093 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1092 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1091 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1090 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1089 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1088 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1087 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1086 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1085 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1084 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1083 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1082 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1081 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1080 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1079 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1078 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1077 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1076 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1075 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1074 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1073 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1072 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1071 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1070 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1069 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1068 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1067 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1066 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1065 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1064 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1063 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1062 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1061 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1060 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1059 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1058 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1057 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1056 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1055 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1054 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1053 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1052 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1051 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1050 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1049 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1048 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1047 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1046 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1045 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1044 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1043 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1042 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1041 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1040 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1039 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1038 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1037 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1036 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1035 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1034 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1033 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1032 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1031 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1030 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1029 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1028 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1027 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1026 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1025 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1024 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1023 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1022 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1021 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1020 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1019 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1018 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1017 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1016 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1015 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1014 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1013 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1012 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1011 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1010 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1009 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1008 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1007 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1006 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1005 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1004 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1003 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1002 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1001 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n1000 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n999 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n998 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n997 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n996 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n995 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n994 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n993 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n992 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n991 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n990 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n989 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n988 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n987 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n986 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n985 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n984 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n983 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n982 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n981 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n980 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n979 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n978 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n977 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n976 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n975 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n974 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n973 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n972 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n971 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n970 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n969 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n968 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n967 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n966 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n965 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n964 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n963 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n962 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n961 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n960 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n959 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n958 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n957 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n956 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n955 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n954 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n953 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n952 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n951 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n950 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n949 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n948 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n947 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n946 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n945 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n944 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n943 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n942 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n941 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n940 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n939 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n938 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n937 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n936 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n935 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n934 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n933 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n932 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n931 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n930 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n929 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n928 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n927 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n926 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n925 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n924 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n923 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n922 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n921 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n920 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n919 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n918 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n917 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n916 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n915 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n914 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n913 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n912 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n911 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n910 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n909 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n908 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n907 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n906 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n905 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n904 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n903 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n902 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n901 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n900 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n899 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n898 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n897 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n896 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n895 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n894 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n893 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n892 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n891 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n890 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n889 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n888 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n887 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n886 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n885 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n884 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n883 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n882 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n881 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n880 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n879 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n878 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n877 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n876 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n875 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n874 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n873 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n872 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n871 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n870 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n869 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n868 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n867 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n866 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n865 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n864 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n863 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n862 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n861 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n860 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n859 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n858 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n857 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n856 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n855 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n854 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n853 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n852 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n851 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n850 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n849 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n848 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n847 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n846 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n845 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n844 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n843 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n842 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n841 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n840 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n839 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n838 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n837 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n836 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n835 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n834 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n833 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n832 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n831 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n830 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n829 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n828 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n827 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n826 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n825 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n824 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n823 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n822 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n821 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n820 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n819 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n818 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n817 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n816 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n815 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n814 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n813 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n812 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n811 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n810 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n809 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n808 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n807 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n806 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n805 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n804 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n803 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n802 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n801 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n800 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n799 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n798 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n797 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n796 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n795 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n794 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n793 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n792 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n791 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n790 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n789 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n788 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n787 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n786 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n785 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n784 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n783 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n782 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n781 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n780 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n779 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n778 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n777 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n776 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n775 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n774 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n773 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n772 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n771 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n770 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n769 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n768 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n767 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n766 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n765 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n764 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n763 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n762 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n761 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n760 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n759 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n758 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n757 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n756 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n755 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n754 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n753 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n752 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n751 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n750 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n749 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n748 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n747 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n746 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n745 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n744 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n743 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n742 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n741 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n740 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n739 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n738 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n737 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n736 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n735 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n734 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n733 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n732 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n731 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n730 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n729 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n728 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n727 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n726 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n725 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n724 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n723 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n722 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n721 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n720 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n719 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n718 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n717 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n716 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n715 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n714 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n713 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n712 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n711 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n710 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n709 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n708 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n707 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n706 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n705 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n704 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n703 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n702 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n701 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n700 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n699 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n698 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n697 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n696 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n695 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n694 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n693 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n692 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n691 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n690 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n689 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n688 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n687 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n686 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n685 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n684 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n683 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n682 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n681 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n680 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n679 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n678 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n677 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n676 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n675 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n674 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n673 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n672 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n671 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n670 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n669 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n668 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n667 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n666 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n665 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n664 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n663 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n662 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n661 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n660 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n659 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n658 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n657 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n656 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n655 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n654 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n653 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n652 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n651 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n650 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n649 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n648 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n647 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n646 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n645 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n644 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n643 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n642 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n641 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n640 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n639 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n638 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n637 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n636 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n635 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n634 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n633 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n632 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n631 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n630 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n629 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n628 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n627 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n626 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n625 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n624 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n623 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n622 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n621 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n620 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n619 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n618 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n617 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n616 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n615 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n614 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n613 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n612 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n611 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n610 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n609 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n608 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n607 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n606 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n605 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n604 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n603 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n602 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n601 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n600 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n599 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n598 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n597 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n596 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n595 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n594 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n593 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n592 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n591 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n590 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n589 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n588 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n587 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n586 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n585 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n584 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n583 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n582 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n581 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n580 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n579 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n578 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n577 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n576 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n575 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n574 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n573 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n572 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n571 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n570 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n569 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n568 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n567 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n566 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n565 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n564 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n563 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n562 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n561 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n560 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n559 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n558 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n557 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n556 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n555 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n554 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n553 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n552 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n551 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n550 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n549 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n548 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n547 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n546 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n545 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n544 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n543 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n542 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n541 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n540 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n539 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n538 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n537 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n536 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n535 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n534 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n533 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n532 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n531 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n530 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n529 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n528 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n527 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n526 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n525 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n524 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n523 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n522 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n521 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n520 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n519 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n518 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n517 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n516 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n515 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n514 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n513 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n512 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n511 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n510 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n509 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n508 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n507 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n506 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n505 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n504 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n503 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n502 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n501 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n500 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n499 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n498 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n497 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n496 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n495 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n494 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n493 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n492 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n491 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n490 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n489 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n488 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n487 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n486 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n485 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n484 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n483 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n482 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n481 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n480 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n479 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n478 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n477 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n476 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n475 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n474 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n473 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n472 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n471 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n470 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n469 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n468 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n467 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n466 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n465 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n464 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n463 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n462 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n461 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n460 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n459 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n458 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n457 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n456 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n455 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n454 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n453 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n452 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n451 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n450 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n449 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n448 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n447 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n446 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n445 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n444 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n443 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n442 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n441 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n440 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n439 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n438 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n437 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n436 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n435 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n434 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n433 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n432 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n431 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n430 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n429 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n428 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n427 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n426 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n425 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n424 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n423 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n422 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n421 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n420 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n419 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n418 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n417 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n416 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n415 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n414 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n413 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n412 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n411 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n410 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n409 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n408 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n407 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n406 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n405 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n404 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n403 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n402 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n401 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n400 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n399 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n398 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n397 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n396 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n395 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n394 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n393 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n392 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n391 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n390 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n389 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n388 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n387 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n386 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n385 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n384 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n383 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n382 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n381 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n380 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n379 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n378 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n377 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n376 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n375 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n374 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n373 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n372 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n371 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n370 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n369 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n368 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n367 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n366 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n365 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n364 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n363 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n362 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n361 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n360 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n359 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n358 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n357 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n356 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n355 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n354 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n353 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n352 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n351 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n350 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n349 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n348 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n347 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n346 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n345 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n344 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n343 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n342 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n341 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n340 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n339 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n338 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n337 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n336 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n335 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n334 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n333 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n332 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n331 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n330 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n329 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n328 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n327 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n326 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n325 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n324 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n323 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n322 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n321 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n320 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n319 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n318 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n317 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n316 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n315 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n314 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n313 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n312 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n311 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n310 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n309 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n308 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n307 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n306 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n305 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n304 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n303 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n302 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n301 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n300 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n299 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n298 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n297 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n296 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n295 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n294 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n293 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n292 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n291 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n290 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n289 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n288 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n287 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n286 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n285 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n284 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n283 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n282 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n281 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n280 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n279 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n278 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n277 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n276 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n275 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n274 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n273 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n272 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n271 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n270 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n269 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n268 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n267 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n266 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n265 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n264 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n263 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n262 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n261 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n260 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n259 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n258 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n257 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n256 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n255 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n254 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n253 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n252 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n251 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n250 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n249 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n248 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n247 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n246 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n245 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n244 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n243 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n242 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n241 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n240 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n239 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n238 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n237 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n236 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n235 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n234 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n233 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n232 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n231 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n230 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n229 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n228 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n227 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n226 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n225 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n224 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n223 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n222 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n221 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n220 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n219 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n218 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n217 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n216 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n215 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n214 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n213 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n212 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n211 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n210 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n209 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n208 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n207 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n206 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n205 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n204 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n203 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n202 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n201 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n200 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n199 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n198 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n197 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n196 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n195 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n194 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n193 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n192 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n191 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n190 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n189 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n188 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n187 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n186 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n185 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n184 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n183 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n182 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n181 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n180 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n179 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n178 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n177 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n176 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n175 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n174 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n173 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n172 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n171 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n170 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n169 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n168 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n167 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n166 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n165 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n164 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n163 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n162 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n161 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n160 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n159 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n158 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n157 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n156 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n155 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n154 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n153 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n152 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n151 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n150 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n149 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n148 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n147 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n146 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n145 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n144 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n143 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n142 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n141 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n140 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n139 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n138 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n137 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n136 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n135 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n134 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n133 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n132 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n131 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n130 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n129 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n128 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n127 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n126 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n125 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n124 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n123 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n122 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n121 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n120 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n119 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n118 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n117 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n116 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n115 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n114 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n113 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n112 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n111 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n110 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n109 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n108 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n107 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n106 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n105 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n104 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n103 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n102 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n101 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n100 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n99 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n98 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n97 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n96 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n95 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n94 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n93 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n92 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n91 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n90 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n89 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n88 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n87 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n86 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n85 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n84 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n83 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n82 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n81 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n80 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n79 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n78 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n77 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n76 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n75 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n74 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n73 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n72 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n71 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n70 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n69 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n68 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n67 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n66 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n65 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n64 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n63 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n62 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n61 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n60 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n59 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n58 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n57 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n56 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n55 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n54 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n53 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n52 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n51 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n50 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n49 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n48 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n47 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n46 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n45 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n44 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n43 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n42 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n41 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n40 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n39 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n38 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n37 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n36 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n35 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n34 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n33 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n32 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n31 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n30 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n29 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n28 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n27 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n26 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n25 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n24 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n23 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n22 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n21 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n20 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n19 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n18 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n17 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n16 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n15 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n14 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n13 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n12 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n11 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n10 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n9 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n8 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n7 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n6 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n5 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n4 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n3 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/n2 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N429 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N428 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N427 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N426 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N425 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N424 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N423 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N422 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N421 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N420 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N419 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N418 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N417 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N416 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N415 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N414 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N413 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N412 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N411 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N410 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N409 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N408 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N407 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N406 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N405 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N404 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N403 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N402 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N401 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N400 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N399 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N398 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N397 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N396 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N359 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N358 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N357 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N356 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N355 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N354 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N353 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N352 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N351 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N350 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N349 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N348 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N347 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N346 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N345 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N344 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N343 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N342 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N341 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N340 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N339 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N338 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N337 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N336 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N335 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N334 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N333 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N332 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N331 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N330 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N329 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/N328 ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][31] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][0] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][1] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][2] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][3] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][4] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][5] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][6] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][7] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][8] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][9] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][10] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][11] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][12] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][13] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][14] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][15] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][16] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][17] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][18] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][19] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][20] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][21] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][22] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][23] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][24] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][25] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][26] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][27] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][28] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][29] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][30] ,
         \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][31] ,
         \dp/ex_stage/n10 , \dp/ex_stage/n9 , \dp/ex_stage/n8 ,
         \dp/ex_stage/n7 , \dp/ex_stage/n6 , \dp/ex_stage/n5 ,
         \dp/ex_stage/n4 , \dp/ex_stage/n3 , \dp/ex_stage/n2 ,
         \dp/ex_stage/n1 , \dp/ex_stage/muxA/n110 , \dp/ex_stage/muxA/n109 ,
         \dp/ex_stage/muxA/n108 , \dp/ex_stage/muxA/n107 ,
         \dp/ex_stage/muxA/n106 , \dp/ex_stage/muxA/n105 ,
         \dp/ex_stage/muxA/n104 , \dp/ex_stage/muxA/n103 ,
         \dp/ex_stage/muxA/n102 , \dp/ex_stage/muxA/n101 ,
         \dp/ex_stage/muxA/n100 , \dp/ex_stage/muxA/n99 ,
         \dp/ex_stage/muxA/n98 , \dp/ex_stage/muxA/n97 ,
         \dp/ex_stage/muxA/n96 , \dp/ex_stage/muxA/n95 ,
         \dp/ex_stage/muxA/n94 , \dp/ex_stage/muxA/n93 ,
         \dp/ex_stage/muxA/n92 , \dp/ex_stage/muxA/n91 ,
         \dp/ex_stage/muxA/n90 , \dp/ex_stage/muxA/n89 ,
         \dp/ex_stage/muxA/n88 , \dp/ex_stage/muxA/n87 ,
         \dp/ex_stage/muxA/n86 , \dp/ex_stage/muxA/n85 ,
         \dp/ex_stage/muxA/n84 , \dp/ex_stage/muxA/n83 ,
         \dp/ex_stage/muxA/n82 , \dp/ex_stage/muxA/n81 ,
         \dp/ex_stage/muxA/n80 , \dp/ex_stage/muxA/n79 ,
         \dp/ex_stage/muxA/n14 , \dp/ex_stage/muxA/n13 ,
         \dp/ex_stage/muxA/n12 , \dp/ex_stage/muxA/n11 ,
         \dp/ex_stage/muxA/n10 , \dp/ex_stage/muxA/n9 , \dp/ex_stage/muxA/n8 ,
         \dp/ex_stage/muxA/n7 , \dp/ex_stage/muxA/n6 , \dp/ex_stage/muxA/n5 ,
         \dp/ex_stage/muxA/n4 , \dp/ex_stage/muxA/n3 , \dp/ex_stage/muxA/n2 ,
         \dp/ex_stage/muxA/n1 , \dp/ex_stage/muxB/n110 ,
         \dp/ex_stage/muxB/n109 , \dp/ex_stage/muxB/n108 ,
         \dp/ex_stage/muxB/n107 , \dp/ex_stage/muxB/n106 ,
         \dp/ex_stage/muxB/n105 , \dp/ex_stage/muxB/n104 ,
         \dp/ex_stage/muxB/n103 , \dp/ex_stage/muxB/n102 ,
         \dp/ex_stage/muxB/n101 , \dp/ex_stage/muxB/n100 ,
         \dp/ex_stage/muxB/n99 , \dp/ex_stage/muxB/n98 ,
         \dp/ex_stage/muxB/n97 , \dp/ex_stage/muxB/n96 ,
         \dp/ex_stage/muxB/n95 , \dp/ex_stage/muxB/n94 ,
         \dp/ex_stage/muxB/n93 , \dp/ex_stage/muxB/n92 ,
         \dp/ex_stage/muxB/n91 , \dp/ex_stage/muxB/n90 ,
         \dp/ex_stage/muxB/n89 , \dp/ex_stage/muxB/n88 ,
         \dp/ex_stage/muxB/n87 , \dp/ex_stage/muxB/n86 ,
         \dp/ex_stage/muxB/n85 , \dp/ex_stage/muxB/n84 ,
         \dp/ex_stage/muxB/n83 , \dp/ex_stage/muxB/n82 ,
         \dp/ex_stage/muxB/n81 , \dp/ex_stage/muxB/n80 ,
         \dp/ex_stage/muxB/n79 , \dp/ex_stage/muxB/n14 ,
         \dp/ex_stage/muxB/n13 , \dp/ex_stage/muxB/n12 ,
         \dp/ex_stage/muxB/n11 , \dp/ex_stage/muxB/n10 , \dp/ex_stage/muxB/n9 ,
         \dp/ex_stage/muxB/n8 , \dp/ex_stage/muxB/n7 , \dp/ex_stage/muxB/n6 ,
         \dp/ex_stage/muxB/n5 , \dp/ex_stage/muxB/n4 , \dp/ex_stage/muxB/n3 ,
         \dp/ex_stage/muxB/n2 , \dp/ex_stage/muxB/n1 , \dp/ex_stage/alu/n227 ,
         \dp/ex_stage/alu/n226 , \dp/ex_stage/alu/n225 ,
         \dp/ex_stage/alu/n224 , \dp/ex_stage/alu/n223 ,
         \dp/ex_stage/alu/n222 , \dp/ex_stage/alu/n221 ,
         \dp/ex_stage/alu/n220 , \dp/ex_stage/alu/n219 ,
         \dp/ex_stage/alu/n218 , \dp/ex_stage/alu/n217 ,
         \dp/ex_stage/alu/n216 , \dp/ex_stage/alu/n215 ,
         \dp/ex_stage/alu/n214 , \dp/ex_stage/alu/n213 ,
         \dp/ex_stage/alu/n212 , \dp/ex_stage/alu/n211 ,
         \dp/ex_stage/alu/n210 , \dp/ex_stage/alu/n209 , \dp/ex_stage/alu/n87 ,
         \dp/ex_stage/alu/n86 , \dp/ex_stage/alu/n85 , \dp/ex_stage/alu/n84 ,
         \dp/ex_stage/alu/n83 , \dp/ex_stage/alu/n82 , \dp/ex_stage/alu/n81 ,
         \dp/ex_stage/alu/n80 , \dp/ex_stage/alu/n79 , \dp/ex_stage/alu/n78 ,
         \dp/ex_stage/alu/n77 , \dp/ex_stage/alu/n76 , \dp/ex_stage/alu/n75 ,
         \dp/ex_stage/alu/n74 , \dp/ex_stage/alu/n73 , \dp/ex_stage/alu/n72 ,
         \dp/ex_stage/alu/n71 , \dp/ex_stage/alu/n70 , \dp/ex_stage/alu/n69 ,
         \dp/ex_stage/alu/n68 , \dp/ex_stage/alu/n67 , \dp/ex_stage/alu/n66 ,
         \dp/ex_stage/alu/n65 , \dp/ex_stage/alu/n64 , \dp/ex_stage/alu/n63 ,
         \dp/ex_stage/alu/n62 , \dp/ex_stage/alu/n61 , \dp/ex_stage/alu/n60 ,
         \dp/ex_stage/alu/n59 , \dp/ex_stage/alu/n58 , \dp/ex_stage/alu/n57 ,
         \dp/ex_stage/alu/n56 , \dp/ex_stage/alu/n55 , \dp/ex_stage/alu/n54 ,
         \dp/ex_stage/alu/n53 , \dp/ex_stage/alu/n52 , \dp/ex_stage/alu/n51 ,
         \dp/ex_stage/alu/n50 , \dp/ex_stage/alu/n49 , \dp/ex_stage/alu/n48 ,
         \dp/ex_stage/alu/n47 , \dp/ex_stage/alu/n46 , \dp/ex_stage/alu/n45 ,
         \dp/ex_stage/alu/n44 , \dp/ex_stage/alu/n43 , \dp/ex_stage/alu/n42 ,
         \dp/ex_stage/alu/n41 , \dp/ex_stage/alu/n40 , \dp/ex_stage/alu/n39 ,
         \dp/ex_stage/alu/n38 , \dp/ex_stage/alu/n37 , \dp/ex_stage/alu/n36 ,
         \dp/ex_stage/alu/n35 , \dp/ex_stage/alu/n34 , \dp/ex_stage/alu/n33 ,
         \dp/ex_stage/alu/n32 , \dp/ex_stage/alu/n31 , \dp/ex_stage/alu/n30 ,
         \dp/ex_stage/alu/n29 , \dp/ex_stage/alu/n28 , \dp/ex_stage/alu/n27 ,
         \dp/ex_stage/alu/n26 , \dp/ex_stage/alu/n25 , \dp/ex_stage/alu/n24 ,
         \dp/ex_stage/alu/n23 , \dp/ex_stage/alu/n22 , \dp/ex_stage/alu/n21 ,
         \dp/ex_stage/alu/n20 , \dp/ex_stage/alu/n19 , \dp/ex_stage/alu/n18 ,
         \dp/ex_stage/alu/n17 , \dp/ex_stage/alu/n16 , \dp/ex_stage/alu/n15 ,
         \dp/ex_stage/alu/n14 , \dp/ex_stage/alu/n11 , \dp/ex_stage/alu/n10 ,
         \dp/ex_stage/alu/n9 , \dp/ex_stage/alu/n8 , \dp/ex_stage/alu/n7 ,
         \dp/ex_stage/alu/n6 , \dp/ex_stage/alu/n5 , \dp/ex_stage/alu/n4 ,
         \dp/ex_stage/alu/n3 , \dp/ex_stage/alu/n2 , \dp/ex_stage/alu/n1 ,
         \dp/ex_stage/alu/n208 , \dp/ex_stage/alu/n207 ,
         \dp/ex_stage/alu/n206 , \dp/ex_stage/alu/n205 ,
         \dp/ex_stage/alu/n204 , \dp/ex_stage/alu/n203 ,
         \dp/ex_stage/alu/n202 , \dp/ex_stage/alu/n201 ,
         \dp/ex_stage/alu/n200 , \dp/ex_stage/alu/n199 ,
         \dp/ex_stage/alu/n198 , \dp/ex_stage/alu/n197 ,
         \dp/ex_stage/alu/n196 , \dp/ex_stage/alu/n195 ,
         \dp/ex_stage/alu/n194 , \dp/ex_stage/alu/n193 ,
         \dp/ex_stage/alu/n192 , \dp/ex_stage/alu/n191 ,
         \dp/ex_stage/alu/n190 , \dp/ex_stage/alu/n189 ,
         \dp/ex_stage/alu/n188 , \dp/ex_stage/alu/n187 ,
         \dp/ex_stage/alu/n186 , \dp/ex_stage/alu/n185 ,
         \dp/ex_stage/alu/n184 , \dp/ex_stage/alu/n183 ,
         \dp/ex_stage/alu/n182 , \dp/ex_stage/alu/n181 ,
         \dp/ex_stage/alu/n180 , \dp/ex_stage/alu/n179 ,
         \dp/ex_stage/alu/n178 , \dp/ex_stage/alu/n177 ,
         \dp/ex_stage/alu/n176 , \dp/ex_stage/alu/n175 ,
         \dp/ex_stage/alu/n174 , \dp/ex_stage/alu/n173 ,
         \dp/ex_stage/alu/n172 , \dp/ex_stage/alu/n171 ,
         \dp/ex_stage/alu/n170 , \dp/ex_stage/alu/n169 ,
         \dp/ex_stage/alu/n168 , \dp/ex_stage/alu/n167 ,
         \dp/ex_stage/alu/n166 , \dp/ex_stage/alu/n165 ,
         \dp/ex_stage/alu/n164 , \dp/ex_stage/alu/n163 ,
         \dp/ex_stage/alu/n162 , \dp/ex_stage/alu/n161 ,
         \dp/ex_stage/alu/n160 , \dp/ex_stage/alu/n159 ,
         \dp/ex_stage/alu/n158 , \dp/ex_stage/alu/n157 ,
         \dp/ex_stage/alu/n156 , \dp/ex_stage/alu/n155 ,
         \dp/ex_stage/alu/n154 , \dp/ex_stage/alu/n153 ,
         \dp/ex_stage/alu/n152 , \dp/ex_stage/alu/n151 ,
         \dp/ex_stage/alu/n150 , \dp/ex_stage/alu/n149 ,
         \dp/ex_stage/alu/n148 , \dp/ex_stage/alu/n147 ,
         \dp/ex_stage/alu/n146 , \dp/ex_stage/alu/n145 ,
         \dp/ex_stage/alu/n144 , \dp/ex_stage/alu/n143 ,
         \dp/ex_stage/alu/n142 , \dp/ex_stage/alu/n141 ,
         \dp/ex_stage/alu/n140 , \dp/ex_stage/alu/n139 ,
         \dp/ex_stage/alu/n138 , \dp/ex_stage/alu/n137 ,
         \dp/ex_stage/alu/n136 , \dp/ex_stage/alu/n135 ,
         \dp/ex_stage/alu/n134 , \dp/ex_stage/alu/n133 ,
         \dp/ex_stage/alu/n132 , \dp/ex_stage/alu/n131 ,
         \dp/ex_stage/alu/n130 , \dp/ex_stage/alu/n129 ,
         \dp/ex_stage/alu/n128 , \dp/ex_stage/alu/n127 ,
         \dp/ex_stage/alu/n126 , \dp/ex_stage/alu/n125 ,
         \dp/ex_stage/alu/n124 , \dp/ex_stage/alu/n123 ,
         \dp/ex_stage/alu/n122 , \dp/ex_stage/alu/n121 ,
         \dp/ex_stage/alu/n120 , \dp/ex_stage/alu/n119 ,
         \dp/ex_stage/alu/n118 , \dp/ex_stage/alu/n117 ,
         \dp/ex_stage/alu/n116 , \dp/ex_stage/alu/n115 ,
         \dp/ex_stage/alu/n114 , \dp/ex_stage/alu/n113 ,
         \dp/ex_stage/alu/n112 , \dp/ex_stage/alu/n111 ,
         \dp/ex_stage/alu/n110 , \dp/ex_stage/alu/n109 ,
         \dp/ex_stage/alu/n108 , \dp/ex_stage/alu/n107 ,
         \dp/ex_stage/alu/n106 , \dp/ex_stage/alu/n105 ,
         \dp/ex_stage/alu/n104 , \dp/ex_stage/alu/n103 ,
         \dp/ex_stage/alu/n102 , \dp/ex_stage/alu/n101 ,
         \dp/ex_stage/alu/n100 , \dp/ex_stage/alu/n99 , \dp/ex_stage/alu/n98 ,
         \dp/ex_stage/alu/n97 , \dp/ex_stage/alu/n96 , \dp/ex_stage/alu/n95 ,
         \dp/ex_stage/alu/n94 , \dp/ex_stage/alu/n93 , \dp/ex_stage/alu/n92 ,
         \dp/ex_stage/alu/n91 , \dp/ex_stage/alu/n90 , \dp/ex_stage/alu/n89 ,
         \dp/ex_stage/alu/n88 , \dp/ex_stage/alu/N23 ,
         \dp/ex_stage/alu/shift_arith_i , \dp/ex_stage/alu/N22 ,
         \dp/ex_stage/alu/N21 , \dp/ex_stage/alu/N20 , \dp/ex_stage/alu/N19 ,
         \dp/ex_stage/alu/N18 , \dp/ex_stage/alu/N17 , \dp/ex_stage/alu/N16 ,
         \dp/ex_stage/alu/adder/n3 , \dp/ex_stage/alu/adder/n2 ,
         \dp/ex_stage/alu/adder/n1 , \dp/ex_stage/alu/adder/B_xor[0] ,
         \dp/ex_stage/alu/adder/B_xor[1] , \dp/ex_stage/alu/adder/B_xor[2] ,
         \dp/ex_stage/alu/adder/B_xor[3] , \dp/ex_stage/alu/adder/B_xor[4] ,
         \dp/ex_stage/alu/adder/B_xor[5] , \dp/ex_stage/alu/adder/B_xor[6] ,
         \dp/ex_stage/alu/adder/B_xor[7] , \dp/ex_stage/alu/adder/B_xor[8] ,
         \dp/ex_stage/alu/adder/B_xor[9] , \dp/ex_stage/alu/adder/B_xor[10] ,
         \dp/ex_stage/alu/adder/B_xor[11] , \dp/ex_stage/alu/adder/B_xor[12] ,
         \dp/ex_stage/alu/adder/B_xor[13] , \dp/ex_stage/alu/adder/B_xor[14] ,
         \dp/ex_stage/alu/adder/B_xor[15] , \dp/ex_stage/alu/adder/B_xor[16] ,
         \dp/ex_stage/alu/adder/B_xor[17] , \dp/ex_stage/alu/adder/B_xor[18] ,
         \dp/ex_stage/alu/adder/B_xor[19] , \dp/ex_stage/alu/adder/B_xor[20] ,
         \dp/ex_stage/alu/adder/B_xor[21] , \dp/ex_stage/alu/adder/B_xor[22] ,
         \dp/ex_stage/alu/adder/B_xor[23] , \dp/ex_stage/alu/adder/B_xor[24] ,
         \dp/ex_stage/alu/adder/B_xor[25] , \dp/ex_stage/alu/adder/B_xor[26] ,
         \dp/ex_stage/alu/adder/B_xor[27] , \dp/ex_stage/alu/adder/B_xor[28] ,
         \dp/ex_stage/alu/adder/B_xor[29] , \dp/ex_stage/alu/adder/B_xor[30] ,
         \dp/ex_stage/alu/adder/B_xor[31] , \dp/ex_stage/alu/adder/Cout ,
         \dp/ex_stage/alu/adder/SparseTree/prop[2][2] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[3][3] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[4][3] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[4][4] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[5][5] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[6][5] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[6][6] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[7][7] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[8][5] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[8][7] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[8][8] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[9][9] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[10][9] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[10][10] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[11][11] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[12][9] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[12][11] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[12][12] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[13][13] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[14][13] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[14][14] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[15][15] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[16][9] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[16][13] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[16][15] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[16][16] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[17][17] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[18][17] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[18][18] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[19][19] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[20][17] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[20][19] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[20][20] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[21][21] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[22][21] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[22][22] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[23][23] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[24][17] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[24][21] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[24][23] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[24][24] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[25][25] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[26][25] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[26][26] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[27][27] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[28][17] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[28][25] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[28][27] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[28][28] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[29][29] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[30][29] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[30][30] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[31][31] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[32][17] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[32][25] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[32][29] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[32][31] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[32][32] ,
         \dp/ex_stage/alu/adder/SparseTree/prop[1][1] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[2][0] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[2][2] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[3][3] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[4][3] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[4][4] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[5][5] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[6][5] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[6][6] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[7][7] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[8][5] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[8][7] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[8][8] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[9][9] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[10][9] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[10][10] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[11][11] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[12][9] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[12][11] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[12][12] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[13][13] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[14][13] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[14][14] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[15][15] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[16][9] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[16][13] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[16][15] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[16][16] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[17][17] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[18][17] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[18][18] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[19][19] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[20][17] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[20][19] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[20][20] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[21][21] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[22][21] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[22][22] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[23][23] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[24][17] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[24][21] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[24][23] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[24][24] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[25][25] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[26][25] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[26][26] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[27][27] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[28][17] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[28][25] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[28][27] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[28][28] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[29][29] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[30][29] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[30][30] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[31][31] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[32][17] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[32][25] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[32][29] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[32][31] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[32][32] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[1][0] ,
         \dp/ex_stage/alu/adder/SparseTree/gen[1][1] ,
         \dp/ex_stage/alu/adder/SparseTree/G10/n2 ,
         \dp/ex_stage/alu/adder/SparseTree/G20_1/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_0/n2 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_1/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_2/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_3/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_4/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_5/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_6/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_7/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_8/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_9/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_10/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_11/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_12/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_13/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_14/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_2/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_0/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_1/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_2/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_3/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_4/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_5/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_6/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_3/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_0/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_1/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_2/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_4/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/G_2n_0_4_1/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_0_0/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_1_0/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_5/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_1/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_2/n3 ,
         \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_3/n3 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n5 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n9 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n8 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n7 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n6 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n13 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n12 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n11 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n10 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n5 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n13 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n12 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n11 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n10 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n5 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n13 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n12 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n11 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n10 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n5 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n13 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n12 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n11 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n10 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n5 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n13 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n12 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n11 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n10 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n5 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n13 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n12 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n11 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n10 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n5 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[1] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[2] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[3] ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/Co ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n13 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n12 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n11 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n10 ,
         \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n5 ,
         \dp/ex_stage/alu/shifter/n101 , \dp/ex_stage/alu/shifter/n100 ,
         \dp/ex_stage/alu/shifter/n99 , \dp/ex_stage/alu/shifter/n98 ,
         \dp/ex_stage/alu/shifter/n97 , \dp/ex_stage/alu/shifter/n96 ,
         \dp/ex_stage/alu/shifter/n95 , \dp/ex_stage/alu/shifter/n94 ,
         \dp/ex_stage/alu/shifter/n93 , \dp/ex_stage/alu/shifter/n20 ,
         \dp/ex_stage/alu/shifter/n19 , \dp/ex_stage/alu/shifter/n12 ,
         \dp/ex_stage/alu/shifter/n11 , \dp/ex_stage/alu/shifter/n10 ,
         \dp/ex_stage/alu/shifter/n9 , \dp/ex_stage/alu/shifter/n8 ,
         \dp/ex_stage/alu/shifter/n7 , \dp/ex_stage/alu/shifter/n6 ,
         \dp/ex_stage/alu/shifter/n5 , \dp/ex_stage/alu/shifter/n4 ,
         \dp/ex_stage/alu/shifter/n3 , \dp/ex_stage/alu/shifter/n2 ,
         \dp/ex_stage/alu/shifter/n1 , \dp/ex_stage/alu/shifter/n92 ,
         \dp/ex_stage/alu/shifter/n91 , \dp/ex_stage/alu/shifter/n90 ,
         \dp/ex_stage/alu/shifter/n89 , \dp/ex_stage/alu/shifter/n88 ,
         \dp/ex_stage/alu/shifter/n87 , \dp/ex_stage/alu/shifter/n86 ,
         \dp/ex_stage/alu/shifter/n85 , \dp/ex_stage/alu/shifter/n84 ,
         \dp/ex_stage/alu/shifter/n83 , \dp/ex_stage/alu/shifter/n82 ,
         \dp/ex_stage/alu/shifter/n81 , \dp/ex_stage/alu/shifter/n80 ,
         \dp/ex_stage/alu/shifter/n79 , \dp/ex_stage/alu/shifter/n78 ,
         \dp/ex_stage/alu/shifter/n77 , \dp/ex_stage/alu/shifter/n76 ,
         \dp/ex_stage/alu/shifter/n75 , \dp/ex_stage/alu/shifter/n74 ,
         \dp/ex_stage/alu/shifter/n73 , \dp/ex_stage/alu/shifter/n72 ,
         \dp/ex_stage/alu/shifter/n71 , \dp/ex_stage/alu/shifter/n70 ,
         \dp/ex_stage/alu/shifter/n69 , \dp/ex_stage/alu/shifter/n68 ,
         \dp/ex_stage/alu/shifter/n67 , \dp/ex_stage/alu/shifter/n66 ,
         \dp/ex_stage/alu/shifter/n65 , \dp/ex_stage/alu/shifter/n64 ,
         \dp/ex_stage/alu/shifter/n63 , \dp/ex_stage/alu/shifter/n62 ,
         \dp/ex_stage/alu/shifter/n61 , \dp/ex_stage/alu/shifter/n60 ,
         \dp/ex_stage/alu/shifter/n59 , \dp/ex_stage/alu/shifter/n58 ,
         \dp/ex_stage/alu/shifter/n57 , \dp/ex_stage/alu/shifter/n56 ,
         \dp/ex_stage/alu/shifter/n55 , \dp/ex_stage/alu/shifter/n54 ,
         \dp/ex_stage/alu/shifter/n53 , \dp/ex_stage/alu/shifter/n52 ,
         \dp/ex_stage/alu/shifter/n51 , \dp/ex_stage/alu/shifter/n50 ,
         \dp/ex_stage/alu/shifter/n49 , \dp/ex_stage/alu/shifter/n48 ,
         \dp/ex_stage/alu/shifter/n47 , \dp/ex_stage/alu/shifter/n46 ,
         \dp/ex_stage/alu/shifter/n45 , \dp/ex_stage/alu/shifter/n44 ,
         \dp/ex_stage/alu/shifter/n43 , \dp/ex_stage/alu/shifter/n42 ,
         \dp/ex_stage/alu/shifter/n41 , \dp/ex_stage/alu/shifter/n40 ,
         \dp/ex_stage/alu/shifter/n39 , \dp/ex_stage/alu/shifter/n38 ,
         \dp/ex_stage/alu/shifter/n37 , \dp/ex_stage/alu/shifter/n36 ,
         \dp/ex_stage/alu/shifter/n35 , \dp/ex_stage/alu/shifter/n34 ,
         \dp/ex_stage/alu/shifter/n33 , \dp/ex_stage/alu/shifter/n32 ,
         \dp/ex_stage/alu/shifter/n31 , \dp/ex_stage/alu/shifter/n30 ,
         \dp/ex_stage/alu/shifter/n29 , \dp/ex_stage/alu/shifter/n28 ,
         \dp/ex_stage/alu/shifter/n27 , \dp/ex_stage/alu/shifter/n26 ,
         \dp/ex_stage/alu/shifter/n25 , \dp/ex_stage/alu/shifter/n24 ,
         \dp/ex_stage/alu/shifter/n23 , \dp/ex_stage/alu/shifter/n22 ,
         \dp/ex_stage/alu/shifter/n21 , \dp/ex_stage/alu/shifter/N265 ,
         \dp/ex_stage/alu/shifter/N264 , \dp/ex_stage/alu/shifter/N263 ,
         \dp/ex_stage/alu/shifter/N262 , \dp/ex_stage/alu/shifter/N261 ,
         \dp/ex_stage/alu/shifter/N260 , \dp/ex_stage/alu/shifter/N259 ,
         \dp/ex_stage/alu/shifter/N258 , \dp/ex_stage/alu/shifter/N257 ,
         \dp/ex_stage/alu/shifter/N256 , \dp/ex_stage/alu/shifter/N255 ,
         \dp/ex_stage/alu/shifter/N254 , \dp/ex_stage/alu/shifter/N253 ,
         \dp/ex_stage/alu/shifter/N252 , \dp/ex_stage/alu/shifter/N251 ,
         \dp/ex_stage/alu/shifter/N250 , \dp/ex_stage/alu/shifter/N249 ,
         \dp/ex_stage/alu/shifter/N248 , \dp/ex_stage/alu/shifter/N247 ,
         \dp/ex_stage/alu/shifter/N246 , \dp/ex_stage/alu/shifter/N245 ,
         \dp/ex_stage/alu/shifter/N244 , \dp/ex_stage/alu/shifter/N243 ,
         \dp/ex_stage/alu/shifter/N242 , \dp/ex_stage/alu/shifter/N241 ,
         \dp/ex_stage/alu/shifter/N240 , \dp/ex_stage/alu/shifter/N239 ,
         \dp/ex_stage/alu/shifter/N238 , \dp/ex_stage/alu/shifter/N237 ,
         \dp/ex_stage/alu/shifter/N236 , \dp/ex_stage/alu/shifter/N235 ,
         \dp/ex_stage/alu/shifter/N234 , \dp/ex_stage/alu/shifter/N233 ,
         \dp/ex_stage/alu/shifter/N232 , \dp/ex_stage/alu/shifter/N231 ,
         \dp/ex_stage/alu/shifter/N230 , \dp/ex_stage/alu/shifter/N229 ,
         \dp/ex_stage/alu/shifter/N228 , \dp/ex_stage/alu/shifter/N227 ,
         \dp/ex_stage/alu/shifter/N226 , \dp/ex_stage/alu/shifter/N225 ,
         \dp/ex_stage/alu/shifter/N224 , \dp/ex_stage/alu/shifter/N223 ,
         \dp/ex_stage/alu/shifter/N222 , \dp/ex_stage/alu/shifter/N221 ,
         \dp/ex_stage/alu/shifter/N220 , \dp/ex_stage/alu/shifter/N219 ,
         \dp/ex_stage/alu/shifter/N218 , \dp/ex_stage/alu/shifter/N217 ,
         \dp/ex_stage/alu/shifter/N216 , \dp/ex_stage/alu/shifter/N215 ,
         \dp/ex_stage/alu/shifter/N214 , \dp/ex_stage/alu/shifter/N213 ,
         \dp/ex_stage/alu/shifter/N212 , \dp/ex_stage/alu/shifter/N211 ,
         \dp/ex_stage/alu/shifter/N210 , \dp/ex_stage/alu/shifter/N209 ,
         \dp/ex_stage/alu/shifter/N208 , \dp/ex_stage/alu/shifter/N207 ,
         \dp/ex_stage/alu/shifter/N206 , \dp/ex_stage/alu/shifter/N205 ,
         \dp/ex_stage/alu/shifter/N204 , \dp/ex_stage/alu/shifter/N203 ,
         \dp/ex_stage/alu/shifter/N202 , \dp/ex_stage/alu/shifter/N168 ,
         \dp/ex_stage/alu/shifter/N167 , \dp/ex_stage/alu/shifter/N166 ,
         \dp/ex_stage/alu/shifter/N165 , \dp/ex_stage/alu/shifter/N164 ,
         \dp/ex_stage/alu/shifter/N163 , \dp/ex_stage/alu/shifter/N162 ,
         \dp/ex_stage/alu/shifter/N161 , \dp/ex_stage/alu/shifter/N160 ,
         \dp/ex_stage/alu/shifter/N159 , \dp/ex_stage/alu/shifter/N158 ,
         \dp/ex_stage/alu/shifter/N157 , \dp/ex_stage/alu/shifter/N156 ,
         \dp/ex_stage/alu/shifter/N155 , \dp/ex_stage/alu/shifter/N154 ,
         \dp/ex_stage/alu/shifter/N153 , \dp/ex_stage/alu/shifter/N152 ,
         \dp/ex_stage/alu/shifter/N151 , \dp/ex_stage/alu/shifter/N150 ,
         \dp/ex_stage/alu/shifter/N149 , \dp/ex_stage/alu/shifter/N148 ,
         \dp/ex_stage/alu/shifter/N147 , \dp/ex_stage/alu/shifter/N146 ,
         \dp/ex_stage/alu/shifter/N145 , \dp/ex_stage/alu/shifter/N144 ,
         \dp/ex_stage/alu/shifter/N143 , \dp/ex_stage/alu/shifter/N142 ,
         \dp/ex_stage/alu/shifter/N141 , \dp/ex_stage/alu/shifter/N140 ,
         \dp/ex_stage/alu/shifter/N139 , \dp/ex_stage/alu/shifter/N138 ,
         \dp/ex_stage/alu/shifter/N137 , \dp/ex_stage/alu/shifter/N136 ,
         \dp/ex_stage/alu/shifter/N135 , \dp/ex_stage/alu/shifter/N134 ,
         \dp/ex_stage/alu/shifter/N133 , \dp/ex_stage/alu/shifter/N132 ,
         \dp/ex_stage/alu/shifter/N131 , \dp/ex_stage/alu/shifter/N130 ,
         \dp/ex_stage/alu/shifter/N129 , \dp/ex_stage/alu/shifter/N128 ,
         \dp/ex_stage/alu/shifter/N127 , \dp/ex_stage/alu/shifter/N126 ,
         \dp/ex_stage/alu/shifter/N125 , \dp/ex_stage/alu/shifter/N124 ,
         \dp/ex_stage/alu/shifter/N123 , \dp/ex_stage/alu/shifter/N122 ,
         \dp/ex_stage/alu/shifter/N121 , \dp/ex_stage/alu/shifter/N120 ,
         \dp/ex_stage/alu/shifter/N119 , \dp/ex_stage/alu/shifter/N118 ,
         \dp/ex_stage/alu/shifter/N117 , \dp/ex_stage/alu/shifter/N116 ,
         \dp/ex_stage/alu/shifter/N115 , \dp/ex_stage/alu/shifter/N114 ,
         \dp/ex_stage/alu/shifter/N113 , \dp/ex_stage/alu/shifter/N112 ,
         \dp/ex_stage/alu/shifter/N111 , \dp/ex_stage/alu/shifter/N110 ,
         \dp/ex_stage/alu/shifter/N109 , \dp/ex_stage/alu/shifter/N108 ,
         \dp/ex_stage/alu/shifter/N107 , \dp/ex_stage/alu/shifter/N106 ,
         \dp/ex_stage/alu/shifter/N105 , \dp/ex_stage/alu/shifter/N70 ,
         \dp/ex_stage/alu/shifter/N69 , \dp/ex_stage/alu/shifter/N68 ,
         \dp/ex_stage/alu/shifter/N67 , \dp/ex_stage/alu/shifter/N66 ,
         \dp/ex_stage/alu/shifter/N65 , \dp/ex_stage/alu/shifter/N64 ,
         \dp/ex_stage/alu/shifter/N63 , \dp/ex_stage/alu/shifter/N62 ,
         \dp/ex_stage/alu/shifter/N61 , \dp/ex_stage/alu/shifter/N60 ,
         \dp/ex_stage/alu/shifter/N59 , \dp/ex_stage/alu/shifter/N58 ,
         \dp/ex_stage/alu/shifter/N57 , \dp/ex_stage/alu/shifter/N56 ,
         \dp/ex_stage/alu/shifter/N55 , \dp/ex_stage/alu/shifter/N54 ,
         \dp/ex_stage/alu/shifter/N53 , \dp/ex_stage/alu/shifter/N52 ,
         \dp/ex_stage/alu/shifter/N51 , \dp/ex_stage/alu/shifter/N50 ,
         \dp/ex_stage/alu/shifter/N49 , \dp/ex_stage/alu/shifter/N48 ,
         \dp/ex_stage/alu/shifter/N47 , \dp/ex_stage/alu/shifter/N46 ,
         \dp/ex_stage/alu/shifter/N45 , \dp/ex_stage/alu/shifter/N44 ,
         \dp/ex_stage/alu/shifter/N43 , \dp/ex_stage/alu/shifter/N42 ,
         \dp/ex_stage/alu/shifter/N41 , \dp/ex_stage/alu/shifter/N40 ,
         \dp/ex_stage/alu/shifter/N39 , \dp/ex_stage/alu/shifter/N38 ,
         \dp/ex_stage/alu/shifter/N37 , \dp/ex_stage/alu/shifter/N36 ,
         \dp/ex_stage/alu/shifter/N35 , \dp/ex_stage/alu/shifter/N34 ,
         \dp/ex_stage/alu/shifter/N33 , \dp/ex_stage/alu/shifter/N32 ,
         \dp/ex_stage/alu/shifter/N31 , \dp/ex_stage/alu/shifter/N30 ,
         \dp/ex_stage/alu/shifter/N29 , \dp/ex_stage/alu/shifter/N28 ,
         \dp/ex_stage/alu/shifter/N27 , \dp/ex_stage/alu/shifter/N26 ,
         \dp/ex_stage/alu/shifter/N25 , \dp/ex_stage/alu/shifter/N24 ,
         \dp/ex_stage/alu/shifter/N23 , \dp/ex_stage/alu/shifter/N22 ,
         \dp/ex_stage/alu/shifter/N21 , \dp/ex_stage/alu/shifter/N20 ,
         \dp/ex_stage/alu/shifter/N19 , \dp/ex_stage/alu/shifter/N18 ,
         \dp/ex_stage/alu/shifter/N17 , \dp/ex_stage/alu/shifter/N16 ,
         \dp/ex_stage/alu/shifter/N15 , \dp/ex_stage/alu/shifter/N14 ,
         \dp/ex_stage/alu/shifter/N13 , \dp/ex_stage/alu/shifter/N12 ,
         \dp/ex_stage/alu/shifter/N11 , \dp/ex_stage/alu/shifter/N10 ,
         \dp/ex_stage/alu/shifter/N9 , \dp/ex_stage/alu/shifter/N8 ,
         \dp/ex_stage/alu/shifter/N7 , \dp/ex_stage/alu/shifter/sll_48/n29 ,
         \dp/ex_stage/alu/shifter/sll_48/n28 ,
         \dp/ex_stage/alu/shifter/sll_48/n27 ,
         \dp/ex_stage/alu/shifter/sll_48/n26 ,
         \dp/ex_stage/alu/shifter/sll_48/n25 ,
         \dp/ex_stage/alu/shifter/sll_48/n24 ,
         \dp/ex_stage/alu/shifter/sll_48/n23 ,
         \dp/ex_stage/alu/shifter/sll_48/n22 ,
         \dp/ex_stage/alu/shifter/sll_48/n21 ,
         \dp/ex_stage/alu/shifter/sll_48/n20 ,
         \dp/ex_stage/alu/shifter/sll_48/n19 ,
         \dp/ex_stage/alu/shifter/sll_48/n18 ,
         \dp/ex_stage/alu/shifter/sll_48/n17 ,
         \dp/ex_stage/alu/shifter/sll_48/n16 ,
         \dp/ex_stage/alu/shifter/sll_48/n15 ,
         \dp/ex_stage/alu/shifter/sll_48/n14 ,
         \dp/ex_stage/alu/shifter/sll_48/n13 ,
         \dp/ex_stage/alu/shifter/sll_48/n12 ,
         \dp/ex_stage/alu/shifter/sll_48/n11 ,
         \dp/ex_stage/alu/shifter/sll_48/n10 ,
         \dp/ex_stage/alu/shifter/sll_48/n9 ,
         \dp/ex_stage/alu/shifter/sll_48/n8 ,
         \dp/ex_stage/alu/shifter/sll_48/n7 ,
         \dp/ex_stage/alu/shifter/sll_48/n6 ,
         \dp/ex_stage/alu/shifter/sll_48/n5 ,
         \dp/ex_stage/alu/shifter/sll_48/n4 ,
         \dp/ex_stage/alu/shifter/sll_48/n3 ,
         \dp/ex_stage/alu/shifter/sll_48/n2 ,
         \dp/ex_stage/alu/shifter/sll_48/n1 ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][8] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][9] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][10] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][11] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][12] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][13] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][14] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][15] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][16] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][17] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][18] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][19] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][20] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][21] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][22] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][23] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][24] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][25] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][26] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][27] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][28] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][29] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][30] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[4][31] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][0] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][1] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][2] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][3] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][4] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][5] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][6] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][7] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][8] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][9] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][10] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][11] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][12] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][13] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][14] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][15] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][16] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][17] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][18] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][19] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][20] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][21] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][22] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][23] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][24] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][25] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][26] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][27] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][28] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][29] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][30] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[3][31] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][0] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][1] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][2] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][3] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][4] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][5] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][6] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][7] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][8] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][9] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][10] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][11] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][12] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][13] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][14] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][15] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][16] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][17] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][18] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][19] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][20] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][21] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][22] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][23] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][24] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][25] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][26] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][27] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][28] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][29] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][30] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[2][31] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][0] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][1] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][2] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][3] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][4] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][5] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][6] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][7] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][8] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][9] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][10] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][11] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][12] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][13] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][14] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][15] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][16] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][17] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][18] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][19] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][20] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][21] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][22] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][23] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][24] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][25] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][26] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][27] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][28] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][29] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][30] ,
         \dp/ex_stage/alu/shifter/sll_48/ML_int[1][31] ,
         \dp/ex_stage/alu/shifter/sla_46/n189 ,
         \dp/ex_stage/alu/shifter/sla_46/n188 ,
         \dp/ex_stage/alu/shifter/sla_46/n187 ,
         \dp/ex_stage/alu/shifter/sla_46/n186 ,
         \dp/ex_stage/alu/shifter/sla_46/n185 ,
         \dp/ex_stage/alu/shifter/sla_46/n184 ,
         \dp/ex_stage/alu/shifter/sla_46/n183 ,
         \dp/ex_stage/alu/shifter/sla_46/n182 ,
         \dp/ex_stage/alu/shifter/sla_46/n181 ,
         \dp/ex_stage/alu/shifter/sla_46/n180 ,
         \dp/ex_stage/alu/shifter/sla_46/n179 ,
         \dp/ex_stage/alu/shifter/sla_46/n178 ,
         \dp/ex_stage/alu/shifter/sla_46/n177 ,
         \dp/ex_stage/alu/shifter/sla_46/n176 ,
         \dp/ex_stage/alu/shifter/sla_46/n175 ,
         \dp/ex_stage/alu/shifter/sla_46/n174 ,
         \dp/ex_stage/alu/shifter/sla_46/n173 ,
         \dp/ex_stage/alu/shifter/sla_46/n172 ,
         \dp/ex_stage/alu/shifter/sla_46/n171 ,
         \dp/ex_stage/alu/shifter/sla_46/n170 ,
         \dp/ex_stage/alu/shifter/sla_46/n169 ,
         \dp/ex_stage/alu/shifter/sla_46/n168 ,
         \dp/ex_stage/alu/shifter/sla_46/n167 ,
         \dp/ex_stage/alu/shifter/sla_46/n166 ,
         \dp/ex_stage/alu/shifter/sla_46/n165 ,
         \dp/ex_stage/alu/shifter/sla_46/n164 ,
         \dp/ex_stage/alu/shifter/sla_46/n163 ,
         \dp/ex_stage/alu/shifter/sla_46/n162 ,
         \dp/ex_stage/alu/shifter/sla_46/n161 ,
         \dp/ex_stage/alu/shifter/sla_46/n160 ,
         \dp/ex_stage/alu/shifter/sla_46/n159 ,
         \dp/ex_stage/alu/shifter/sla_46/n158 ,
         \dp/ex_stage/alu/shifter/sla_46/n157 ,
         \dp/ex_stage/alu/shifter/sla_46/n156 ,
         \dp/ex_stage/alu/shifter/sla_46/n155 ,
         \dp/ex_stage/alu/shifter/sla_46/n154 ,
         \dp/ex_stage/alu/shifter/sla_46/n153 ,
         \dp/ex_stage/alu/shifter/sla_46/n152 ,
         \dp/ex_stage/alu/shifter/sla_46/n151 ,
         \dp/ex_stage/alu/shifter/sla_46/n150 ,
         \dp/ex_stage/alu/shifter/sla_46/n149 ,
         \dp/ex_stage/alu/shifter/sla_46/n148 ,
         \dp/ex_stage/alu/shifter/sla_46/n147 ,
         \dp/ex_stage/alu/shifter/sla_46/n146 ,
         \dp/ex_stage/alu/shifter/sla_46/n145 ,
         \dp/ex_stage/alu/shifter/sla_46/n144 ,
         \dp/ex_stage/alu/shifter/sla_46/n143 ,
         \dp/ex_stage/alu/shifter/sla_46/n142 ,
         \dp/ex_stage/alu/shifter/sla_46/n141 ,
         \dp/ex_stage/alu/shifter/sla_46/n140 ,
         \dp/ex_stage/alu/shifter/sla_46/n139 ,
         \dp/ex_stage/alu/shifter/sla_46/n138 ,
         \dp/ex_stage/alu/shifter/sla_46/n137 ,
         \dp/ex_stage/alu/shifter/sla_46/n136 ,
         \dp/ex_stage/alu/shifter/sla_46/n135 ,
         \dp/ex_stage/alu/shifter/sla_46/n134 ,
         \dp/ex_stage/alu/shifter/sla_46/n133 ,
         \dp/ex_stage/alu/shifter/sla_46/n132 ,
         \dp/ex_stage/alu/shifter/sla_46/n131 ,
         \dp/ex_stage/alu/shifter/sla_46/n130 ,
         \dp/ex_stage/alu/shifter/sla_46/n129 ,
         \dp/ex_stage/alu/shifter/sla_46/n128 ,
         \dp/ex_stage/alu/shifter/sla_46/n127 ,
         \dp/ex_stage/alu/shifter/sla_46/n126 ,
         \dp/ex_stage/alu/shifter/sla_46/n125 ,
         \dp/ex_stage/alu/shifter/sla_46/n124 ,
         \dp/ex_stage/alu/shifter/sla_46/n123 ,
         \dp/ex_stage/alu/shifter/sla_46/n122 ,
         \dp/ex_stage/alu/shifter/sla_46/n121 ,
         \dp/ex_stage/alu/shifter/sla_46/n120 ,
         \dp/ex_stage/alu/shifter/sla_46/n119 ,
         \dp/ex_stage/alu/shifter/sla_46/n118 ,
         \dp/ex_stage/alu/shifter/sla_46/n117 ,
         \dp/ex_stage/alu/shifter/sla_46/n116 ,
         \dp/ex_stage/alu/shifter/sla_46/n115 ,
         \dp/ex_stage/alu/shifter/sla_46/n114 ,
         \dp/ex_stage/alu/shifter/sla_46/n113 ,
         \dp/ex_stage/alu/shifter/sla_46/n112 ,
         \dp/ex_stage/alu/shifter/sla_46/n111 ,
         \dp/ex_stage/alu/shifter/sla_46/n110 ,
         \dp/ex_stage/alu/shifter/sla_46/n109 ,
         \dp/ex_stage/alu/shifter/sla_46/n108 ,
         \dp/ex_stage/alu/shifter/sla_46/n107 ,
         \dp/ex_stage/alu/shifter/sla_46/n106 ,
         \dp/ex_stage/alu/shifter/sla_46/n105 ,
         \dp/ex_stage/alu/shifter/sla_46/n104 ,
         \dp/ex_stage/alu/shifter/sla_46/n103 ,
         \dp/ex_stage/alu/shifter/sla_46/n102 ,
         \dp/ex_stage/alu/shifter/sla_46/n101 ,
         \dp/ex_stage/alu/shifter/sla_46/n100 ,
         \dp/ex_stage/alu/shifter/sla_46/n99 ,
         \dp/ex_stage/alu/shifter/sla_46/n98 ,
         \dp/ex_stage/alu/shifter/sla_46/n97 ,
         \dp/ex_stage/alu/shifter/sla_46/n96 ,
         \dp/ex_stage/alu/shifter/sla_46/n95 ,
         \dp/ex_stage/alu/shifter/sla_46/n94 ,
         \dp/ex_stage/alu/shifter/sla_46/n93 ,
         \dp/ex_stage/alu/shifter/sla_46/n92 ,
         \dp/ex_stage/alu/shifter/sla_46/n91 ,
         \dp/ex_stage/alu/shifter/sla_46/n90 ,
         \dp/ex_stage/alu/shifter/sla_46/n89 ,
         \dp/ex_stage/alu/shifter/sla_46/n88 ,
         \dp/ex_stage/alu/shifter/sla_46/n87 ,
         \dp/ex_stage/alu/shifter/sla_46/n86 ,
         \dp/ex_stage/alu/shifter/sla_46/n85 ,
         \dp/ex_stage/alu/shifter/sla_46/n84 ,
         \dp/ex_stage/alu/shifter/sla_46/n83 ,
         \dp/ex_stage/alu/shifter/sla_46/n82 ,
         \dp/ex_stage/alu/shifter/sla_46/n81 ,
         \dp/ex_stage/alu/shifter/sla_46/n80 ,
         \dp/ex_stage/alu/shifter/sla_46/n79 ,
         \dp/ex_stage/alu/shifter/sla_46/n78 ,
         \dp/ex_stage/alu/shifter/sla_46/n77 ,
         \dp/ex_stage/alu/shifter/sla_46/n76 ,
         \dp/ex_stage/alu/shifter/sla_46/n75 ,
         \dp/ex_stage/alu/shifter/sla_46/n74 ,
         \dp/ex_stage/alu/shifter/sla_46/n73 ,
         \dp/ex_stage/alu/shifter/sla_46/n72 ,
         \dp/ex_stage/alu/shifter/sla_46/n71 ,
         \dp/ex_stage/alu/shifter/sla_46/n70 ,
         \dp/ex_stage/alu/shifter/sla_46/n69 ,
         \dp/ex_stage/alu/shifter/sla_46/n68 ,
         \dp/ex_stage/alu/shifter/sla_46/n67 ,
         \dp/ex_stage/alu/shifter/sla_46/n66 ,
         \dp/ex_stage/alu/shifter/sla_46/n65 ,
         \dp/ex_stage/alu/shifter/sla_46/n64 ,
         \dp/ex_stage/alu/shifter/sla_46/n63 ,
         \dp/ex_stage/alu/shifter/sla_46/n62 ,
         \dp/ex_stage/alu/shifter/sla_46/n61 ,
         \dp/ex_stage/alu/shifter/sla_46/n60 ,
         \dp/ex_stage/alu/shifter/sla_46/n59 ,
         \dp/ex_stage/alu/shifter/sla_46/n58 ,
         \dp/ex_stage/alu/shifter/sla_46/n57 ,
         \dp/ex_stage/alu/shifter/sla_46/n56 ,
         \dp/ex_stage/alu/shifter/sla_46/n55 ,
         \dp/ex_stage/alu/shifter/sla_46/n54 ,
         \dp/ex_stage/alu/shifter/sla_46/n53 ,
         \dp/ex_stage/alu/shifter/sla_46/n52 ,
         \dp/ex_stage/alu/shifter/sla_46/n51 ,
         \dp/ex_stage/alu/shifter/sla_46/n50 ,
         \dp/ex_stage/alu/shifter/sla_46/n49 ,
         \dp/ex_stage/alu/shifter/sla_46/n48 ,
         \dp/ex_stage/alu/shifter/sla_46/n47 ,
         \dp/ex_stage/alu/shifter/sla_46/n46 ,
         \dp/ex_stage/alu/shifter/sla_46/n45 ,
         \dp/ex_stage/alu/shifter/sla_46/n44 ,
         \dp/ex_stage/alu/shifter/sla_46/n43 ,
         \dp/ex_stage/alu/shifter/sla_46/n42 ,
         \dp/ex_stage/alu/shifter/sla_46/n41 ,
         \dp/ex_stage/alu/shifter/sla_46/n40 ,
         \dp/ex_stage/alu/shifter/sla_46/n39 ,
         \dp/ex_stage/alu/shifter/sla_46/n38 ,
         \dp/ex_stage/alu/shifter/sla_46/n37 ,
         \dp/ex_stage/alu/shifter/sla_46/n36 ,
         \dp/ex_stage/alu/shifter/sla_46/n35 ,
         \dp/ex_stage/alu/shifter/sla_46/n34 ,
         \dp/ex_stage/alu/shifter/sla_46/n33 ,
         \dp/ex_stage/alu/shifter/sla_46/n32 ,
         \dp/ex_stage/alu/shifter/sla_46/n31 ,
         \dp/ex_stage/alu/shifter/sla_46/n30 ,
         \dp/ex_stage/alu/shifter/sla_46/n29 ,
         \dp/ex_stage/alu/shifter/sla_46/n28 ,
         \dp/ex_stage/alu/shifter/sla_46/n27 ,
         \dp/ex_stage/alu/shifter/sla_46/n26 ,
         \dp/ex_stage/alu/shifter/sla_46/n25 ,
         \dp/ex_stage/alu/shifter/sla_46/n24 ,
         \dp/ex_stage/alu/shifter/sla_46/n23 ,
         \dp/ex_stage/alu/shifter/sla_46/n22 ,
         \dp/ex_stage/alu/shifter/sla_46/n21 ,
         \dp/ex_stage/alu/shifter/sla_46/n20 ,
         \dp/ex_stage/alu/shifter/sla_46/n19 ,
         \dp/ex_stage/alu/shifter/sla_46/n18 ,
         \dp/ex_stage/alu/shifter/sla_46/n17 ,
         \dp/ex_stage/alu/shifter/sla_46/n16 ,
         \dp/ex_stage/alu/shifter/sla_46/n15 ,
         \dp/ex_stage/alu/shifter/sla_46/n14 ,
         \dp/ex_stage/alu/shifter/sla_46/n13 ,
         \dp/ex_stage/alu/shifter/sla_46/n12 ,
         \dp/ex_stage/alu/shifter/sla_46/n11 ,
         \dp/ex_stage/alu/shifter/sla_46/n10 ,
         \dp/ex_stage/alu/shifter/sla_46/n9 ,
         \dp/ex_stage/alu/shifter/sla_46/n8 ,
         \dp/ex_stage/alu/shifter/sla_46/n7 ,
         \dp/ex_stage/alu/shifter/sla_46/n6 ,
         \dp/ex_stage/alu/shifter/sla_46/n5 ,
         \dp/ex_stage/alu/shifter/sla_46/n4 ,
         \dp/ex_stage/alu/shifter/sla_46/n3 ,
         \dp/ex_stage/alu/shifter/sla_46/n2 ,
         \dp/ex_stage/alu/shifter/sla_46/n1 ,
         \dp/ex_stage/alu/shifter/srl_41/n167 ,
         \dp/ex_stage/alu/shifter/srl_41/n166 ,
         \dp/ex_stage/alu/shifter/srl_41/n165 ,
         \dp/ex_stage/alu/shifter/srl_41/n164 ,
         \dp/ex_stage/alu/shifter/srl_41/n163 ,
         \dp/ex_stage/alu/shifter/srl_41/n162 ,
         \dp/ex_stage/alu/shifter/srl_41/n161 ,
         \dp/ex_stage/alu/shifter/srl_41/n160 ,
         \dp/ex_stage/alu/shifter/srl_41/n159 ,
         \dp/ex_stage/alu/shifter/srl_41/n158 ,
         \dp/ex_stage/alu/shifter/srl_41/n157 ,
         \dp/ex_stage/alu/shifter/srl_41/n156 ,
         \dp/ex_stage/alu/shifter/srl_41/n155 ,
         \dp/ex_stage/alu/shifter/srl_41/n154 ,
         \dp/ex_stage/alu/shifter/srl_41/n153 ,
         \dp/ex_stage/alu/shifter/srl_41/n152 ,
         \dp/ex_stage/alu/shifter/srl_41/n151 ,
         \dp/ex_stage/alu/shifter/srl_41/n150 ,
         \dp/ex_stage/alu/shifter/srl_41/n149 ,
         \dp/ex_stage/alu/shifter/srl_41/n148 ,
         \dp/ex_stage/alu/shifter/srl_41/n147 ,
         \dp/ex_stage/alu/shifter/srl_41/n146 ,
         \dp/ex_stage/alu/shifter/srl_41/n145 ,
         \dp/ex_stage/alu/shifter/srl_41/n144 ,
         \dp/ex_stage/alu/shifter/srl_41/n143 ,
         \dp/ex_stage/alu/shifter/srl_41/n142 ,
         \dp/ex_stage/alu/shifter/srl_41/n141 ,
         \dp/ex_stage/alu/shifter/srl_41/n140 ,
         \dp/ex_stage/alu/shifter/srl_41/n139 ,
         \dp/ex_stage/alu/shifter/srl_41/n138 ,
         \dp/ex_stage/alu/shifter/srl_41/n137 ,
         \dp/ex_stage/alu/shifter/srl_41/n136 ,
         \dp/ex_stage/alu/shifter/srl_41/n135 ,
         \dp/ex_stage/alu/shifter/srl_41/n134 ,
         \dp/ex_stage/alu/shifter/srl_41/n133 ,
         \dp/ex_stage/alu/shifter/srl_41/n132 ,
         \dp/ex_stage/alu/shifter/srl_41/n131 ,
         \dp/ex_stage/alu/shifter/srl_41/n130 ,
         \dp/ex_stage/alu/shifter/srl_41/n129 ,
         \dp/ex_stage/alu/shifter/srl_41/n128 ,
         \dp/ex_stage/alu/shifter/srl_41/n127 ,
         \dp/ex_stage/alu/shifter/srl_41/n126 ,
         \dp/ex_stage/alu/shifter/srl_41/n125 ,
         \dp/ex_stage/alu/shifter/srl_41/n124 ,
         \dp/ex_stage/alu/shifter/srl_41/n123 ,
         \dp/ex_stage/alu/shifter/srl_41/n122 ,
         \dp/ex_stage/alu/shifter/srl_41/n121 ,
         \dp/ex_stage/alu/shifter/srl_41/n120 ,
         \dp/ex_stage/alu/shifter/srl_41/n119 ,
         \dp/ex_stage/alu/shifter/srl_41/n118 ,
         \dp/ex_stage/alu/shifter/srl_41/n117 ,
         \dp/ex_stage/alu/shifter/srl_41/n116 ,
         \dp/ex_stage/alu/shifter/srl_41/n115 ,
         \dp/ex_stage/alu/shifter/srl_41/n114 ,
         \dp/ex_stage/alu/shifter/srl_41/n113 ,
         \dp/ex_stage/alu/shifter/srl_41/n112 ,
         \dp/ex_stage/alu/shifter/srl_41/n111 ,
         \dp/ex_stage/alu/shifter/srl_41/n110 ,
         \dp/ex_stage/alu/shifter/srl_41/n109 ,
         \dp/ex_stage/alu/shifter/srl_41/n108 ,
         \dp/ex_stage/alu/shifter/srl_41/n107 ,
         \dp/ex_stage/alu/shifter/srl_41/n106 ,
         \dp/ex_stage/alu/shifter/srl_41/n105 ,
         \dp/ex_stage/alu/shifter/srl_41/n104 ,
         \dp/ex_stage/alu/shifter/srl_41/n103 ,
         \dp/ex_stage/alu/shifter/srl_41/n102 ,
         \dp/ex_stage/alu/shifter/srl_41/n101 ,
         \dp/ex_stage/alu/shifter/srl_41/n100 ,
         \dp/ex_stage/alu/shifter/srl_41/n99 ,
         \dp/ex_stage/alu/shifter/srl_41/n98 ,
         \dp/ex_stage/alu/shifter/srl_41/n97 ,
         \dp/ex_stage/alu/shifter/srl_41/n96 ,
         \dp/ex_stage/alu/shifter/srl_41/n95 ,
         \dp/ex_stage/alu/shifter/srl_41/n94 ,
         \dp/ex_stage/alu/shifter/srl_41/n93 ,
         \dp/ex_stage/alu/shifter/srl_41/n92 ,
         \dp/ex_stage/alu/shifter/srl_41/n91 ,
         \dp/ex_stage/alu/shifter/srl_41/n90 ,
         \dp/ex_stage/alu/shifter/srl_41/n89 ,
         \dp/ex_stage/alu/shifter/srl_41/n88 ,
         \dp/ex_stage/alu/shifter/srl_41/n87 ,
         \dp/ex_stage/alu/shifter/srl_41/n86 ,
         \dp/ex_stage/alu/shifter/srl_41/n85 ,
         \dp/ex_stage/alu/shifter/srl_41/n84 ,
         \dp/ex_stage/alu/shifter/srl_41/n83 ,
         \dp/ex_stage/alu/shifter/srl_41/n82 ,
         \dp/ex_stage/alu/shifter/srl_41/n81 ,
         \dp/ex_stage/alu/shifter/srl_41/n80 ,
         \dp/ex_stage/alu/shifter/srl_41/n79 ,
         \dp/ex_stage/alu/shifter/srl_41/n78 ,
         \dp/ex_stage/alu/shifter/srl_41/n77 ,
         \dp/ex_stage/alu/shifter/srl_41/n76 ,
         \dp/ex_stage/alu/shifter/srl_41/n75 ,
         \dp/ex_stage/alu/shifter/srl_41/n74 ,
         \dp/ex_stage/alu/shifter/srl_41/n73 ,
         \dp/ex_stage/alu/shifter/srl_41/n72 ,
         \dp/ex_stage/alu/shifter/srl_41/n71 ,
         \dp/ex_stage/alu/shifter/srl_41/n70 ,
         \dp/ex_stage/alu/shifter/srl_41/n69 ,
         \dp/ex_stage/alu/shifter/srl_41/n68 ,
         \dp/ex_stage/alu/shifter/srl_41/n67 ,
         \dp/ex_stage/alu/shifter/srl_41/n66 ,
         \dp/ex_stage/alu/shifter/srl_41/n65 ,
         \dp/ex_stage/alu/shifter/srl_41/n64 ,
         \dp/ex_stage/alu/shifter/srl_41/n63 ,
         \dp/ex_stage/alu/shifter/srl_41/n62 ,
         \dp/ex_stage/alu/shifter/srl_41/n61 ,
         \dp/ex_stage/alu/shifter/srl_41/n60 ,
         \dp/ex_stage/alu/shifter/srl_41/n59 ,
         \dp/ex_stage/alu/shifter/srl_41/n58 ,
         \dp/ex_stage/alu/shifter/srl_41/n57 ,
         \dp/ex_stage/alu/shifter/srl_41/n56 ,
         \dp/ex_stage/alu/shifter/srl_41/n55 ,
         \dp/ex_stage/alu/shifter/srl_41/n54 ,
         \dp/ex_stage/alu/shifter/srl_41/n53 ,
         \dp/ex_stage/alu/shifter/srl_41/n52 ,
         \dp/ex_stage/alu/shifter/srl_41/n51 ,
         \dp/ex_stage/alu/shifter/srl_41/n50 ,
         \dp/ex_stage/alu/shifter/srl_41/n49 ,
         \dp/ex_stage/alu/shifter/srl_41/n48 ,
         \dp/ex_stage/alu/shifter/srl_41/n47 ,
         \dp/ex_stage/alu/shifter/srl_41/n46 ,
         \dp/ex_stage/alu/shifter/srl_41/n45 ,
         \dp/ex_stage/alu/shifter/srl_41/n44 ,
         \dp/ex_stage/alu/shifter/srl_41/n43 ,
         \dp/ex_stage/alu/shifter/srl_41/n42 ,
         \dp/ex_stage/alu/shifter/srl_41/n41 ,
         \dp/ex_stage/alu/shifter/srl_41/n40 ,
         \dp/ex_stage/alu/shifter/srl_41/n39 ,
         \dp/ex_stage/alu/shifter/srl_41/n38 ,
         \dp/ex_stage/alu/shifter/srl_41/n37 ,
         \dp/ex_stage/alu/shifter/srl_41/n36 ,
         \dp/ex_stage/alu/shifter/srl_41/n35 ,
         \dp/ex_stage/alu/shifter/srl_41/n34 ,
         \dp/ex_stage/alu/shifter/srl_41/n33 ,
         \dp/ex_stage/alu/shifter/srl_41/n32 ,
         \dp/ex_stage/alu/shifter/srl_41/n31 ,
         \dp/ex_stage/alu/shifter/srl_41/n29 ,
         \dp/ex_stage/alu/shifter/srl_41/n28 ,
         \dp/ex_stage/alu/shifter/srl_41/n27 ,
         \dp/ex_stage/alu/shifter/srl_41/n26 ,
         \dp/ex_stage/alu/shifter/srl_41/n25 ,
         \dp/ex_stage/alu/shifter/srl_41/n24 ,
         \dp/ex_stage/alu/shifter/srl_41/n23 ,
         \dp/ex_stage/alu/shifter/srl_41/n22 ,
         \dp/ex_stage/alu/shifter/srl_41/n21 ,
         \dp/ex_stage/alu/shifter/srl_41/n20 ,
         \dp/ex_stage/alu/shifter/srl_41/n19 ,
         \dp/ex_stage/alu/shifter/srl_41/n18 ,
         \dp/ex_stage/alu/shifter/srl_41/n17 ,
         \dp/ex_stage/alu/shifter/srl_41/n16 ,
         \dp/ex_stage/alu/shifter/srl_41/n15 ,
         \dp/ex_stage/alu/shifter/srl_41/n14 ,
         \dp/ex_stage/alu/shifter/srl_41/n13 ,
         \dp/ex_stage/alu/shifter/srl_41/n12 ,
         \dp/ex_stage/alu/shifter/srl_41/n11 ,
         \dp/ex_stage/alu/shifter/srl_41/n10 ,
         \dp/ex_stage/alu/shifter/srl_41/n9 ,
         \dp/ex_stage/alu/shifter/srl_41/n8 ,
         \dp/ex_stage/alu/shifter/srl_41/n7 ,
         \dp/ex_stage/alu/shifter/srl_41/n6 ,
         \dp/ex_stage/alu/shifter/srl_41/n5 ,
         \dp/ex_stage/alu/shifter/srl_41/n4 ,
         \dp/ex_stage/alu/shifter/srl_41/n3 ,
         \dp/ex_stage/alu/shifter/srl_41/n2 ,
         \dp/ex_stage/alu/shifter/srl_41/n1 ,
         \dp/ex_stage/alu/shifter/sra_39/n174 ,
         \dp/ex_stage/alu/shifter/sra_39/n173 ,
         \dp/ex_stage/alu/shifter/sra_39/n172 ,
         \dp/ex_stage/alu/shifter/sra_39/n171 ,
         \dp/ex_stage/alu/shifter/sra_39/n170 ,
         \dp/ex_stage/alu/shifter/sra_39/n169 ,
         \dp/ex_stage/alu/shifter/sra_39/n168 ,
         \dp/ex_stage/alu/shifter/sra_39/n167 ,
         \dp/ex_stage/alu/shifter/sra_39/n166 ,
         \dp/ex_stage/alu/shifter/sra_39/n165 ,
         \dp/ex_stage/alu/shifter/sra_39/n164 ,
         \dp/ex_stage/alu/shifter/sra_39/n163 ,
         \dp/ex_stage/alu/shifter/sra_39/n162 ,
         \dp/ex_stage/alu/shifter/sra_39/n161 ,
         \dp/ex_stage/alu/shifter/sra_39/n160 ,
         \dp/ex_stage/alu/shifter/sra_39/n159 ,
         \dp/ex_stage/alu/shifter/sra_39/n158 ,
         \dp/ex_stage/alu/shifter/sra_39/n157 ,
         \dp/ex_stage/alu/shifter/sra_39/n156 ,
         \dp/ex_stage/alu/shifter/sra_39/n155 ,
         \dp/ex_stage/alu/shifter/sra_39/n154 ,
         \dp/ex_stage/alu/shifter/sra_39/n153 ,
         \dp/ex_stage/alu/shifter/sra_39/n152 ,
         \dp/ex_stage/alu/shifter/sra_39/n151 ,
         \dp/ex_stage/alu/shifter/sra_39/n150 ,
         \dp/ex_stage/alu/shifter/sra_39/n149 ,
         \dp/ex_stage/alu/shifter/sra_39/n148 ,
         \dp/ex_stage/alu/shifter/sra_39/n147 ,
         \dp/ex_stage/alu/shifter/sra_39/n146 ,
         \dp/ex_stage/alu/shifter/sra_39/n145 ,
         \dp/ex_stage/alu/shifter/sra_39/n144 ,
         \dp/ex_stage/alu/shifter/sra_39/n143 ,
         \dp/ex_stage/alu/shifter/sra_39/n142 ,
         \dp/ex_stage/alu/shifter/sra_39/n141 ,
         \dp/ex_stage/alu/shifter/sra_39/n140 ,
         \dp/ex_stage/alu/shifter/sra_39/n139 ,
         \dp/ex_stage/alu/shifter/sra_39/n138 ,
         \dp/ex_stage/alu/shifter/sra_39/n137 ,
         \dp/ex_stage/alu/shifter/sra_39/n136 ,
         \dp/ex_stage/alu/shifter/sra_39/n135 ,
         \dp/ex_stage/alu/shifter/sra_39/n134 ,
         \dp/ex_stage/alu/shifter/sra_39/n133 ,
         \dp/ex_stage/alu/shifter/sra_39/n132 ,
         \dp/ex_stage/alu/shifter/sra_39/n131 ,
         \dp/ex_stage/alu/shifter/sra_39/n130 ,
         \dp/ex_stage/alu/shifter/sra_39/n129 ,
         \dp/ex_stage/alu/shifter/sra_39/n128 ,
         \dp/ex_stage/alu/shifter/sra_39/n127 ,
         \dp/ex_stage/alu/shifter/sra_39/n126 ,
         \dp/ex_stage/alu/shifter/sra_39/n125 ,
         \dp/ex_stage/alu/shifter/sra_39/n124 ,
         \dp/ex_stage/alu/shifter/sra_39/n123 ,
         \dp/ex_stage/alu/shifter/sra_39/n122 ,
         \dp/ex_stage/alu/shifter/sra_39/n121 ,
         \dp/ex_stage/alu/shifter/sra_39/n120 ,
         \dp/ex_stage/alu/shifter/sra_39/n119 ,
         \dp/ex_stage/alu/shifter/sra_39/n118 ,
         \dp/ex_stage/alu/shifter/sra_39/n117 ,
         \dp/ex_stage/alu/shifter/sra_39/n116 ,
         \dp/ex_stage/alu/shifter/sra_39/n115 ,
         \dp/ex_stage/alu/shifter/sra_39/n114 ,
         \dp/ex_stage/alu/shifter/sra_39/n113 ,
         \dp/ex_stage/alu/shifter/sra_39/n112 ,
         \dp/ex_stage/alu/shifter/sra_39/n111 ,
         \dp/ex_stage/alu/shifter/sra_39/n110 ,
         \dp/ex_stage/alu/shifter/sra_39/n109 ,
         \dp/ex_stage/alu/shifter/sra_39/n108 ,
         \dp/ex_stage/alu/shifter/sra_39/n107 ,
         \dp/ex_stage/alu/shifter/sra_39/n106 ,
         \dp/ex_stage/alu/shifter/sra_39/n105 ,
         \dp/ex_stage/alu/shifter/sra_39/n104 ,
         \dp/ex_stage/alu/shifter/sra_39/n103 ,
         \dp/ex_stage/alu/shifter/sra_39/n102 ,
         \dp/ex_stage/alu/shifter/sra_39/n101 ,
         \dp/ex_stage/alu/shifter/sra_39/n100 ,
         \dp/ex_stage/alu/shifter/sra_39/n99 ,
         \dp/ex_stage/alu/shifter/sra_39/n98 ,
         \dp/ex_stage/alu/shifter/sra_39/n97 ,
         \dp/ex_stage/alu/shifter/sra_39/n96 ,
         \dp/ex_stage/alu/shifter/sra_39/n95 ,
         \dp/ex_stage/alu/shifter/sra_39/n94 ,
         \dp/ex_stage/alu/shifter/sra_39/n93 ,
         \dp/ex_stage/alu/shifter/sra_39/n92 ,
         \dp/ex_stage/alu/shifter/sra_39/n91 ,
         \dp/ex_stage/alu/shifter/sra_39/n90 ,
         \dp/ex_stage/alu/shifter/sra_39/n89 ,
         \dp/ex_stage/alu/shifter/sra_39/n88 ,
         \dp/ex_stage/alu/shifter/sra_39/n87 ,
         \dp/ex_stage/alu/shifter/sra_39/n86 ,
         \dp/ex_stage/alu/shifter/sra_39/n85 ,
         \dp/ex_stage/alu/shifter/sra_39/n84 ,
         \dp/ex_stage/alu/shifter/sra_39/n83 ,
         \dp/ex_stage/alu/shifter/sra_39/n82 ,
         \dp/ex_stage/alu/shifter/sra_39/n81 ,
         \dp/ex_stage/alu/shifter/sra_39/n80 ,
         \dp/ex_stage/alu/shifter/sra_39/n79 ,
         \dp/ex_stage/alu/shifter/sra_39/n78 ,
         \dp/ex_stage/alu/shifter/sra_39/n77 ,
         \dp/ex_stage/alu/shifter/sra_39/n76 ,
         \dp/ex_stage/alu/shifter/sra_39/n75 ,
         \dp/ex_stage/alu/shifter/sra_39/n74 ,
         \dp/ex_stage/alu/shifter/sra_39/n73 ,
         \dp/ex_stage/alu/shifter/sra_39/n72 ,
         \dp/ex_stage/alu/shifter/sra_39/n71 ,
         \dp/ex_stage/alu/shifter/sra_39/n70 ,
         \dp/ex_stage/alu/shifter/sra_39/n69 ,
         \dp/ex_stage/alu/shifter/sra_39/n68 ,
         \dp/ex_stage/alu/shifter/sra_39/n67 ,
         \dp/ex_stage/alu/shifter/sra_39/n66 ,
         \dp/ex_stage/alu/shifter/sra_39/n65 ,
         \dp/ex_stage/alu/shifter/sra_39/n64 ,
         \dp/ex_stage/alu/shifter/sra_39/n63 ,
         \dp/ex_stage/alu/shifter/sra_39/n62 ,
         \dp/ex_stage/alu/shifter/sra_39/n61 ,
         \dp/ex_stage/alu/shifter/sra_39/n60 ,
         \dp/ex_stage/alu/shifter/sra_39/n59 ,
         \dp/ex_stage/alu/shifter/sra_39/n58 ,
         \dp/ex_stage/alu/shifter/sra_39/n57 ,
         \dp/ex_stage/alu/shifter/sra_39/n56 ,
         \dp/ex_stage/alu/shifter/sra_39/n55 ,
         \dp/ex_stage/alu/shifter/sra_39/n54 ,
         \dp/ex_stage/alu/shifter/sra_39/n53 ,
         \dp/ex_stage/alu/shifter/sra_39/n52 ,
         \dp/ex_stage/alu/shifter/sra_39/n51 ,
         \dp/ex_stage/alu/shifter/sra_39/n50 ,
         \dp/ex_stage/alu/shifter/sra_39/n49 ,
         \dp/ex_stage/alu/shifter/sra_39/n48 ,
         \dp/ex_stage/alu/shifter/sra_39/n47 ,
         \dp/ex_stage/alu/shifter/sra_39/n46 ,
         \dp/ex_stage/alu/shifter/sra_39/n45 ,
         \dp/ex_stage/alu/shifter/sra_39/n44 ,
         \dp/ex_stage/alu/shifter/sra_39/n43 ,
         \dp/ex_stage/alu/shifter/sra_39/n42 ,
         \dp/ex_stage/alu/shifter/sra_39/n41 ,
         \dp/ex_stage/alu/shifter/sra_39/n40 ,
         \dp/ex_stage/alu/shifter/sra_39/n39 ,
         \dp/ex_stage/alu/shifter/sra_39/n38 ,
         \dp/ex_stage/alu/shifter/sra_39/n37 ,
         \dp/ex_stage/alu/shifter/sra_39/n36 ,
         \dp/ex_stage/alu/shifter/sra_39/n35 ,
         \dp/ex_stage/alu/shifter/sra_39/n34 ,
         \dp/ex_stage/alu/shifter/sra_39/n33 ,
         \dp/ex_stage/alu/shifter/sra_39/n32 ,
         \dp/ex_stage/alu/shifter/sra_39/n31 ,
         \dp/ex_stage/alu/shifter/sra_39/n30 ,
         \dp/ex_stage/alu/shifter/sra_39/n29 ,
         \dp/ex_stage/alu/shifter/sra_39/n28 ,
         \dp/ex_stage/alu/shifter/sra_39/n27 ,
         \dp/ex_stage/alu/shifter/sra_39/n26 ,
         \dp/ex_stage/alu/shifter/sra_39/n25 ,
         \dp/ex_stage/alu/shifter/sra_39/n24 ,
         \dp/ex_stage/alu/shifter/sra_39/n23 ,
         \dp/ex_stage/alu/shifter/sra_39/n22 ,
         \dp/ex_stage/alu/shifter/sra_39/n21 ,
         \dp/ex_stage/alu/shifter/sra_39/n20 ,
         \dp/ex_stage/alu/shifter/sra_39/n19 ,
         \dp/ex_stage/alu/shifter/sra_39/n18 ,
         \dp/ex_stage/alu/shifter/sra_39/n17 ,
         \dp/ex_stage/alu/shifter/sra_39/n16 ,
         \dp/ex_stage/alu/shifter/sra_39/n15 ,
         \dp/ex_stage/alu/shifter/sra_39/n14 ,
         \dp/ex_stage/alu/shifter/sra_39/n13 ,
         \dp/ex_stage/alu/shifter/sra_39/n12 ,
         \dp/ex_stage/alu/shifter/sra_39/n11 ,
         \dp/ex_stage/alu/shifter/sra_39/n10 ,
         \dp/ex_stage/alu/shifter/sra_39/n9 ,
         \dp/ex_stage/alu/shifter/sra_39/n8 ,
         \dp/ex_stage/alu/shifter/sra_39/n7 ,
         \dp/ex_stage/alu/shifter/sra_39/n6 ,
         \dp/ex_stage/alu/shifter/sra_39/n5 ,
         \dp/ex_stage/alu/shifter/sra_39/n4 ,
         \dp/ex_stage/alu/shifter/sra_39/n3 ,
         \dp/ex_stage/alu/shifter/sra_39/n2 ,
         \dp/ex_stage/alu/shifter/sra_39/n1 ,
         \dp/ex_stage/alu/shifter/rol_32/n15 ,
         \dp/ex_stage/alu/shifter/rol_32/n14 ,
         \dp/ex_stage/alu/shifter/rol_32/n13 ,
         \dp/ex_stage/alu/shifter/rol_32/n12 ,
         \dp/ex_stage/alu/shifter/rol_32/n11 ,
         \dp/ex_stage/alu/shifter/rol_32/n10 ,
         \dp/ex_stage/alu/shifter/rol_32/n9 ,
         \dp/ex_stage/alu/shifter/rol_32/n8 ,
         \dp/ex_stage/alu/shifter/rol_32/n7 ,
         \dp/ex_stage/alu/shifter/rol_32/n6 ,
         \dp/ex_stage/alu/shifter/rol_32/n5 ,
         \dp/ex_stage/alu/shifter/rol_32/n4 ,
         \dp/ex_stage/alu/shifter/rol_32/n3 ,
         \dp/ex_stage/alu/shifter/rol_32/n2 ,
         \dp/ex_stage/alu/shifter/rol_32/n1 ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][0] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][1] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][2] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][3] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][4] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][5] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][6] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][7] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][8] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][9] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][10] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][11] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][12] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][13] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][14] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][15] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][16] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][17] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][18] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][19] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][20] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][21] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][22] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][23] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][24] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][25] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][26] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][27] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][28] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][29] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][30] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[4][31] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][0] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][1] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][2] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][3] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][4] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][5] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][6] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][7] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][8] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][9] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][10] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][11] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][12] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][13] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][14] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][15] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][16] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][17] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][18] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][19] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][20] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][21] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][22] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][23] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][24] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][25] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][26] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][27] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][28] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][29] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][30] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[3][31] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][0] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][1] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][2] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][3] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][4] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][5] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][6] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][7] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][8] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][9] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][10] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][11] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][12] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][13] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][14] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][15] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][16] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][17] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][18] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][19] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][20] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][21] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][22] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][23] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][24] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][25] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][26] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][27] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][28] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][29] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][30] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[2][31] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][0] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][1] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][2] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][3] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][4] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][5] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][6] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][7] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][8] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][9] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][10] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][11] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][12] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][13] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][14] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][15] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][16] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][17] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][18] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][19] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][20] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][21] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][22] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][23] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][24] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][25] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][26] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][27] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][28] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][29] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][30] ,
         \dp/ex_stage/alu/shifter/rol_32/ML_int[1][31] ,
         \dp/ex_stage/alu/shifter/ror_30/n15 ,
         \dp/ex_stage/alu/shifter/ror_30/n14 ,
         \dp/ex_stage/alu/shifter/ror_30/n13 ,
         \dp/ex_stage/alu/shifter/ror_30/n12 ,
         \dp/ex_stage/alu/shifter/ror_30/n11 ,
         \dp/ex_stage/alu/shifter/ror_30/n10 ,
         \dp/ex_stage/alu/shifter/ror_30/n9 ,
         \dp/ex_stage/alu/shifter/ror_30/n8 ,
         \dp/ex_stage/alu/shifter/ror_30/n7 ,
         \dp/ex_stage/alu/shifter/ror_30/n6 ,
         \dp/ex_stage/alu/shifter/ror_30/n5 ,
         \dp/ex_stage/alu/shifter/ror_30/n4 ,
         \dp/ex_stage/alu/shifter/ror_30/n3 ,
         \dp/ex_stage/alu/shifter/ror_30/n2 ,
         \dp/ex_stage/alu/shifter/ror_30/n1 ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][0] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][1] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][2] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][3] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][4] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][5] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][6] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][7] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][8] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][9] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][10] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][11] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][12] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][13] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][14] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][15] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][16] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][17] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][18] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][19] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][20] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][21] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][22] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][23] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][24] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][25] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][26] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][27] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][28] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][29] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][30] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[4][31] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][0] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][1] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][2] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][3] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][4] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][5] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][6] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][7] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][8] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][9] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][10] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][11] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][12] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][13] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][14] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][15] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][16] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][17] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][18] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][19] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][20] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][21] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][22] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][23] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][24] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][25] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][26] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][27] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][28] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][29] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][30] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[3][31] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][0] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][1] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][2] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][3] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][4] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][5] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][6] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][7] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][8] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][9] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][10] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][11] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][12] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][13] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][14] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][15] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][16] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][17] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][18] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][19] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][20] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][21] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][22] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][23] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][24] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][25] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][26] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][27] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][28] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][29] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][30] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[2][31] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][0] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][1] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][2] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][3] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][4] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][5] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][6] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][7] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][8] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][9] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][10] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][11] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][12] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][13] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][14] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][15] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][16] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][17] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][18] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][19] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][20] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][21] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][22] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][23] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][24] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][25] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][26] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][27] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][28] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][29] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][30] ,
         \dp/ex_stage/alu/shifter/ror_30/MR_int[1][31] ,
         \dp/ex_stage/alu/r61/n110 , \dp/ex_stage/alu/r61/n109 ,
         \dp/ex_stage/alu/r61/n108 , \dp/ex_stage/alu/r61/n107 ,
         \dp/ex_stage/alu/r61/n106 , \dp/ex_stage/alu/r61/n105 ,
         \dp/ex_stage/alu/r61/n104 , \dp/ex_stage/alu/r61/n103 ,
         \dp/ex_stage/alu/r61/n102 , \dp/ex_stage/alu/r61/n101 ,
         \dp/ex_stage/alu/r61/n100 , \dp/ex_stage/alu/r61/n99 ,
         \dp/ex_stage/alu/r61/n98 , \dp/ex_stage/alu/r61/n97 ,
         \dp/ex_stage/alu/r61/n96 , \dp/ex_stage/alu/r61/n95 ,
         \dp/ex_stage/alu/r61/n94 , \dp/ex_stage/alu/r61/n93 ,
         \dp/ex_stage/alu/r61/n92 , \dp/ex_stage/alu/r61/n91 ,
         \dp/ex_stage/alu/r61/n90 , \dp/ex_stage/alu/r61/n89 ,
         \dp/ex_stage/alu/r61/n88 , \dp/ex_stage/alu/r61/n87 ,
         \dp/ex_stage/alu/r61/n86 , \dp/ex_stage/alu/r61/n85 ,
         \dp/ex_stage/alu/r61/n84 , \dp/ex_stage/alu/r61/n83 ,
         \dp/ex_stage/alu/r61/n82 , \dp/ex_stage/alu/r61/n81 ,
         \dp/ex_stage/alu/r61/n80 , \dp/ex_stage/alu/r61/n79 ,
         \dp/ex_stage/alu/r61/n78 , \dp/ex_stage/alu/r61/n77 ,
         \dp/ex_stage/alu/r61/n76 , \dp/ex_stage/alu/r61/n75 ,
         \dp/ex_stage/alu/r61/n74 , \dp/ex_stage/alu/r61/n73 ,
         \dp/ex_stage/alu/r61/n72 , \dp/ex_stage/alu/r61/n71 ,
         \dp/ex_stage/alu/r61/n70 , \dp/ex_stage/alu/r61/n69 ,
         \dp/ex_stage/alu/r61/n68 , \dp/ex_stage/alu/r61/n67 ,
         \dp/ex_stage/alu/r61/n66 , \dp/ex_stage/alu/r61/n65 ,
         \dp/ex_stage/alu/r61/n64 , \dp/ex_stage/alu/r61/n63 ,
         \dp/ex_stage/alu/r61/n62 , \dp/ex_stage/alu/r61/n61 ,
         \dp/ex_stage/alu/r61/n60 , \dp/ex_stage/alu/r61/n59 ,
         \dp/ex_stage/alu/r61/n58 , \dp/ex_stage/alu/r61/n57 ,
         \dp/ex_stage/alu/r61/n56 , \dp/ex_stage/alu/r61/n55 ,
         \dp/ex_stage/alu/r61/n54 , \dp/ex_stage/alu/r61/n53 ,
         \dp/ex_stage/alu/r61/n52 , \dp/ex_stage/alu/r61/n51 ,
         \dp/ex_stage/alu/r61/n50 , \dp/ex_stage/alu/r61/n49 ,
         \dp/ex_stage/alu/r61/n48 , \dp/ex_stage/alu/r61/n47 ,
         \dp/ex_stage/alu/r61/n46 , \dp/ex_stage/alu/r61/n45 ,
         \dp/ex_stage/alu/r61/n44 , \dp/ex_stage/alu/r61/n43 ,
         \dp/ex_stage/alu/r61/n42 , \dp/ex_stage/alu/r61/n41 ,
         \dp/ex_stage/alu/r61/n40 , \dp/ex_stage/alu/r61/n39 ,
         \dp/ex_stage/alu/r61/n38 , \dp/ex_stage/alu/r61/n37 ,
         \dp/ex_stage/alu/r61/n36 , \dp/ex_stage/alu/r61/n35 ,
         \dp/ex_stage/alu/r61/n34 , \dp/ex_stage/alu/r61/n33 ,
         \dp/ex_stage/alu/r61/n32 , \dp/ex_stage/alu/r61/n31 ,
         \dp/ex_stage/alu/r61/n30 , \dp/ex_stage/alu/r61/n29 ,
         \dp/ex_stage/alu/r61/n28 , \dp/ex_stage/alu/r61/n27 ,
         \dp/ex_stage/alu/r61/n26 , \dp/ex_stage/alu/r61/n25 ,
         \dp/ex_stage/alu/r61/n24 , \dp/ex_stage/alu/r61/n23 ,
         \dp/ex_stage/alu/r61/n22 , \dp/ex_stage/alu/r61/n21 ,
         \dp/ex_stage/alu/r61/n20 , \dp/ex_stage/alu/r61/n19 ,
         \dp/ex_stage/alu/r61/n18 , \dp/ex_stage/alu/r61/n17 ,
         \dp/ex_stage/alu/r61/n16 , \dp/ex_stage/alu/r61/n15 ,
         \dp/ex_stage/alu/r61/n14 , \dp/ex_stage/alu/r61/n13 ,
         \dp/ex_stage/alu/r61/n11 , \dp/ex_stage/alu/r61/n10 ,
         \dp/ex_stage/alu/r61/n9 , \dp/ex_stage/alu/r61/n8 ,
         \dp/ex_stage/alu/r61/n7 , \dp/ex_stage/alu/r61/n6 ,
         \dp/ex_stage/alu/r61/n5 , \dp/ex_stage/alu/r61/n4 ,
         \dp/ex_stage/alu/r61/n3 , \dp/ex_stage/alu/r61/n2 ,
         \dp/ex_stage/alu/r61/n1 , \dp/ex_stage/alu/r60/n202 ,
         \dp/ex_stage/alu/r60/n201 , \dp/ex_stage/alu/r60/n200 ,
         \dp/ex_stage/alu/r60/n199 , \dp/ex_stage/alu/r60/n198 ,
         \dp/ex_stage/alu/r60/n197 , \dp/ex_stage/alu/r60/n196 ,
         \dp/ex_stage/alu/r60/n195 , \dp/ex_stage/alu/r60/n194 ,
         \dp/ex_stage/alu/r60/n193 , \dp/ex_stage/alu/r60/n192 ,
         \dp/ex_stage/alu/r60/n191 , \dp/ex_stage/alu/r60/n190 ,
         \dp/ex_stage/alu/r60/n189 , \dp/ex_stage/alu/r60/n188 ,
         \dp/ex_stage/alu/r60/n187 , \dp/ex_stage/alu/r60/n186 ,
         \dp/ex_stage/alu/r60/n185 , \dp/ex_stage/alu/r60/n184 ,
         \dp/ex_stage/alu/r60/n183 , \dp/ex_stage/alu/r60/n182 ,
         \dp/ex_stage/alu/r60/n181 , \dp/ex_stage/alu/r60/n180 ,
         \dp/ex_stage/alu/r60/n179 , \dp/ex_stage/alu/r60/n178 ,
         \dp/ex_stage/alu/r60/n177 , \dp/ex_stage/alu/r60/n176 ,
         \dp/ex_stage/alu/r60/n175 , \dp/ex_stage/alu/r60/n174 ,
         \dp/ex_stage/alu/r60/n173 , \dp/ex_stage/alu/r60/n172 ,
         \dp/ex_stage/alu/r60/n171 , \dp/ex_stage/alu/r60/n170 ,
         \dp/ex_stage/alu/r60/n169 , \dp/ex_stage/alu/r60/n168 ,
         \dp/ex_stage/alu/r60/n167 , \dp/ex_stage/alu/r60/n166 ,
         \dp/ex_stage/alu/r60/n165 , \dp/ex_stage/alu/r60/n164 ,
         \dp/ex_stage/alu/r60/n163 , \dp/ex_stage/alu/r60/n162 ,
         \dp/ex_stage/alu/r60/n161 , \dp/ex_stage/alu/r60/n160 ,
         \dp/ex_stage/alu/r60/n159 , \dp/ex_stage/alu/r60/n158 ,
         \dp/ex_stage/alu/r60/n157 , \dp/ex_stage/alu/r60/n156 ,
         \dp/ex_stage/alu/r60/n155 , \dp/ex_stage/alu/r60/n154 ,
         \dp/ex_stage/alu/r60/n153 , \dp/ex_stage/alu/r60/n152 ,
         \dp/ex_stage/alu/r60/n151 , \dp/ex_stage/alu/r60/n150 ,
         \dp/ex_stage/alu/r60/n149 , \dp/ex_stage/alu/r60/n148 ,
         \dp/ex_stage/alu/r60/n147 , \dp/ex_stage/alu/r60/n146 ,
         \dp/ex_stage/alu/r60/n145 , \dp/ex_stage/alu/r60/n144 ,
         \dp/ex_stage/alu/r60/n143 , \dp/ex_stage/alu/r60/n142 ,
         \dp/ex_stage/alu/r60/n141 , \dp/ex_stage/alu/r60/n140 ,
         \dp/ex_stage/alu/r60/n139 , \dp/ex_stage/alu/r60/n138 ,
         \dp/ex_stage/alu/r60/n137 , \dp/ex_stage/alu/r60/n136 ,
         \dp/ex_stage/alu/r60/n135 , \dp/ex_stage/alu/r60/n134 ,
         \dp/ex_stage/alu/r60/n133 , \dp/ex_stage/alu/r60/n132 ,
         \dp/ex_stage/alu/r60/n131 , \dp/ex_stage/alu/r60/n130 ,
         \dp/ex_stage/alu/r60/n129 , \dp/ex_stage/alu/r60/n128 ,
         \dp/ex_stage/alu/r60/n127 , \dp/ex_stage/alu/r60/n126 ,
         \dp/ex_stage/alu/r60/n125 , \dp/ex_stage/alu/r60/n124 ,
         \dp/ex_stage/alu/r60/n123 , \dp/ex_stage/alu/r60/n122 ,
         \dp/ex_stage/alu/r60/n121 , \dp/ex_stage/alu/r60/n120 ,
         \dp/ex_stage/alu/r60/n119 , \dp/ex_stage/alu/r60/n118 ,
         \dp/ex_stage/alu/r60/n117 , \dp/ex_stage/alu/r60/n116 ,
         \dp/ex_stage/alu/r60/n115 , \dp/ex_stage/alu/r60/n114 ,
         \dp/ex_stage/alu/r60/n113 , \dp/ex_stage/alu/r60/n112 ,
         \dp/ex_stage/alu/r60/n111 , \dp/ex_stage/alu/r60/n110 ,
         \dp/ex_stage/alu/r60/n109 , \dp/ex_stage/alu/r60/n108 ,
         \dp/ex_stage/alu/r60/n107 , \dp/ex_stage/alu/r60/n106 ,
         \dp/ex_stage/alu/r60/n105 , \dp/ex_stage/alu/r60/n104 ,
         \dp/ex_stage/alu/r60/n103 , \dp/ex_stage/alu/r60/n102 ,
         \dp/ex_stage/alu/r60/n101 , \dp/ex_stage/alu/r60/n100 ,
         \dp/ex_stage/alu/r60/n99 , \dp/ex_stage/alu/r60/n98 ,
         \dp/ex_stage/alu/r60/n97 , \dp/ex_stage/alu/r60/n96 ,
         \dp/ex_stage/alu/r60/n95 , \dp/ex_stage/alu/r60/n94 ,
         \dp/ex_stage/alu/r60/n93 , \dp/ex_stage/alu/r60/n92 ,
         \dp/ex_stage/alu/r60/n91 , \dp/ex_stage/alu/r60/n90 ,
         \dp/ex_stage/alu/r60/n89 , \dp/ex_stage/alu/r60/n88 ,
         \dp/ex_stage/alu/r60/n87 , \dp/ex_stage/alu/r60/n86 ,
         \dp/ex_stage/alu/r60/n85 , \dp/ex_stage/alu/r60/n84 ,
         \dp/ex_stage/alu/r60/n83 , \dp/ex_stage/alu/r60/n82 ,
         \dp/ex_stage/alu/r60/n81 , \dp/ex_stage/alu/r60/n80 ,
         \dp/ex_stage/alu/r60/n79 , \dp/ex_stage/alu/r60/n78 ,
         \dp/ex_stage/alu/r60/n77 , \dp/ex_stage/alu/r60/n76 ,
         \dp/ex_stage/alu/r60/n75 , \dp/ex_stage/alu/r60/n74 ,
         \dp/ex_stage/alu/r60/n73 , \dp/ex_stage/alu/r60/n72 ,
         \dp/ex_stage/alu/r60/n71 , \dp/ex_stage/alu/r60/n70 ,
         \dp/ex_stage/alu/r60/n69 , \dp/ex_stage/alu/r60/n68 ,
         \dp/ex_stage/alu/r60/n67 , \dp/ex_stage/alu/r60/n66 ,
         \dp/ex_stage/alu/r60/n65 , \dp/ex_stage/alu/r60/n64 ,
         \dp/ex_stage/alu/r60/n63 , \dp/ex_stage/alu/r60/n62 ,
         \dp/ex_stage/alu/r60/n61 , \dp/ex_stage/alu/r60/n60 ,
         \dp/ex_stage/alu/r60/n59 , \dp/ex_stage/alu/r60/n58 ,
         \dp/ex_stage/alu/r60/n57 , \dp/ex_stage/alu/r60/n56 ,
         \dp/ex_stage/alu/r60/n55 , \dp/ex_stage/alu/r60/n54 ,
         \dp/ex_stage/alu/r60/n53 , \dp/ex_stage/alu/r60/n52 ,
         \dp/ex_stage/alu/r60/n51 , \dp/ex_stage/alu/r60/n50 ,
         \dp/ex_stage/alu/r60/n49 , \dp/ex_stage/alu/r60/n48 ,
         \dp/ex_stage/alu/r60/n47 , \dp/ex_stage/alu/r60/n46 ,
         \dp/ex_stage/alu/r60/n45 , \dp/ex_stage/alu/r60/n44 ,
         \dp/ex_stage/alu/r60/n43 , \dp/ex_stage/alu/r60/n42 ,
         \dp/ex_stage/alu/r60/n41 , \dp/ex_stage/alu/r60/n40 ,
         \dp/ex_stage/alu/r60/n39 , \dp/ex_stage/alu/r60/n38 ,
         \dp/ex_stage/alu/r60/n37 , \dp/ex_stage/alu/r60/n36 ,
         \dp/ex_stage/alu/r60/n35 , \dp/ex_stage/alu/r60/n34 ,
         \dp/ex_stage/alu/r60/n33 , \dp/ex_stage/alu/r60/n32 ,
         \dp/ex_stage/alu/r60/n31 , \dp/ex_stage/alu/r60/n30 ,
         \dp/ex_stage/alu/r60/n29 , \dp/ex_stage/alu/r60/n28 ,
         \dp/ex_stage/alu/r60/n27 , \dp/ex_stage/alu/r60/n26 ,
         \dp/ex_stage/alu/r60/n25 , \dp/ex_stage/alu/r60/n24 ,
         \dp/ex_stage/alu/r60/n23 , \dp/ex_stage/alu/r60/n22 ,
         \dp/ex_stage/alu/r60/n21 , \dp/ex_stage/alu/r60/n20 ,
         \dp/ex_stage/alu/r60/n19 , \dp/ex_stage/alu/r60/n18 ,
         \dp/ex_stage/alu/r60/n17 , \dp/ex_stage/alu/r60/n16 ,
         \dp/ex_stage/alu/r60/n15 , \dp/ex_stage/alu/r60/n14 ,
         \dp/ex_stage/alu/r60/n12 , \dp/ex_stage/alu/r60/n10 ,
         \dp/ex_stage/alu/r60/n9 , \dp/ex_stage/alu/r60/n8 ,
         \dp/ex_stage/alu/r60/n7 , \dp/ex_stage/alu/r60/n6 ,
         \dp/ex_stage/alu/r60/n5 , \dp/ex_stage/alu/r60/n4 ,
         \dp/ex_stage/alu/r60/n3 , \dp/ex_stage/alu/r60/n2 ,
         \dp/ex_stage/alu/r60/n1 ;
  wire   [31:0] instr_i;
  wire   [4:0] alu_op_i;
  wire   [7:1] \CU_I/cw2 ;
  wire   [4:0] \dp/rd_fwd_ex_o ;
  wire   [31:0] \dp/data_mem_ex_o ;
  wire   [31:0] \dp/alu_out_ex_o ;
  wire   [31:0] \dp/npc_ex_i ;
  wire   [31:0] \dp/imm_ex_i ;
  wire   [31:0] \dp/rf_out1_ex_i ;
  wire   [4:0] \dp/rd_fwd_id_o ;
  wire   [31:0] \dp/npc_id_o ;
  wire   [31:0] \dp/imm_id_o ;
  wire   [31:0] \dp/rf_out2_id_o ;
  wire   [31:0] \dp/rf_out1_id_o ;
  wire   [31:0] \dp/wr_data_id_i ;
  wire   [4:0] \dp/rd_fwd_wb_i ;
  wire   [31:0] \dp/npc_if_o ;
  wire   [31:0] \dp/if_stage/NPC_4_i ;
  wire   [31:0] \dp/id_stage/out2_i ;
  wire   [31:0] \dp/id_stage/out1_i ;
  wire   [4:0] \dp/id_stage/p_addr_wRD ;
  wire   [4:0] \dp/id_stage/p_addr_wRS2 ;
  wire   [4:0] \dp/id_stage/p_addr_wRS1 ;
  wire   [3:0] \dp/id_stage/regfile/ControlUnit/next_state ;
  wire   [5:0] \dp/id_stage/regfile/DataPath/mux_wr_out ;
  wire   [5:0] \dp/id_stage/regfile/DataPath/mux_rd_out ;
  wire   [5:0] \dp/id_stage/regfile/DataPath/addr_w_p ;
  wire   [5:0] \dp/id_stage/regfile/DataPath/addr_rd2_p ;
  wire   [5:0] \dp/id_stage/regfile/DataPath/addr_rd1_p ;
  wire   [31:0] \dp/ex_stage/muxB_out ;
  wire   [31:0] \dp/ex_stage/muxA_out ;
  wire   [31:0] \dp/ex_stage/alu/shifter_out ;
  wire   [31:0] \dp/ex_stage/alu/adder_out ;
  wire   [7:0] \dp/ex_stage/alu/adder/carries ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 ;
  wire   [3:0] \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 ;
  tri   [31:0] DRAM_DATA;
  tri   [31:0] \dp/z_word ;
  assign instr_i[31] = IRAM_DATA[31];
  assign instr_i[30] = IRAM_DATA[30];
  assign instr_i[29] = IRAM_DATA[29];
  assign instr_i[28] = IRAM_DATA[28];
  assign instr_i[27] = IRAM_DATA[27];
  assign instr_i[26] = IRAM_DATA[26];
  assign instr_i[25] = IRAM_DATA[25];
  assign instr_i[24] = IRAM_DATA[24];
  assign instr_i[23] = IRAM_DATA[23];
  assign instr_i[22] = IRAM_DATA[22];
  assign instr_i[21] = IRAM_DATA[21];
  assign instr_i[20] = IRAM_DATA[20];
  assign instr_i[19] = IRAM_DATA[19];
  assign instr_i[18] = IRAM_DATA[18];
  assign instr_i[17] = IRAM_DATA[17];
  assign instr_i[16] = IRAM_DATA[16];
  assign instr_i[15] = IRAM_DATA[15];
  assign instr_i[14] = IRAM_DATA[14];
  assign instr_i[13] = IRAM_DATA[13];
  assign instr_i[12] = IRAM_DATA[12];
  assign instr_i[11] = IRAM_DATA[11];
  assign instr_i[10] = IRAM_DATA[10];
  assign instr_i[9] = IRAM_DATA[9];
  assign instr_i[8] = IRAM_DATA[8];
  assign instr_i[7] = IRAM_DATA[7];
  assign instr_i[6] = IRAM_DATA[6];
  assign instr_i[5] = IRAM_DATA[5];
  assign instr_i[4] = IRAM_DATA[4];
  assign instr_i[3] = IRAM_DATA[3];
  assign instr_i[2] = IRAM_DATA[2];
  assign instr_i[1] = IRAM_DATA[1];
  assign instr_i[0] = IRAM_DATA[0];
  assign IRAM_ADDRESS[1] = \dp/if_stage/NPC_4_i  [1];
  assign IRAM_ADDRESS[0] = \dp/if_stage/NPC_4_i  [0];

  CLKBUF_X1 \CU_I/U249  ( .A(\CU_I/n56 ), .Z(\CU_I/n26 ) );
  CLKBUF_X1 \CU_I/U248  ( .A(\CU_I/n56 ), .Z(\CU_I/n25 ) );
  CLKBUF_X1 \CU_I/U247  ( .A(\CU_I/n56 ), .Z(\CU_I/n24 ) );
  CLKBUF_X1 \CU_I/U246  ( .A(\CU_I/n56 ), .Z(\CU_I/n20 ) );
  AOI22_X1 \CU_I/U245  ( .A1(\CU_I/n272 ), .A2(instr_i[2]), .B1(\CU_I/n270 ), 
        .B2(\CU_I/n94 ), .ZN(\CU_I/n93 ) );
  OR2_X1 \CU_I/U244  ( .A1(\CU_I/n93 ), .A2(instr_i[3]), .ZN(\CU_I/n88 ) );
  INV_X1 \CU_I/U243  ( .A(RST), .ZN(\CU_I/n56 ) );
  INV_X1 \CU_I/U242  ( .A(instr_i[26]), .ZN(\CU_I/n263 ) );
  INV_X1 \CU_I/U241  ( .A(instr_i[4]), .ZN(\CU_I/n267 ) );
  INV_X1 \CU_I/U240  ( .A(\CU_I/n126 ), .ZN(\CU_I/n266 ) );
  OR3_X1 \CU_I/U239  ( .A1(\CU_I/n157 ), .A2(instr_i[28]), .A3(\CU_I/n76 ), 
        .ZN(\CU_I/n116 ) );
  NAND2_X1 \CU_I/U238  ( .A1(\CU_I/n91 ), .A2(\CU_I/n92 ), .ZN(\CU_I/n90 ) );
  INV_X1 \CU_I/U237  ( .A(instr_i[5]), .ZN(\CU_I/n265 ) );
  INV_X1 \CU_I/U236  ( .A(instr_i[31]), .ZN(\CU_I/n67 ) );
  INV_X1 \CU_I/U235  ( .A(instr_i[27]), .ZN(\CU_I/n260 ) );
  NAND4_X1 \CU_I/U234  ( .A1(\CU_I/n91 ), .A2(instr_i[1]), .A3(instr_i[0]), 
        .A4(\CU_I/n270 ), .ZN(\CU_I/n128 ) );
  NAND2_X1 \CU_I/U233  ( .A1(\CU_I/n127 ), .A2(\CU_I/n128 ), .ZN(\CU_I/n105 )
         );
  NOR2_X1 \CU_I/U232  ( .A1(instr_i[2]), .A2(\CU_I/n272 ), .ZN(\CU_I/n144 ) );
  OAI22_X1 \CU_I/U215  ( .A1(instr_i[0]), .A2(\CU_I/n271 ), .B1(\CU_I/n272 ), 
        .B2(\CU_I/n119 ), .ZN(\CU_I/n135 ) );
  NAND4_X1 \CU_I/U214  ( .A1(\CU_I/n107 ), .A2(instr_i[5]), .A3(\CU_I/n135 ), 
        .A4(\CU_I/n269 ), .ZN(\CU_I/n129 ) );
  NAND4_X1 \CU_I/U213  ( .A1(\CU_I/n107 ), .A2(instr_i[5]), .A3(instr_i[0]), 
        .A4(\CU_I/n108 ), .ZN(\CU_I/n103 ) );
  INV_X1 \CU_I/U212  ( .A(instr_i[1]), .ZN(\CU_I/n271 ) );
  NAND2_X1 \CU_I/U211  ( .A1(instr_i[2]), .A2(instr_i[1]), .ZN(\CU_I/n108 ) );
  NOR2_X1 \CU_I/U210  ( .A1(instr_i[28]), .A2(instr_i[29]), .ZN(\CU_I/n201 )
         );
  AOI21_X1 \CU_I/U209  ( .B1(\CU_I/n259 ), .B2(\CU_I/n257 ), .A(instr_i[30]), 
        .ZN(\CU_I/n162 ) );
  AOI21_X1 \CU_I/U208  ( .B1(instr_i[29]), .B2(\CU_I/n262 ), .A(\CU_I/n76 ), 
        .ZN(\CU_I/n163 ) );
  INV_X1 \CU_I/U207  ( .A(instr_i[2]), .ZN(\CU_I/n270 ) );
  INV_X1 \CU_I/U206  ( .A(instr_i[30]), .ZN(\CU_I/n76 ) );
  NOR2_X1 \CU_I/U205  ( .A1(\CU_I/n67 ), .A2(instr_i[30]), .ZN(\CU_I/n161 ) );
  NAND4_X1 \CU_I/U204  ( .A1(\CU_I/n161 ), .A2(\CU_I/n154 ), .A3(instr_i[29]), 
        .A4(\CU_I/n257 ), .ZN(\CU_I/n187 ) );
  NAND2_X1 \CU_I/U203  ( .A1(instr_i[29]), .A2(\CU_I/n67 ), .ZN(\CU_I/n157 )
         );
  NOR2_X1 \CU_I/U202  ( .A1(\CU_I/n114 ), .A2(instr_i[4]), .ZN(\CU_I/n107 ) );
  OAI221_X1 \CU_I/U201  ( .B1(instr_i[27]), .B2(\CU_I/n256 ), .C1(\CU_I/n157 ), 
        .C2(\CU_I/n258 ), .A(\CU_I/n158 ), .ZN(\CU_I/n156 ) );
  INV_X1 \CU_I/U200  ( .A(instr_i[29]), .ZN(\CU_I/n255 ) );
  NOR3_X1 \CU_I/U199  ( .A1(\CU_I/n76 ), .A2(\CU_I/n255 ), .A3(\CU_I/n67 ), 
        .ZN(\CU_I/n205 ) );
  NOR3_X1 \CU_I/U198  ( .A1(instr_i[30]), .A2(instr_i[31]), .A3(instr_i[29]), 
        .ZN(\CU_I/n202 ) );
  INV_X1 \CU_I/U197  ( .A(instr_i[3]), .ZN(\CU_I/n269 ) );
  NOR3_X1 \CU_I/U196  ( .A1(\CU_I/n76 ), .A2(instr_i[31]), .A3(\CU_I/n256 ), 
        .ZN(\CU_I/n153 ) );
  AOI211_X1 \CU_I/U195  ( .C1(\CU_I/n122 ), .C2(\CU_I/n272 ), .A(instr_i[4]), 
        .B(\CU_I/n94 ), .ZN(\CU_I/n121 ) );
  AOI21_X1 \CU_I/U194  ( .B1(\CU_I/n272 ), .B2(\CU_I/n269 ), .A(\CU_I/n108 ), 
        .ZN(\CU_I/n120 ) );
  OAI222_X1 \CU_I/U193  ( .A1(\CU_I/n269 ), .A2(\CU_I/n119 ), .B1(instr_i[5]), 
        .B2(\CU_I/n120 ), .C1(\CU_I/n121 ), .C2(\CU_I/n270 ), .ZN(\CU_I/n118 )
         );
  AOI221_X1 \CU_I/U192  ( .B1(\CU_I/n106 ), .B2(instr_i[1]), .C1(instr_i[4]), 
        .C2(\CU_I/n269 ), .A(\CU_I/n118 ), .ZN(\CU_I/n113 ) );
  OAI22_X1 \CU_I/U191  ( .A1(instr_i[3]), .A2(\CU_I/n272 ), .B1(\CU_I/n144 ), 
        .B2(\CU_I/n264 ), .ZN(\CU_I/n142 ) );
  AOI21_X1 \CU_I/U190  ( .B1(\CU_I/n106 ), .B2(\CU_I/n119 ), .A(\CU_I/n267 ), 
        .ZN(\CU_I/n143 ) );
  OAI211_X1 \CU_I/U189  ( .C1(instr_i[1]), .C2(\CU_I/n269 ), .A(\CU_I/n272 ), 
        .B(instr_i[2]), .ZN(\CU_I/n141 ) );
  AOI221_X1 \CU_I/U188  ( .B1(\CU_I/n141 ), .B2(\CU_I/n265 ), .C1(instr_i[1]), 
        .C2(\CU_I/n142 ), .A(\CU_I/n143 ), .ZN(\CU_I/n139 ) );
  INV_X1 \CU_I/U187  ( .A(instr_i[28]), .ZN(\CU_I/n257 ) );
  NOR4_X1 \CU_I/U186  ( .A1(instr_i[30]), .A2(instr_i[29]), .A3(\CU_I/n257 ), 
        .A4(\CU_I/n260 ), .ZN(\CU_I/n150 ) );
  NOR3_X1 \CU_I/U185  ( .A1(\CU_I/n73 ), .A2(instr_i[5]), .A3(\CU_I/n108 ), 
        .ZN(\CU_I/n85 ) );
  INV_X1 \CU_I/U184  ( .A(instr_i[0]), .ZN(\CU_I/n272 ) );
  NOR2_X1 \CU_I/U183  ( .A1(instr_i[27]), .A2(instr_i[26]), .ZN(\CU_I/n160 )
         );
  NOR2_X1 \CU_I/U182  ( .A1(\CU_I/n260 ), .A2(instr_i[26]), .ZN(\CU_I/n132 )
         );
  NOR3_X1 \CU_I/U181  ( .A1(\CU_I/n157 ), .A2(instr_i[30]), .A3(\CU_I/n257 ), 
        .ZN(\CU_I/n152 ) );
  NOR3_X1 \CU_I/U180  ( .A1(instr_i[28]), .A2(instr_i[30]), .A3(\CU_I/n157 ), 
        .ZN(\CU_I/n133 ) );
  AOI22_X1 \CU_I/U179  ( .A1(\CU_I/n45 ), .A2(\CU_I/cw1[1] ), .B1(\CU_I/n171 ), 
        .B2(\CU_I/n172 ), .ZN(\CU_I/n170 ) );
  INV_X1 \CU_I/U178  ( .A(\CU_I/n170 ), .ZN(\CU_I/n52 ) );
  AOI22_X1 \CU_I/U177  ( .A1(\CU_I/n46 ), .A2(\CU_I/cw3[4] ), .B1(\CU_I/n172 ), 
        .B2(\CU_I/cw2 [4]), .ZN(\CU_I/n210 ) );
  INV_X1 \CU_I/U176  ( .A(\CU_I/n210 ), .ZN(\CU_I/n50 ) );
  AOI22_X1 \CU_I/U175  ( .A1(\CU_I/n45 ), .A2(\CU_I/cw3[5] ), .B1(\CU_I/n172 ), 
        .B2(\CU_I/cw2 [5]), .ZN(\CU_I/n208 ) );
  INV_X1 \CU_I/U174  ( .A(\CU_I/n208 ), .ZN(\CU_I/n51 ) );
  NAND2_X1 \CU_I/U173  ( .A1(regrd_sel_i), .A2(\CU_I/n42 ), .ZN(\CU_I/n190 )
         );
  INV_X1 \CU_I/U172  ( .A(\CU_I/n185 ), .ZN(\CU_I/n60 ) );
  OAI21_X1 \CU_I/U171  ( .B1(\CU_I/n60 ), .B2(\CU_I/n1 ), .A(\CU_I/n190 ), 
        .ZN(\CU_I/n247 ) );
  NAND2_X1 \CU_I/U170  ( .A1(rf_rs2_en_i), .A2(\CU_I/n43 ), .ZN(\CU_I/n198 )
         );
  AND3_X1 \CU_I/U169  ( .A1(\CU_I/n114 ), .A2(\CU_I/n196 ), .A3(\CU_I/n187 ), 
        .ZN(\CU_I/n197 ) );
  OAI21_X1 \CU_I/U168  ( .B1(\CU_I/n197 ), .B2(\CU_I/n1 ), .A(\CU_I/n198 ), 
        .ZN(\CU_I/n251 ) );
  NAND2_X1 \CU_I/U167  ( .A1(imm_uns_i), .A2(\CU_I/n43 ), .ZN(\CU_I/n193 ) );
  NOR2_X1 \CU_I/U166  ( .A1(\CU_I/n68 ), .A2(\CU_I/n194 ), .ZN(\CU_I/n192 ) );
  OAI21_X1 \CU_I/U165  ( .B1(\CU_I/n192 ), .B2(\CU_I/n1 ), .A(\CU_I/n193 ), 
        .ZN(\CU_I/n249 ) );
  NAND2_X1 \CU_I/U164  ( .A1(imm_isoff_i), .A2(\CU_I/n43 ), .ZN(\CU_I/n195 )
         );
  OAI21_X1 \CU_I/U163  ( .B1(\CU_I/n69 ), .B2(\CU_I/n1 ), .A(\CU_I/n195 ), 
        .ZN(\CU_I/n250 ) );
  NAND2_X1 \CU_I/U162  ( .A1(rf_rs1_en_i), .A2(\CU_I/n44 ), .ZN(\CU_I/n200 )
         );
  NOR4_X1 \CU_I/U161  ( .A1(\CU_I/n68 ), .A2(\CU_I/n179 ), .A3(\CU_I/n184 ), 
        .A4(\CU_I/n181 ), .ZN(\CU_I/n199 ) );
  OAI21_X1 \CU_I/U160  ( .B1(\CU_I/n199 ), .B2(\CU_I/n1 ), .A(\CU_I/n200 ), 
        .ZN(\CU_I/n252 ) );
  OAI21_X1 \CU_I/U159  ( .B1(pipe_if_id_en_i), .B2(\CU_I/n6 ), .A(\CU_I/n182 ), 
        .ZN(\CU_I/n243 ) );
  OAI21_X1 \CU_I/U158  ( .B1(\CU_I/n2 ), .B2(pc_latch_en_i), .A(\CU_I/n182 ), 
        .ZN(\CU_I/n248 ) );
  NAND2_X1 \CU_I/U157  ( .A1(DRAM_READNOTWRITE), .A2(\CU_I/n44 ), .ZN(
        \CU_I/n209 ) );
  OAI211_X1 \CU_I/U156  ( .C1(\CU_I/n46 ), .C2(\CU_I/n16 ), .A(\CU_I/n80 ), 
        .B(\CU_I/n209 ), .ZN(\CU_I/n253 ) );
  NAND2_X1 \CU_I/U155  ( .A1(alu_op_i[4]), .A2(\CU_I/n41 ), .ZN(\CU_I/n83 ) );
  OAI211_X1 \CU_I/U154  ( .C1(\CU_I/n46 ), .C2(\CU_I/n33 ), .A(\CU_I/n80 ), 
        .B(\CU_I/n83 ), .ZN(\CU_I/n215 ) );
  NAND2_X1 \CU_I/U153  ( .A1(alu_op_i[2]), .A2(\CU_I/n40 ), .ZN(\CU_I/n81 ) );
  OAI211_X1 \CU_I/U152  ( .C1(\CU_I/n46 ), .C2(\CU_I/n35 ), .A(\CU_I/n80 ), 
        .B(\CU_I/n81 ), .ZN(\CU_I/n213 ) );
  NAND2_X1 \CU_I/U151  ( .A1(muxA_sel_i), .A2(\CU_I/n41 ), .ZN(\CU_I/n166 ) );
  OAI21_X1 \CU_I/U150  ( .B1(\CU_I/n18 ), .B2(\CU_I/n3 ), .A(\CU_I/n166 ), 
        .ZN(\CU_I/n226 ) );
  NAND2_X1 \CU_I/U149  ( .A1(muxB_sel_i), .A2(\CU_I/n43 ), .ZN(\CU_I/n167 ) );
  OAI21_X1 \CU_I/U148  ( .B1(\CU_I/n18 ), .B2(\CU_I/n4 ), .A(\CU_I/n167 ), 
        .ZN(\CU_I/n227 ) );
  NAND2_X1 \CU_I/U147  ( .A1(mem_in_en_i), .A2(\CU_I/n42 ), .ZN(\CU_I/n168 )
         );
  OAI21_X1 \CU_I/U146  ( .B1(\CU_I/n18 ), .B2(\CU_I/n5 ), .A(\CU_I/n168 ), 
        .ZN(\CU_I/n228 ) );
  NAND2_X1 \CU_I/U145  ( .A1(npc_wb_en_i), .A2(\CU_I/n42 ), .ZN(\CU_I/n169 )
         );
  OAI21_X1 \CU_I/U144  ( .B1(\CU_I/n18 ), .B2(\CU_I/n6 ), .A(\CU_I/n169 ), 
        .ZN(\CU_I/n229 ) );
  NAND2_X1 \CU_I/U143  ( .A1(wb_mux_sel_i), .A2(\CU_I/n41 ), .ZN(\CU_I/n165 )
         );
  OAI21_X1 \CU_I/U142  ( .B1(\CU_I/n18 ), .B2(\CU_I/n31 ), .A(\CU_I/n165 ), 
        .ZN(\CU_I/n222 ) );
  NAND2_X1 \CU_I/U141  ( .A1(rf_we_i), .A2(\CU_I/n41 ), .ZN(\CU_I/n164 ) );
  OAI21_X1 \CU_I/U140  ( .B1(\CU_I/n18 ), .B2(\CU_I/n32 ), .A(\CU_I/n164 ), 
        .ZN(\CU_I/n221 ) );
  NAND2_X1 \CU_I/U139  ( .A1(alu_op_i[3]), .A2(\CU_I/n40 ), .ZN(\CU_I/n82 ) );
  OAI21_X1 \CU_I/U138  ( .B1(\CU_I/n18 ), .B2(\CU_I/n34 ), .A(\CU_I/n82 ), 
        .ZN(\CU_I/n214 ) );
  NAND2_X1 \CU_I/U137  ( .A1(alu_op_i[1]), .A2(\CU_I/n40 ), .ZN(\CU_I/n79 ) );
  OAI21_X1 \CU_I/U136  ( .B1(\CU_I/n18 ), .B2(\CU_I/n36 ), .A(\CU_I/n79 ), 
        .ZN(\CU_I/n212 ) );
  NAND2_X1 \CU_I/U135  ( .A1(alu_op_i[0]), .A2(\CU_I/n42 ), .ZN(\CU_I/n77 ) );
  OAI21_X1 \CU_I/U134  ( .B1(\CU_I/n18 ), .B2(\CU_I/n37 ), .A(\CU_I/n77 ), 
        .ZN(\CU_I/n211 ) );
  NAND2_X1 \CU_I/U133  ( .A1(pipe_clear_n_i), .A2(\CU_I/n30 ), .ZN(jump_en_i)
         );
  INV_X1 \CU_I/U132  ( .A(\CU_I/n187 ), .ZN(\CU_I/n57 ) );
  NOR4_X1 \CU_I/U131  ( .A1(\CU_I/n57 ), .A2(\CU_I/n184 ), .A3(\CU_I/n185 ), 
        .A4(\CU_I/n186 ), .ZN(\CU_I/n183 ) );
  OAI22_X1 \CU_I/U130  ( .A1(pipe_if_id_en_i), .A2(\CU_I/n4 ), .B1(\CU_I/n183 ), .B2(\CU_I/n1 ), .ZN(\CU_I/n245 ) );
  OAI22_X1 \CU_I/U129  ( .A1(pc_latch_en_i), .A2(\CU_I/n23 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n13 ), .ZN(\CU_I/n236 ) );
  NOR4_X1 \CU_I/U128  ( .A1(\CU_I/n96 ), .A2(\CU_I/n97 ), .A3(\CU_I/n98 ), 
        .A4(\CU_I/n99 ), .ZN(\CU_I/n95 ) );
  OAI22_X1 \CU_I/U127  ( .A1(pc_latch_en_i), .A2(\CU_I/n36 ), .B1(\CU_I/n95 ), 
        .B2(\CU_I/n1 ), .ZN(\CU_I/n217 ) );
  OAI211_X1 \CU_I/U126  ( .C1(\CU_I/n73 ), .C2(\CU_I/n88 ), .A(\CU_I/n89 ), 
        .B(\CU_I/n90 ), .ZN(\CU_I/n86 ) );
  INV_X1 \CU_I/U125  ( .A(\CU_I/n87 ), .ZN(\CU_I/n61 ) );
  AOI211_X1 \CU_I/U124  ( .C1(\CU_I/n85 ), .C2(\CU_I/n272 ), .A(\CU_I/n86 ), 
        .B(\CU_I/n61 ), .ZN(\CU_I/n84 ) );
  OAI22_X1 \CU_I/U123  ( .A1(pc_latch_en_i), .A2(\CU_I/n37 ), .B1(\CU_I/n84 ), 
        .B2(\CU_I/n1 ), .ZN(\CU_I/n216 ) );
  OAI22_X1 \CU_I/U122  ( .A1(pc_latch_en_i), .A2(\CU_I/n11 ), .B1(\CU_I/n69 ), 
        .B2(\CU_I/n1 ), .ZN(\CU_I/n238 ) );
  OAI22_X1 \CU_I/U121  ( .A1(pc_latch_en_i), .A2(\CU_I/n12 ), .B1(\CU_I/n62 ), 
        .B2(\CU_I/n1 ), .ZN(\CU_I/n237 ) );
  INV_X1 \CU_I/U120  ( .A(\CU_I/n181 ), .ZN(\CU_I/n58 ) );
  OAI22_X1 \CU_I/U119  ( .A1(pipe_if_id_en_i), .A2(\CU_I/n7 ), .B1(\CU_I/n58 ), 
        .B2(\CU_I/n1 ), .ZN(\CU_I/n242 ) );
  NOR4_X1 \CU_I/U118  ( .A1(\CU_I/n64 ), .A2(\CU_I/n149 ), .A3(\CU_I/n150 ), 
        .A4(\CU_I/n66 ), .ZN(\CU_I/n148 ) );
  AOI22_X1 \CU_I/U117  ( .A1(\CU_I/n59 ), .A2(\CU_I/n257 ), .B1(instr_i[30]), 
        .B2(\CU_I/n156 ), .ZN(\CU_I/n147 ) );
  OAI21_X1 \CU_I/U116  ( .B1(\CU_I/n162 ), .B2(\CU_I/n163 ), .A(instr_i[31]), 
        .ZN(\CU_I/n146 ) );
  NAND4_X1 \CU_I/U115  ( .A1(\CU_I/n145 ), .A2(\CU_I/n146 ), .A3(\CU_I/n147 ), 
        .A4(\CU_I/n148 ), .ZN(\CU_I/n112 ) );
  OAI22_X1 \CU_I/U114  ( .A1(pipe_if_id_en_i), .A2(\CU_I/n27 ), .B1(\CU_I/n14 ), .B2(\CU_I/n15 ), .ZN(\CU_I/n254 ) );
  OAI22_X1 \CU_I/U113  ( .A1(pc_latch_en_i), .A2(\CU_I/n22 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n12 ), .ZN(\CU_I/n235 ) );
  OAI22_X1 \CU_I/U112  ( .A1(pc_latch_en_i), .A2(\CU_I/n21 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n11 ), .ZN(\CU_I/n234 ) );
  OAI22_X1 \CU_I/U111  ( .A1(pc_latch_en_i), .A2(\CU_I/n19 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n10 ), .ZN(\CU_I/n233 ) );
  OAI22_X1 \CU_I/U110  ( .A1(pc_latch_en_i), .A2(\CU_I/n17 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n9 ), .ZN(\CU_I/n232 ) );
  OAI22_X1 \CU_I/U109  ( .A1(pc_latch_en_i), .A2(\CU_I/n15 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n7 ), .ZN(\CU_I/n230 ) );
  OAI22_X1 \CU_I/U108  ( .A1(pc_latch_en_i), .A2(\CU_I/n30 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n21 ), .ZN(\CU_I/n225 ) );
  OAI22_X1 \CU_I/U107  ( .A1(pc_latch_en_i), .A2(\CU_I/n31 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n22 ), .ZN(\CU_I/n224 ) );
  OAI22_X1 \CU_I/U106  ( .A1(pc_latch_en_i), .A2(\CU_I/n32 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n23 ), .ZN(\CU_I/n223 ) );
  INV_X1 \CU_I/U105  ( .A(\CU_I/n145 ), .ZN(\CU_I/n48 ) );
  NOR4_X1 \CU_I/U104  ( .A1(\CU_I/n68 ), .A2(\CU_I/n176 ), .A3(\CU_I/n48 ), 
        .A4(\CU_I/n171 ), .ZN(\CU_I/n175 ) );
  OAI22_X1 \CU_I/U103  ( .A1(pc_latch_en_i), .A2(\CU_I/n8 ), .B1(\CU_I/n175 ), 
        .B2(\CU_I/n44 ), .ZN(\CU_I/n241 ) );
  INV_X1 \CU_I/U102  ( .A(\CU_I/n99 ), .ZN(\CU_I/n63 ) );
  OAI211_X1 \CU_I/U101  ( .C1(\CU_I/n113 ), .C2(\CU_I/n114 ), .A(\CU_I/n115 ), 
        .B(\CU_I/n63 ), .ZN(\CU_I/n110 ) );
  NOR3_X1 \CU_I/U100  ( .A1(\CU_I/n110 ), .A2(\CU_I/n111 ), .A3(\CU_I/n112 ), 
        .ZN(\CU_I/n109 ) );
  OAI22_X1 \CU_I/U99  ( .A1(pc_latch_en_i), .A2(\CU_I/n35 ), .B1(\CU_I/n109 ), 
        .B2(\CU_I/n45 ), .ZN(\CU_I/n218 ) );
  OAI211_X1 \CU_I/U98  ( .C1(\CU_I/n259 ), .C2(\CU_I/n116 ), .A(\CU_I/n70 ), 
        .B(\CU_I/n101 ), .ZN(\CU_I/n137 ) );
  OAI21_X1 \CU_I/U97  ( .B1(\CU_I/n139 ), .B2(\CU_I/n114 ), .A(\CU_I/n140 ), 
        .ZN(\CU_I/n138 ) );
  NOR3_X1 \CU_I/U96  ( .A1(\CU_I/n137 ), .A2(\CU_I/n112 ), .A3(\CU_I/n138 ), 
        .ZN(\CU_I/n136 ) );
  OAI22_X1 \CU_I/U95  ( .A1(pc_latch_en_i), .A2(\CU_I/n33 ), .B1(\CU_I/n136 ), 
        .B2(\CU_I/n44 ), .ZN(\CU_I/n220 ) );
  NOR3_X1 \CU_I/U94  ( .A1(\CU_I/n124 ), .A2(\CU_I/n105 ), .A3(\CU_I/n125 ), 
        .ZN(\CU_I/n123 ) );
  OAI22_X1 \CU_I/U93  ( .A1(pc_latch_en_i), .A2(\CU_I/n34 ), .B1(\CU_I/n123 ), 
        .B2(\CU_I/n1 ), .ZN(\CU_I/n219 ) );
  OAI22_X1 \CU_I/U92  ( .A1(pc_latch_en_i), .A2(\CU_I/n9 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n174 ), .ZN(\CU_I/n240 ) );
  OAI22_X1 \CU_I/U91  ( .A1(pc_latch_en_i), .A2(\CU_I/n10 ), .B1(\CU_I/n14 ), 
        .B2(\CU_I/n173 ), .ZN(\CU_I/n239 ) );
  OAI22_X1 \CU_I/U90  ( .A1(pipe_if_id_en_i), .A2(\CU_I/n5 ), .B1(\CU_I/n18 ), 
        .B2(\CU_I/n178 ), .ZN(\CU_I/n244 ) );
  OAI221_X1 \CU_I/U89  ( .B1(\CU_I/n40 ), .B2(\CU_I/n8 ), .C1(pipe_if_id_en_i), 
        .C2(\CU_I/n16 ), .A(\CU_I/n80 ), .ZN(\CU_I/n231 ) );
  INV_X1 \CU_I/U88  ( .A(\CU_I/n189 ), .ZN(\CU_I/n75 ) );
  NOR2_X1 \CU_I/U87  ( .A1(\CU_I/n75 ), .A2(\CU_I/n184 ), .ZN(\CU_I/n188 ) );
  OAI221_X1 \CU_I/U86  ( .B1(\CU_I/n188 ), .B2(\CU_I/n18 ), .C1(
        pipe_if_id_en_i), .C2(\CU_I/n3 ), .A(\CU_I/n182 ), .ZN(\CU_I/n246 ) );
  INV_X1 \CU_I/U85  ( .A(is_zero_i), .ZN(\CU_I/n54 ) );
  AOI22_X1 \CU_I/U84  ( .A1(is_zero_i), .A2(\CU_I/cw3[4] ), .B1(\CU_I/n54 ), 
        .B2(\CU_I/cw3[5] ), .ZN(pipe_clear_n_i) );
  NAND2_X1 \CU_I/U83  ( .A1(IRAM_READY), .A2(IRAM_ISSUE), .ZN(\CU_I/n78 ) );
  NOR2_X1 \CU_I/U82  ( .A1(DRAM_READY), .A2(\CU_I/n27 ), .ZN(DRAM_ISSUE) );
  BUF_X1 \CU_I/U81  ( .A(\CU_I/n273 ), .Z(wb_mux_sel_i) );
  OAI21_X1 \CU_I/U80  ( .B1(\CU_I/n152 ), .B2(\CU_I/n153 ), .A(\CU_I/n154 ), 
        .ZN(\CU_I/n151 ) );
  INV_X1 \CU_I/U79  ( .A(\CU_I/n151 ), .ZN(\CU_I/n66 ) );
  AOI22_X1 \CU_I/U78  ( .A1(\CU_I/n157 ), .A2(\CU_I/n117 ), .B1(\CU_I/n160 ), 
        .B2(\CU_I/n161 ), .ZN(\CU_I/n159 ) );
  INV_X1 \CU_I/U77  ( .A(\CU_I/n159 ), .ZN(\CU_I/n59 ) );
  INV_X1 \CU_I/U76  ( .A(\CU_I/n201 ), .ZN(\CU_I/n256 ) );
  INV_X1 \CU_I/U75  ( .A(\CU_I/n85 ), .ZN(\CU_I/n72 ) );
  INV_X1 \CU_I/U74  ( .A(\CU_I/n107 ), .ZN(\CU_I/n73 ) );
  NOR2_X1 \CU_I/U73  ( .A1(\CU_I/n133 ), .A2(\CU_I/n194 ), .ZN(\CU_I/n203 ) );
  AND4_X1 \CU_I/U72  ( .A1(\CU_I/n89 ), .A2(\CU_I/n115 ), .A3(\CU_I/n116 ), 
        .A4(\CU_I/n203 ), .ZN(\CU_I/n191 ) );
  NAND2_X1 \CU_I/U71  ( .A1(\CU_I/n176 ), .A2(\CU_I/n132 ), .ZN(\CU_I/n189 )
         );
  NOR2_X1 \CU_I/U70  ( .A1(\CU_I/n262 ), .A2(\CU_I/n116 ), .ZN(\CU_I/n149 ) );
  INV_X1 \CU_I/U69  ( .A(\CU_I/n132 ), .ZN(\CU_I/n259 ) );
  NAND2_X1 \CU_I/U68  ( .A1(\CU_I/n153 ), .A2(\CU_I/n132 ), .ZN(\CU_I/n196 )
         );
  INV_X1 \CU_I/U67  ( .A(\CU_I/n160 ), .ZN(\CU_I/n262 ) );
  NAND2_X1 \CU_I/U66  ( .A1(\CU_I/n271 ), .A2(\CU_I/n270 ), .ZN(\CU_I/n119 )
         );
  INV_X1 \CU_I/U65  ( .A(\CU_I/n134 ), .ZN(\CU_I/n65 ) );
  AOI21_X1 \CU_I/U64  ( .B1(\CU_I/n132 ), .B2(\CU_I/n133 ), .A(\CU_I/n65 ), 
        .ZN(\CU_I/n131 ) );
  INV_X1 \CU_I/U63  ( .A(\CU_I/n106 ), .ZN(\CU_I/n268 ) );
  AOI21_X1 \CU_I/U62  ( .B1(\CU_I/n85 ), .B2(\CU_I/n268 ), .A(\CU_I/n105 ), 
        .ZN(\CU_I/n104 ) );
  INV_X1 \CU_I/U61  ( .A(\CU_I/n180 ), .ZN(\CU_I/n71 ) );
  NAND2_X1 \CU_I/U60  ( .A1(\CU_I/n207 ), .A2(\CU_I/n117 ), .ZN(\CU_I/n89 ) );
  NAND2_X1 \CU_I/U59  ( .A1(\CU_I/n178 ), .A2(\CU_I/n187 ), .ZN(\CU_I/n181 )
         );
  NAND2_X1 \CU_I/U58  ( .A1(\CU_I/n160 ), .A2(\CU_I/n207 ), .ZN(\CU_I/n115 )
         );
  NAND2_X1 \CU_I/U57  ( .A1(\CU_I/n132 ), .A2(\CU_I/n152 ), .ZN(\CU_I/n134 )
         );
  NAND2_X1 \CU_I/U56  ( .A1(\CU_I/n152 ), .A2(\CU_I/n117 ), .ZN(\CU_I/n100 )
         );
  AND2_X1 \CU_I/U55  ( .A1(\CU_I/n202 ), .A2(\CU_I/n257 ), .ZN(\CU_I/n176 ) );
  NAND2_X1 \CU_I/U54  ( .A1(\CU_I/n180 ), .A2(\CU_I/n132 ), .ZN(\CU_I/n102 )
         );
  NAND2_X1 \CU_I/U53  ( .A1(\CU_I/n154 ), .A2(\CU_I/n133 ), .ZN(\CU_I/n101 )
         );
  NAND2_X1 \CU_I/U52  ( .A1(\CU_I/n174 ), .A2(\CU_I/n173 ), .ZN(\CU_I/n184 )
         );
  NAND2_X1 \CU_I/U51  ( .A1(\CU_I/n133 ), .A2(\CU_I/n117 ), .ZN(\CU_I/n155 )
         );
  NOR2_X1 \CU_I/U50  ( .A1(\CU_I/n269 ), .A2(\CU_I/n265 ), .ZN(\CU_I/n122 ) );
  INV_X1 \CU_I/U49  ( .A(\CU_I/n117 ), .ZN(\CU_I/n261 ) );
  NOR2_X1 \CU_I/U48  ( .A1(\CU_I/n116 ), .A2(\CU_I/n261 ), .ZN(\CU_I/n99 ) );
  NAND2_X1 \CU_I/U47  ( .A1(\CU_I/n176 ), .A2(\CU_I/n160 ), .ZN(\CU_I/n114 )
         );
  AND2_X1 \CU_I/U46  ( .A1(\CU_I/n102 ), .A2(\CU_I/n127 ), .ZN(\CU_I/n206 ) );
  OAI211_X1 \CU_I/U45  ( .C1(\CU_I/n71 ), .C2(\CU_I/n262 ), .A(\CU_I/n130 ), 
        .B(\CU_I/n206 ), .ZN(\CU_I/n111 ) );
  NOR2_X1 \CU_I/U44  ( .A1(\CU_I/n269 ), .A2(\CU_I/n272 ), .ZN(\CU_I/n106 ) );
  NOR3_X1 \CU_I/U43  ( .A1(\CU_I/n257 ), .A2(\CU_I/n157 ), .A3(\CU_I/n76 ), 
        .ZN(\CU_I/n207 ) );
  NOR3_X1 \CU_I/U42  ( .A1(\CU_I/n271 ), .A2(\CU_I/n272 ), .A3(\CU_I/n265 ), 
        .ZN(\CU_I/n94 ) );
  AOI211_X1 \CU_I/U41  ( .C1(\CU_I/n152 ), .C2(\CU_I/n160 ), .A(\CU_I/n111 ), 
        .B(\CU_I/n204 ), .ZN(\CU_I/n87 ) );
  NOR2_X1 \CU_I/U40  ( .A1(\CU_I/n260 ), .A2(\CU_I/n263 ), .ZN(\CU_I/n154 ) );
  BUF_X1 \CU_I/U39  ( .A(\CU_I/n78 ), .Z(\CU_I/n29 ) );
  BUF_X1 \CU_I/U38  ( .A(\CU_I/n78 ), .Z(\CU_I/n28 ) );
  INV_X1 \CU_I/U37  ( .A(pipe_clear_n_i), .ZN(\CU_I/n53 ) );
  AOI21_X1 \CU_I/U36  ( .B1(\CU_I/n117 ), .B2(\CU_I/n180 ), .A(\CU_I/n53 ), 
        .ZN(\CU_I/n145 ) );
  INV_X1 \CU_I/U35  ( .A(DRAM_ISSUE), .ZN(IRAM_ISSUE) );
  INV_X1 \CU_I/U34  ( .A(\CU_I/n155 ), .ZN(\CU_I/n64 ) );
  INV_X1 \CU_I/U33  ( .A(\CU_I/n122 ), .ZN(\CU_I/n264 ) );
  NAND2_X1 \CU_I/U32  ( .A1(\CU_I/n176 ), .A2(\CU_I/n154 ), .ZN(\CU_I/n177 )
         );
  INV_X1 \CU_I/U31  ( .A(\CU_I/n196 ), .ZN(\CU_I/n68 ) );
  NAND2_X1 \CU_I/U30  ( .A1(\CU_I/n191 ), .A2(\CU_I/n114 ), .ZN(\CU_I/n179 )
         );
  INV_X1 \CU_I/U29  ( .A(\CU_I/n154 ), .ZN(\CU_I/n258 ) );
  NAND2_X1 \CU_I/U28  ( .A1(\CU_I/n191 ), .A2(\CU_I/n178 ), .ZN(\CU_I/n185 )
         );
  NOR2_X1 \CU_I/U27  ( .A1(\CU_I/n71 ), .A2(\CU_I/n258 ), .ZN(\CU_I/n98 ) );
  NAND4_X1 \CU_I/U26  ( .A1(\CU_I/n87 ), .A2(\CU_I/n70 ), .A3(\CU_I/n100 ), 
        .A4(\CU_I/n155 ), .ZN(\CU_I/n194 ) );
  NOR2_X1 \CU_I/U25  ( .A1(\CU_I/n264 ), .A2(\CU_I/n114 ), .ZN(\CU_I/n91 ) );
  BUF_X1 \CU_I/U24  ( .A(\CU_I/n29 ), .Z(\CU_I/n45 ) );
  BUF_X1 \CU_I/U23  ( .A(\CU_I/n29 ), .Z(\CU_I/n44 ) );
  BUF_X1 \CU_I/U22  ( .A(\CU_I/n28 ), .Z(\CU_I/n41 ) );
  BUF_X1 \CU_I/U21  ( .A(\CU_I/n29 ), .Z(\CU_I/n43 ) );
  BUF_X1 \CU_I/U20  ( .A(\CU_I/n28 ), .Z(\CU_I/n42 ) );
  BUF_X1 \CU_I/U19  ( .A(\CU_I/n28 ), .Z(\CU_I/n40 ) );
  BUF_X1 \CU_I/U18  ( .A(\CU_I/n29 ), .Z(\CU_I/n46 ) );
  NAND2_X1 \CU_I/U17  ( .A1(pipe_if_id_en_i), .A2(\CU_I/n53 ), .ZN(\CU_I/n80 )
         );
  NOR2_X1 \CU_I/U16  ( .A1(\CU_I/n45 ), .A2(\CU_I/n53 ), .ZN(\CU_I/n172 ) );
  INV_X1 \CU_I/U15  ( .A(\CU_I/n91 ), .ZN(\CU_I/n74 ) );
  INV_X1 \CU_I/U14  ( .A(\CU_I/n179 ), .ZN(\CU_I/n62 ) );
  INV_X1 \CU_I/U13  ( .A(\CU_I/n98 ), .ZN(\CU_I/n70 ) );
  INV_X1 \CU_I/U12  ( .A(\CU_I/n186 ), .ZN(\CU_I/n69 ) );
  INV_X1 \CU_I/U11  ( .A(\CU_I/n172 ), .ZN(\CU_I/n49 ) );
  OR2_X1 \CU_I/U10  ( .A1(\CU_I/n177 ), .A2(\CU_I/n18 ), .ZN(\CU_I/n182 ) );
  INV_X1 \CU_I/U9  ( .A(\CU_I/n46 ), .ZN(pc_latch_en_i) );
  INV_X1 \CU_I/U8  ( .A(\CU_I/n78 ), .ZN(pipe_if_id_en_i) );
  BUF_X1 \CU_I/U7  ( .A(\CU_I/n49 ), .Z(\CU_I/n14 ) );
  BUF_X1 \CU_I/U6  ( .A(\CU_I/n49 ), .Z(\CU_I/n1 ) );
  BUF_X1 \CU_I/U5  ( .A(\CU_I/n49 ), .Z(\CU_I/n18 ) );
  NOR2_X1 \CU_I/U4  ( .A1(\CU_I/n263 ), .A2(instr_i[27]), .ZN(\CU_I/n117 ) );
  NOR4_X1 \CU_I/U3  ( .A1(\CU_I/n76 ), .A2(\CU_I/n257 ), .A3(instr_i[29]), 
        .A4(instr_i[31]), .ZN(\CU_I/n180 ) );
  DFFR_X1 \CU_I/cw1_reg[13]  ( .D(\CU_I/n248 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        reg31_sel_i), .QN(\CU_I/n2 ) );
  DFFR_X1 \CU_I/cw2_reg[4]  ( .D(\CU_I/n233 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        \CU_I/cw2 [4]), .QN(\CU_I/n19 ) );
  DFFR_X1 \CU_I/cw2_reg[5]  ( .D(\CU_I/n232 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        \CU_I/cw2 [5]), .QN(\CU_I/n17 ) );
  DFFR_X1 \CU_I/cw1_reg[1]  ( .D(\CU_I/n52 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        \CU_I/cw1[1] ), .QN(\CU_I/n13 ) );
  DFFR_X1 \CU_I/cw1_reg[12]  ( .D(\CU_I/n247 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        regrd_sel_i) );
  DFFR_X1 \CU_I/cw1_reg[14]  ( .D(\CU_I/n249 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        imm_uns_i) );
  DFFR_X1 \CU_I/cw1_reg[15]  ( .D(\CU_I/n250 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        imm_isoff_i) );
  DFFR_X1 \CU_I/cw1_reg[16]  ( .D(\CU_I/n251 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        rf_rs2_en_i) );
  DFFR_X1 \CU_I/cw1_reg[17]  ( .D(\CU_I/n252 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        rf_rs1_en_i) );
  DFFR_X1 \CU_I/aluOpcode2_reg[0]  ( .D(\CU_I/n211 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(alu_op_i[0]) );
  DFFR_X1 \CU_I/aluOpcode2_reg[1]  ( .D(\CU_I/n212 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(alu_op_i[1]) );
  DFFR_X1 \CU_I/aluOpcode2_reg[3]  ( .D(\CU_I/n214 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(alu_op_i[3]) );
  DFFR_X1 \CU_I/cw2_reg[8]  ( .D(\CU_I/n229 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        npc_wb_en_i) );
  DFFR_X1 \CU_I/cw2_reg[9]  ( .D(\CU_I/n228 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        mem_in_en_i) );
  DFFR_X1 \CU_I/cw2_reg[10]  ( .D(\CU_I/n227 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        muxB_sel_i) );
  DFFR_X1 \CU_I/cw2_reg[11]  ( .D(\CU_I/n226 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        muxA_sel_i) );
  DFFR_X1 \CU_I/cw4_reg[1]  ( .D(\CU_I/n221 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        rf_we_i) );
  DFFR_X1 \CU_I/cw4_reg[2]  ( .D(\CU_I/n222 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        \CU_I/n273 ) );
  DFFR_X1 \CU_I/cw3_reg[4]  ( .D(\CU_I/n50 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        \CU_I/cw3[4] ) );
  DFFR_X1 \CU_I/cw3_reg[5]  ( .D(\CU_I/n51 ), .CK(CLK), .RN(\CU_I/n56 ), .Q(
        \CU_I/cw3[5] ) );
  NAND3_X1 \CU_I/U231  ( .A1(\CU_I/n117 ), .A2(instr_i[28]), .A3(\CU_I/n205 ), 
        .ZN(\CU_I/n130 ) );
  NAND3_X1 \CU_I/U230  ( .A1(\CU_I/n154 ), .A2(\CU_I/n257 ), .A3(\CU_I/n205 ), 
        .ZN(\CU_I/n127 ) );
  NAND3_X1 \CU_I/U229  ( .A1(\CU_I/n132 ), .A2(\CU_I/n257 ), .A3(\CU_I/n205 ), 
        .ZN(\CU_I/n140 ) );
  NAND3_X1 \CU_I/U228  ( .A1(\CU_I/n140 ), .A2(\CU_I/n101 ), .A3(\CU_I/n134 ), 
        .ZN(\CU_I/n204 ) );
  NAND3_X1 \CU_I/U227  ( .A1(\CU_I/n160 ), .A2(instr_i[28]), .A3(\CU_I/n202 ), 
        .ZN(\CU_I/n174 ) );
  NAND3_X1 \CU_I/U226  ( .A1(\CU_I/n117 ), .A2(instr_i[28]), .A3(\CU_I/n202 ), 
        .ZN(\CU_I/n173 ) );
  NAND3_X1 \CU_I/U225  ( .A1(\CU_I/n201 ), .A2(\CU_I/n154 ), .A3(\CU_I/n161 ), 
        .ZN(\CU_I/n178 ) );
  NAND3_X1 \CU_I/U224  ( .A1(\CU_I/n189 ), .A2(\CU_I/n196 ), .A3(\CU_I/n177 ), 
        .ZN(\CU_I/n186 ) );
  NAND3_X1 \CU_I/U223  ( .A1(\CU_I/n177 ), .A2(\CU_I/n178 ), .A3(\CU_I/n62 ), 
        .ZN(\CU_I/n171 ) );
  NAND3_X1 \CU_I/U222  ( .A1(instr_i[28]), .A2(instr_i[29]), .A3(instr_i[27]), 
        .ZN(\CU_I/n158 ) );
  NAND3_X1 \CU_I/U221  ( .A1(\CU_I/n129 ), .A2(\CU_I/n130 ), .A3(\CU_I/n131 ), 
        .ZN(\CU_I/n124 ) );
  OAI33_X1 \CU_I/U220  ( .A1(\CU_I/n267 ), .A2(\CU_I/n272 ), .A3(\CU_I/n270 ), 
        .B1(instr_i[0]), .B2(instr_i[4]), .B3(instr_i[2]), .ZN(\CU_I/n126 ) );
  OAI33_X1 \CU_I/U219  ( .A1(\CU_I/n72 ), .A2(instr_i[0]), .A3(\CU_I/n269 ), 
        .B1(\CU_I/n74 ), .B2(instr_i[1]), .B3(\CU_I/n266 ), .ZN(\CU_I/n125 )
         );
  NAND3_X1 \CU_I/U218  ( .A1(\CU_I/n103 ), .A2(\CU_I/n89 ), .A3(\CU_I/n104 ), 
        .ZN(\CU_I/n96 ) );
  NAND3_X1 \CU_I/U217  ( .A1(\CU_I/n100 ), .A2(\CU_I/n101 ), .A3(\CU_I/n102 ), 
        .ZN(\CU_I/n97 ) );
  OAI33_X1 \CU_I/U216  ( .A1(\CU_I/n267 ), .A2(instr_i[2]), .A3(\CU_I/n271 ), 
        .B1(\CU_I/n270 ), .B2(instr_i[1]), .B3(\CU_I/n272 ), .ZN(\CU_I/n92 )
         );
  DFFS_X1 \CU_I/aluOpcode2_reg[2]  ( .D(\CU_I/n213 ), .CK(CLK), .SN(\CU_I/n26 ), .Q(alu_op_i[2]) );
  DFFS_X1 \CU_I/aluOpcode2_reg[4]  ( .D(\CU_I/n215 ), .CK(CLK), .SN(\CU_I/n25 ), .Q(alu_op_i[4]) );
  DFFR_X1 \CU_I/aluOpcode1_reg[0]  ( .D(\CU_I/n216 ), .CK(CLK), .RN(\CU_I/n20 ), .QN(\CU_I/n37 ) );
  DFFR_X1 \CU_I/aluOpcode1_reg[1]  ( .D(\CU_I/n217 ), .CK(CLK), .RN(\CU_I/n20 ), .QN(\CU_I/n36 ) );
  DFFS_X1 \CU_I/aluOpcode1_reg[2]  ( .D(\CU_I/n218 ), .CK(CLK), .SN(\CU_I/n25 ), .QN(\CU_I/n35 ) );
  DFFR_X1 \CU_I/aluOpcode1_reg[3]  ( .D(\CU_I/n219 ), .CK(CLK), .RN(\CU_I/n20 ), .QN(\CU_I/n34 ) );
  DFFS_X1 \CU_I/aluOpcode1_reg[4]  ( .D(\CU_I/n220 ), .CK(CLK), .SN(\CU_I/n25 ), .QN(\CU_I/n33 ) );
  DFFR_X1 \CU_I/cw3_reg[1]  ( .D(\CU_I/n223 ), .CK(CLK), .RN(\CU_I/n20 ), .QN(
        \CU_I/n32 ) );
  DFFR_X1 \CU_I/cw3_reg[2]  ( .D(\CU_I/n224 ), .CK(CLK), .RN(\CU_I/n20 ), .QN(
        \CU_I/n31 ) );
  DFFR_X1 \CU_I/cw3_reg[3]  ( .D(\CU_I/n225 ), .CK(CLK), .RN(\CU_I/n20 ), .QN(
        \CU_I/n30 ) );
  DFFR_X1 \CU_I/cw2_reg[1]  ( .D(\CU_I/n236 ), .CK(CLK), .RN(\CU_I/n56 ), .QN(
        \CU_I/n23 ) );
  DFFS_X1 \CU_I/cw3_reg[6]  ( .D(\CU_I/n253 ), .CK(CLK), .SN(\CU_I/n25 ), .Q(
        DRAM_READNOTWRITE) );
  DFFS_X1 \CU_I/cw2_reg[6]  ( .D(\CU_I/n231 ), .CK(CLK), .SN(\CU_I/n25 ), .QN(
        \CU_I/n16 ) );
  DFFS_X1 \CU_I/cw1_reg[6]  ( .D(\CU_I/n241 ), .CK(CLK), .SN(\CU_I/n26 ), .QN(
        \CU_I/n8 ) );
  DFFR_X1 \CU_I/cw1_reg[11]  ( .D(\CU_I/n246 ), .CK(CLK), .RN(\CU_I/n24 ), 
        .QN(\CU_I/n3 ) );
  DFFR_X1 \CU_I/cw1_reg[10]  ( .D(\CU_I/n245 ), .CK(CLK), .RN(\CU_I/n24 ), 
        .QN(\CU_I/n4 ) );
  DFFR_X1 \CU_I/cw1_reg[9]  ( .D(\CU_I/n244 ), .CK(CLK), .RN(\CU_I/n24 ), .QN(
        \CU_I/n5 ) );
  DFFR_X1 \CU_I/cw1_reg[8]  ( .D(\CU_I/n243 ), .CK(CLK), .RN(\CU_I/n24 ), .QN(
        \CU_I/n6 ) );
  DFFR_X1 \CU_I/cw2_reg[7]  ( .D(\CU_I/n230 ), .CK(CLK), .RN(\CU_I/n24 ), .QN(
        \CU_I/n15 ) );
  DFFR_X1 \CU_I/cw1_reg[7]  ( .D(\CU_I/n242 ), .CK(CLK), .RN(\CU_I/n25 ), .QN(
        \CU_I/n7 ) );
  DFFR_X1 \CU_I/cw1_reg[5]  ( .D(\CU_I/n240 ), .CK(CLK), .RN(\CU_I/n25 ), .QN(
        \CU_I/n9 ) );
  DFFR_X1 \CU_I/cw1_reg[4]  ( .D(\CU_I/n239 ), .CK(CLK), .RN(\CU_I/n25 ), .QN(
        \CU_I/n10 ) );
  DFFR_X1 \CU_I/cw2_reg[3]  ( .D(\CU_I/n234 ), .CK(CLK), .RN(\CU_I/n25 ), .QN(
        \CU_I/n21 ) );
  DFFR_X1 \CU_I/cw1_reg[3]  ( .D(\CU_I/n238 ), .CK(CLK), .RN(\CU_I/n24 ), .QN(
        \CU_I/n11 ) );
  DFFR_X1 \CU_I/cw2_reg[2]  ( .D(\CU_I/n235 ), .CK(CLK), .RN(\CU_I/n25 ), .QN(
        \CU_I/n22 ) );
  DFFR_X1 \CU_I/cw1_reg[2]  ( .D(\CU_I/n237 ), .CK(CLK), .RN(\CU_I/n25 ), .QN(
        \CU_I/n12 ) );
  DFFR_X1 \CU_I/cw3_reg[7]  ( .D(\CU_I/n254 ), .CK(CLK), .RN(\CU_I/n25 ), .QN(
        \CU_I/n27 ) );
  CLKBUF_X1 \dp/U764  ( .A(\dp/n69 ), .Z(\dp/n76 ) );
  CLKBUF_X1 \dp/U763  ( .A(\dp/n56 ), .Z(\dp/n70 ) );
  CLKBUF_X1 \dp/U762  ( .A(\dp/n132 ), .Z(\dp/n42 ) );
  CLKBUF_X1 \dp/U761  ( .A(\dp/n132 ), .Z(\dp/n41 ) );
  CLKBUF_X1 \dp/U760  ( .A(\dp/n132 ), .Z(\dp/n40 ) );
  CLKBUF_X1 \dp/U759  ( .A(\dp/n132 ), .Z(\dp/n39 ) );
  INV_X1 \dp/U758  ( .A(mem_in_en_i), .ZN(\dp/n632 ) );
  INV_X1 \dp/U757  ( .A(DRAM_DATA[0]), .ZN(\dp/n400 ) );
  INV_X1 \dp/U756  ( .A(DRAM_DATA[1]), .ZN(\dp/n365 ) );
  INV_X1 \dp/U755  ( .A(DRAM_DATA[2]), .ZN(\dp/n364 ) );
  INV_X1 \dp/U754  ( .A(DRAM_DATA[3]), .ZN(\dp/n363 ) );
  INV_X1 \dp/U752  ( .A(DRAM_DATA[4]), .ZN(\dp/n362 ) );
  INV_X1 \dp/U751  ( .A(DRAM_DATA[5]), .ZN(\dp/n361 ) );
  INV_X1 \dp/U750  ( .A(DRAM_DATA[6]), .ZN(\dp/n360 ) );
  INV_X1 \dp/U749  ( .A(DRAM_DATA[7]), .ZN(\dp/n359 ) );
  INV_X1 \dp/U748  ( .A(DRAM_DATA[8]), .ZN(\dp/n358 ) );
  INV_X1 \dp/U747  ( .A(DRAM_DATA[9]), .ZN(\dp/n357 ) );
  INV_X1 \dp/U746  ( .A(DRAM_DATA[10]), .ZN(\dp/n356 ) );
  INV_X1 \dp/U745  ( .A(DRAM_DATA[11]), .ZN(\dp/n355 ) );
  INV_X1 \dp/U744  ( .A(DRAM_DATA[12]), .ZN(\dp/n354 ) );
  INV_X1 \dp/U743  ( .A(DRAM_DATA[13]), .ZN(\dp/n353 ) );
  INV_X1 \dp/U742  ( .A(DRAM_DATA[14]), .ZN(\dp/n352 ) );
  INV_X1 \dp/U741  ( .A(DRAM_DATA[15]), .ZN(\dp/n351 ) );
  INV_X1 \dp/U740  ( .A(DRAM_DATA[16]), .ZN(\dp/n350 ) );
  INV_X1 \dp/U739  ( .A(DRAM_DATA[17]), .ZN(\dp/n349 ) );
  INV_X1 \dp/U738  ( .A(DRAM_DATA[18]), .ZN(\dp/n348 ) );
  INV_X1 \dp/U737  ( .A(DRAM_DATA[19]), .ZN(\dp/n347 ) );
  INV_X1 \dp/U736  ( .A(DRAM_DATA[20]), .ZN(\dp/n346 ) );
  INV_X1 \dp/U735  ( .A(DRAM_DATA[21]), .ZN(\dp/n345 ) );
  INV_X1 \dp/U734  ( .A(DRAM_DATA[22]), .ZN(\dp/n344 ) );
  INV_X1 \dp/U733  ( .A(DRAM_DATA[23]), .ZN(\dp/n343 ) );
  INV_X1 \dp/U732  ( .A(DRAM_DATA[24]), .ZN(\dp/n342 ) );
  INV_X1 \dp/U731  ( .A(DRAM_DATA[25]), .ZN(\dp/n341 ) );
  INV_X1 \dp/U730  ( .A(DRAM_DATA[26]), .ZN(\dp/n340 ) );
  INV_X1 \dp/U729  ( .A(DRAM_DATA[27]), .ZN(\dp/n339 ) );
  INV_X1 \dp/U728  ( .A(DRAM_DATA[28]), .ZN(\dp/n338 ) );
  INV_X1 \dp/U727  ( .A(DRAM_DATA[29]), .ZN(\dp/n337 ) );
  INV_X1 \dp/U726  ( .A(DRAM_DATA[30]), .ZN(\dp/n336 ) );
  INV_X1 \dp/U725  ( .A(DRAM_DATA[31]), .ZN(\dp/n335 ) );
  OAI22_X1 \dp/U724  ( .A1(\dp/n444 ), .A2(\dp/n59 ), .B1(\dp/n48 ), .B2(
        \dp/n597 ), .ZN(\dp/n774 ) );
  OAI22_X1 \dp/U723  ( .A1(\dp/n445 ), .A2(\dp/n59 ), .B1(\dp/n48 ), .B2(
        \dp/n596 ), .ZN(\dp/n775 ) );
  OAI22_X1 \dp/U722  ( .A1(\dp/n446 ), .A2(\dp/n58 ), .B1(\dp/n48 ), .B2(
        \dp/n597 ), .ZN(\dp/n776 ) );
  OAI22_X1 \dp/U721  ( .A1(\dp/n447 ), .A2(\dp/n59 ), .B1(\dp/n48 ), .B2(
        \dp/n597 ), .ZN(\dp/n777 ) );
  INV_X1 \dp/U720  ( .A(\dp/imm_id_o [31]), .ZN(\dp/n596 ) );
  OAI22_X1 \dp/U719  ( .A1(\dp/n448 ), .A2(\dp/n57 ), .B1(\dp/n49 ), .B2(
        \dp/n596 ), .ZN(\dp/n778 ) );
  OAI22_X1 \dp/U718  ( .A1(\dp/n449 ), .A2(\dp/n58 ), .B1(\dp/n49 ), .B2(
        \dp/n596 ), .ZN(\dp/n779 ) );
  INV_X1 \dp/U717  ( .A(\dp/imm_id_o [31]), .ZN(\dp/n597 ) );
  OAI22_X1 \dp/U716  ( .A1(\dp/n450 ), .A2(\dp/n58 ), .B1(\dp/n49 ), .B2(
        \dp/n597 ), .ZN(\dp/n780 ) );
  OAI221_X1 \dp/U715  ( .B1(\dp/n575 ), .B2(regrd_sel_i), .C1(\dp/n574 ), .C2(
        \dp/n633 ), .A(\dp/n631 ), .ZN(\dp/rd_fwd_id_o [0]) );
  INV_X1 \dp/U714  ( .A(\dp/rd_fwd_id_o [0]), .ZN(\dp/n412 ) );
  OAI22_X1 \dp/U713  ( .A1(\dp/n59 ), .A2(\dp/n414 ), .B1(\dp/n43 ), .B2(
        \dp/n412 ), .ZN(\dp/n712 ) );
  OAI221_X1 \dp/U712  ( .B1(\dp/n577 ), .B2(regrd_sel_i), .C1(\dp/n576 ), .C2(
        \dp/n633 ), .A(\dp/n631 ), .ZN(\dp/rd_fwd_id_o [1]) );
  INV_X1 \dp/U711  ( .A(\dp/rd_fwd_id_o [1]), .ZN(\dp/n517 ) );
  OAI22_X1 \dp/U710  ( .A1(\dp/n70 ), .A2(\dp/n415 ), .B1(\dp/n43 ), .B2(
        \dp/n517 ), .ZN(\dp/n713 ) );
  OAI221_X1 \dp/U709  ( .B1(\dp/n579 ), .B2(regrd_sel_i), .C1(\dp/n578 ), .C2(
        \dp/n633 ), .A(\dp/n631 ), .ZN(\dp/rd_fwd_id_o [2]) );
  INV_X1 \dp/U708  ( .A(\dp/rd_fwd_id_o [2]), .ZN(\dp/n521 ) );
  OAI22_X1 \dp/U707  ( .A1(\dp/n70 ), .A2(\dp/n416 ), .B1(\dp/n43 ), .B2(
        \dp/n521 ), .ZN(\dp/n714 ) );
  OAI221_X1 \dp/U706  ( .B1(\dp/n581 ), .B2(regrd_sel_i), .C1(\dp/n580 ), .C2(
        \dp/n633 ), .A(\dp/n631 ), .ZN(\dp/rd_fwd_id_o [3]) );
  INV_X1 \dp/U705  ( .A(\dp/rd_fwd_id_o [3]), .ZN(\dp/n525 ) );
  OAI22_X1 \dp/U704  ( .A1(\dp/n67 ), .A2(\dp/n417 ), .B1(\dp/n43 ), .B2(
        \dp/n525 ), .ZN(\dp/n715 ) );
  OAI221_X1 \dp/U703  ( .B1(\dp/n583 ), .B2(regrd_sel_i), .C1(\dp/n582 ), .C2(
        \dp/n633 ), .A(\dp/n631 ), .ZN(\dp/rd_fwd_id_o [4]) );
  INV_X1 \dp/U702  ( .A(\dp/rd_fwd_id_o [4]), .ZN(\dp/n585 ) );
  OAI22_X1 \dp/U701  ( .A1(\dp/n67 ), .A2(\dp/n418 ), .B1(\dp/n43 ), .B2(
        \dp/n585 ), .ZN(\dp/n716 ) );
  INV_X1 \dp/U700  ( .A(\dp/npc_id_o [0]), .ZN(\dp/n598 ) );
  OAI22_X1 \dp/U699  ( .A1(\dp/n67 ), .A2(\dp/n230 ), .B1(\dp/n43 ), .B2(
        \dp/n598 ), .ZN(\dp/n717 ) );
  INV_X1 \dp/U698  ( .A(\dp/npc_id_o [1]), .ZN(\dp/n599 ) );
  OAI22_X1 \dp/U697  ( .A1(\dp/n67 ), .A2(\dp/n231 ), .B1(\dp/n43 ), .B2(
        \dp/n599 ), .ZN(\dp/n718 ) );
  INV_X1 \dp/U696  ( .A(\dp/npc_id_o [2]), .ZN(\dp/n600 ) );
  OAI22_X1 \dp/U695  ( .A1(\dp/n67 ), .A2(\dp/n232 ), .B1(\dp/n43 ), .B2(
        \dp/n600 ), .ZN(\dp/n719 ) );
  INV_X1 \dp/U694  ( .A(\dp/npc_id_o [3]), .ZN(\dp/n601 ) );
  OAI22_X1 \dp/U693  ( .A1(\dp/n67 ), .A2(\dp/n233 ), .B1(\dp/n43 ), .B2(
        \dp/n601 ), .ZN(\dp/n720 ) );
  INV_X1 \dp/U692  ( .A(\dp/npc_id_o [4]), .ZN(\dp/n602 ) );
  OAI22_X1 \dp/U691  ( .A1(\dp/n67 ), .A2(\dp/n234 ), .B1(\dp/n43 ), .B2(
        \dp/n602 ), .ZN(\dp/n721 ) );
  INV_X1 \dp/U690  ( .A(\dp/npc_id_o [5]), .ZN(\dp/n603 ) );
  OAI22_X1 \dp/U689  ( .A1(\dp/n67 ), .A2(\dp/n235 ), .B1(\dp/n43 ), .B2(
        \dp/n603 ), .ZN(\dp/n722 ) );
  INV_X1 \dp/U688  ( .A(\dp/npc_id_o [6]), .ZN(\dp/n604 ) );
  OAI22_X1 \dp/U687  ( .A1(\dp/n67 ), .A2(\dp/n236 ), .B1(\dp/n44 ), .B2(
        \dp/n604 ), .ZN(\dp/n723 ) );
  INV_X1 \dp/U686  ( .A(\dp/npc_id_o [7]), .ZN(\dp/n605 ) );
  OAI22_X1 \dp/U685  ( .A1(\dp/n67 ), .A2(\dp/n237 ), .B1(\dp/n44 ), .B2(
        \dp/n605 ), .ZN(\dp/n724 ) );
  INV_X1 \dp/U684  ( .A(\dp/npc_id_o [8]), .ZN(\dp/n606 ) );
  OAI22_X1 \dp/U683  ( .A1(\dp/n67 ), .A2(\dp/n238 ), .B1(\dp/n44 ), .B2(
        \dp/n606 ), .ZN(\dp/n725 ) );
  INV_X1 \dp/U682  ( .A(\dp/npc_id_o [9]), .ZN(\dp/n607 ) );
  OAI22_X1 \dp/U681  ( .A1(\dp/n67 ), .A2(\dp/n239 ), .B1(\dp/n44 ), .B2(
        \dp/n607 ), .ZN(\dp/n726 ) );
  INV_X1 \dp/U680  ( .A(\dp/npc_id_o [10]), .ZN(\dp/n608 ) );
  OAI22_X1 \dp/U679  ( .A1(\dp/n66 ), .A2(\dp/n240 ), .B1(\dp/n44 ), .B2(
        \dp/n608 ), .ZN(\dp/n727 ) );
  INV_X1 \dp/U678  ( .A(\dp/npc_id_o [11]), .ZN(\dp/n609 ) );
  OAI22_X1 \dp/U677  ( .A1(\dp/n66 ), .A2(\dp/n241 ), .B1(\dp/n44 ), .B2(
        \dp/n609 ), .ZN(\dp/n728 ) );
  INV_X1 \dp/U676  ( .A(\dp/npc_id_o [12]), .ZN(\dp/n610 ) );
  OAI22_X1 \dp/U675  ( .A1(\dp/n66 ), .A2(\dp/n242 ), .B1(\dp/n44 ), .B2(
        \dp/n610 ), .ZN(\dp/n729 ) );
  INV_X1 \dp/U674  ( .A(\dp/npc_id_o [13]), .ZN(\dp/n611 ) );
  OAI22_X1 \dp/U673  ( .A1(\dp/n66 ), .A2(\dp/n243 ), .B1(\dp/n44 ), .B2(
        \dp/n611 ), .ZN(\dp/n730 ) );
  INV_X1 \dp/U672  ( .A(\dp/npc_id_o [14]), .ZN(\dp/n612 ) );
  OAI22_X1 \dp/U671  ( .A1(\dp/n66 ), .A2(\dp/n244 ), .B1(\dp/n44 ), .B2(
        \dp/n612 ), .ZN(\dp/n731 ) );
  INV_X1 \dp/U670  ( .A(\dp/npc_id_o [15]), .ZN(\dp/n613 ) );
  OAI22_X1 \dp/U669  ( .A1(\dp/n66 ), .A2(\dp/n245 ), .B1(\dp/n44 ), .B2(
        \dp/n613 ), .ZN(\dp/n732 ) );
  INV_X1 \dp/U668  ( .A(\dp/npc_id_o [16]), .ZN(\dp/n614 ) );
  OAI22_X1 \dp/U667  ( .A1(\dp/n66 ), .A2(\dp/n246 ), .B1(\dp/n44 ), .B2(
        \dp/n614 ), .ZN(\dp/n733 ) );
  INV_X1 \dp/U666  ( .A(\dp/npc_id_o [17]), .ZN(\dp/n615 ) );
  OAI22_X1 \dp/U665  ( .A1(\dp/n66 ), .A2(\dp/n247 ), .B1(\dp/n45 ), .B2(
        \dp/n615 ), .ZN(\dp/n734 ) );
  INV_X1 \dp/U664  ( .A(\dp/npc_id_o [18]), .ZN(\dp/n616 ) );
  OAI22_X1 \dp/U663  ( .A1(\dp/n66 ), .A2(\dp/n248 ), .B1(\dp/n45 ), .B2(
        \dp/n616 ), .ZN(\dp/n735 ) );
  INV_X1 \dp/U662  ( .A(\dp/npc_id_o [19]), .ZN(\dp/n617 ) );
  OAI22_X1 \dp/U661  ( .A1(\dp/n66 ), .A2(\dp/n249 ), .B1(\dp/n45 ), .B2(
        \dp/n617 ), .ZN(\dp/n736 ) );
  INV_X1 \dp/U660  ( .A(\dp/npc_id_o [20]), .ZN(\dp/n618 ) );
  OAI22_X1 \dp/U659  ( .A1(\dp/n66 ), .A2(\dp/n250 ), .B1(\dp/n45 ), .B2(
        \dp/n618 ), .ZN(\dp/n737 ) );
  INV_X1 \dp/U658  ( .A(\dp/npc_id_o [21]), .ZN(\dp/n619 ) );
  OAI22_X1 \dp/U657  ( .A1(\dp/n66 ), .A2(\dp/n251 ), .B1(\dp/n45 ), .B2(
        \dp/n619 ), .ZN(\dp/n738 ) );
  INV_X1 \dp/U656  ( .A(\dp/npc_id_o [22]), .ZN(\dp/n620 ) );
  OAI22_X1 \dp/U655  ( .A1(\dp/n65 ), .A2(\dp/n252 ), .B1(\dp/n45 ), .B2(
        \dp/n620 ), .ZN(\dp/n739 ) );
  INV_X1 \dp/U654  ( .A(\dp/npc_id_o [23]), .ZN(\dp/n621 ) );
  OAI22_X1 \dp/U653  ( .A1(\dp/n65 ), .A2(\dp/n253 ), .B1(\dp/n45 ), .B2(
        \dp/n621 ), .ZN(\dp/n740 ) );
  INV_X1 \dp/U652  ( .A(\dp/npc_id_o [24]), .ZN(\dp/n622 ) );
  OAI22_X1 \dp/U651  ( .A1(\dp/n65 ), .A2(\dp/n254 ), .B1(\dp/n45 ), .B2(
        \dp/n622 ), .ZN(\dp/n741 ) );
  INV_X1 \dp/U650  ( .A(\dp/npc_id_o [25]), .ZN(\dp/n623 ) );
  OAI22_X1 \dp/U649  ( .A1(\dp/n65 ), .A2(\dp/n255 ), .B1(\dp/n45 ), .B2(
        \dp/n623 ), .ZN(\dp/n742 ) );
  INV_X1 \dp/U648  ( .A(\dp/npc_id_o [26]), .ZN(\dp/n624 ) );
  OAI22_X1 \dp/U647  ( .A1(\dp/n65 ), .A2(\dp/n256 ), .B1(\dp/n45 ), .B2(
        \dp/n624 ), .ZN(\dp/n743 ) );
  INV_X1 \dp/U646  ( .A(\dp/npc_id_o [27]), .ZN(\dp/n625 ) );
  OAI22_X1 \dp/U645  ( .A1(\dp/n65 ), .A2(\dp/n257 ), .B1(\dp/n45 ), .B2(
        \dp/n625 ), .ZN(\dp/n744 ) );
  INV_X1 \dp/U644  ( .A(\dp/npc_id_o [28]), .ZN(\dp/n626 ) );
  OAI22_X1 \dp/U643  ( .A1(\dp/n65 ), .A2(\dp/n258 ), .B1(\dp/n46 ), .B2(
        \dp/n626 ), .ZN(\dp/n745 ) );
  INV_X1 \dp/U642  ( .A(\dp/npc_id_o [29]), .ZN(\dp/n627 ) );
  OAI22_X1 \dp/U641  ( .A1(\dp/n65 ), .A2(\dp/n259 ), .B1(\dp/n46 ), .B2(
        \dp/n627 ), .ZN(\dp/n746 ) );
  INV_X1 \dp/U640  ( .A(\dp/npc_id_o [30]), .ZN(\dp/n628 ) );
  OAI22_X1 \dp/U639  ( .A1(\dp/n65 ), .A2(\dp/n260 ), .B1(\dp/n46 ), .B2(
        \dp/n628 ), .ZN(\dp/n747 ) );
  INV_X1 \dp/U638  ( .A(\dp/npc_id_o [31]), .ZN(\dp/n629 ) );
  OAI22_X1 \dp/U637  ( .A1(\dp/n65 ), .A2(\dp/n261 ), .B1(\dp/n46 ), .B2(
        \dp/n629 ), .ZN(\dp/n748 ) );
  INV_X1 \dp/U636  ( .A(\dp/imm_id_o [19]), .ZN(\dp/n590 ) );
  OAI22_X1 \dp/U635  ( .A1(\dp/n438 ), .A2(\dp/n59 ), .B1(\dp/n48 ), .B2(
        \dp/n590 ), .ZN(\dp/n768 ) );
  INV_X1 \dp/U634  ( .A(\dp/imm_id_o [6]), .ZN(\dp/n407 ) );
  OAI22_X1 \dp/U633  ( .A1(\dp/n425 ), .A2(\dp/n57 ), .B1(\dp/n46 ), .B2(
        \dp/n407 ), .ZN(\dp/n755 ) );
  INV_X1 \dp/U632  ( .A(\dp/imm_id_o [7]), .ZN(\dp/n408 ) );
  OAI22_X1 \dp/U631  ( .A1(\dp/n426 ), .A2(\dp/n58 ), .B1(\dp/n47 ), .B2(
        \dp/n408 ), .ZN(\dp/n756 ) );
  INV_X1 \dp/U630  ( .A(\dp/imm_id_o [15]), .ZN(\dp/n586 ) );
  OAI22_X1 \dp/U629  ( .A1(\dp/n434 ), .A2(\dp/n57 ), .B1(\dp/n47 ), .B2(
        \dp/n586 ), .ZN(\dp/n764 ) );
  INV_X1 \dp/U628  ( .A(\dp/imm_id_o [16]), .ZN(\dp/n587 ) );
  OAI22_X1 \dp/U627  ( .A1(\dp/n435 ), .A2(\dp/n59 ), .B1(\dp/n47 ), .B2(
        \dp/n587 ), .ZN(\dp/n765 ) );
  INV_X1 \dp/U626  ( .A(\dp/imm_id_o [17]), .ZN(\dp/n588 ) );
  OAI22_X1 \dp/U625  ( .A1(\dp/n436 ), .A2(\dp/n57 ), .B1(\dp/n47 ), .B2(
        \dp/n588 ), .ZN(\dp/n766 ) );
  INV_X1 \dp/U624  ( .A(\dp/imm_id_o [18]), .ZN(\dp/n589 ) );
  OAI22_X1 \dp/U623  ( .A1(\dp/n437 ), .A2(\dp/n58 ), .B1(\dp/n48 ), .B2(
        \dp/n589 ), .ZN(\dp/n767 ) );
  INV_X1 \dp/U622  ( .A(\dp/imm_id_o [20]), .ZN(\dp/n591 ) );
  OAI22_X1 \dp/U621  ( .A1(\dp/n439 ), .A2(\dp/n59 ), .B1(\dp/n48 ), .B2(
        \dp/n591 ), .ZN(\dp/n769 ) );
  INV_X1 \dp/U620  ( .A(\dp/imm_id_o [21]), .ZN(\dp/n592 ) );
  OAI22_X1 \dp/U619  ( .A1(\dp/n440 ), .A2(\dp/n58 ), .B1(\dp/n48 ), .B2(
        \dp/n592 ), .ZN(\dp/n770 ) );
  INV_X1 \dp/U618  ( .A(\dp/imm_id_o [22]), .ZN(\dp/n593 ) );
  OAI22_X1 \dp/U617  ( .A1(\dp/n441 ), .A2(\dp/n59 ), .B1(\dp/n48 ), .B2(
        \dp/n593 ), .ZN(\dp/n771 ) );
  INV_X1 \dp/U616  ( .A(\dp/imm_id_o [23]), .ZN(\dp/n594 ) );
  OAI22_X1 \dp/U615  ( .A1(\dp/n442 ), .A2(\dp/n59 ), .B1(\dp/n48 ), .B2(
        \dp/n594 ), .ZN(\dp/n772 ) );
  INV_X1 \dp/U614  ( .A(\dp/imm_id_o [24]), .ZN(\dp/n595 ) );
  OAI22_X1 \dp/U613  ( .A1(\dp/n443 ), .A2(\dp/n58 ), .B1(\dp/n48 ), .B2(
        \dp/n595 ), .ZN(\dp/n773 ) );
  INV_X1 \dp/U612  ( .A(\dp/imm_id_o [0]), .ZN(\dp/n334 ) );
  OAI22_X1 \dp/U611  ( .A1(\dp/n419 ), .A2(\dp/n57 ), .B1(\dp/n46 ), .B2(
        \dp/n334 ), .ZN(\dp/n749 ) );
  INV_X1 \dp/U610  ( .A(\dp/imm_id_o [1]), .ZN(\dp/n402 ) );
  OAI22_X1 \dp/U609  ( .A1(\dp/n420 ), .A2(\dp/n58 ), .B1(\dp/n46 ), .B2(
        \dp/n402 ), .ZN(\dp/n750 ) );
  INV_X1 \dp/U608  ( .A(\dp/imm_id_o [2]), .ZN(\dp/n403 ) );
  OAI22_X1 \dp/U607  ( .A1(\dp/n421 ), .A2(\dp/n58 ), .B1(\dp/n46 ), .B2(
        \dp/n403 ), .ZN(\dp/n751 ) );
  INV_X1 \dp/U606  ( .A(\dp/imm_id_o [3]), .ZN(\dp/n404 ) );
  OAI22_X1 \dp/U605  ( .A1(\dp/n422 ), .A2(\dp/n57 ), .B1(\dp/n46 ), .B2(
        \dp/n404 ), .ZN(\dp/n752 ) );
  INV_X1 \dp/U604  ( .A(\dp/imm_id_o [4]), .ZN(\dp/n405 ) );
  OAI22_X1 \dp/U603  ( .A1(\dp/n423 ), .A2(\dp/n58 ), .B1(\dp/n46 ), .B2(
        \dp/n405 ), .ZN(\dp/n753 ) );
  INV_X1 \dp/U602  ( .A(\dp/imm_id_o [5]), .ZN(\dp/n406 ) );
  OAI22_X1 \dp/U601  ( .A1(\dp/n424 ), .A2(\dp/n58 ), .B1(\dp/n46 ), .B2(
        \dp/n406 ), .ZN(\dp/n754 ) );
  INV_X1 \dp/U600  ( .A(\dp/imm_id_o [8]), .ZN(\dp/n409 ) );
  OAI22_X1 \dp/U599  ( .A1(\dp/n427 ), .A2(\dp/n57 ), .B1(\dp/n47 ), .B2(
        \dp/n409 ), .ZN(\dp/n757 ) );
  INV_X1 \dp/U598  ( .A(\dp/imm_id_o [9]), .ZN(\dp/n410 ) );
  OAI22_X1 \dp/U597  ( .A1(\dp/n428 ), .A2(\dp/n57 ), .B1(\dp/n47 ), .B2(
        \dp/n410 ), .ZN(\dp/n758 ) );
  INV_X1 \dp/U596  ( .A(\dp/imm_id_o [10]), .ZN(\dp/n411 ) );
  OAI22_X1 \dp/U595  ( .A1(\dp/n429 ), .A2(\dp/n57 ), .B1(\dp/n47 ), .B2(
        \dp/n411 ), .ZN(\dp/n759 ) );
  INV_X1 \dp/U594  ( .A(\dp/imm_id_o [11]), .ZN(\dp/n413 ) );
  OAI22_X1 \dp/U593  ( .A1(\dp/n430 ), .A2(\dp/n58 ), .B1(\dp/n47 ), .B2(
        \dp/n413 ), .ZN(\dp/n760 ) );
  INV_X1 \dp/U592  ( .A(\dp/imm_id_o [12]), .ZN(\dp/n519 ) );
  OAI22_X1 \dp/U591  ( .A1(\dp/n431 ), .A2(\dp/n57 ), .B1(\dp/n47 ), .B2(
        \dp/n519 ), .ZN(\dp/n761 ) );
  INV_X1 \dp/U590  ( .A(\dp/imm_id_o [13]), .ZN(\dp/n523 ) );
  OAI22_X1 \dp/U589  ( .A1(\dp/n432 ), .A2(\dp/n57 ), .B1(\dp/n47 ), .B2(
        \dp/n523 ), .ZN(\dp/n762 ) );
  INV_X1 \dp/U588  ( .A(\dp/imm_id_o [14]), .ZN(\dp/n584 ) );
  OAI22_X1 \dp/U587  ( .A1(\dp/n433 ), .A2(\dp/n59 ), .B1(\dp/n47 ), .B2(
        \dp/n584 ), .ZN(\dp/n763 ) );
  INV_X1 \dp/U586  ( .A(\dp/rf_out2_id_o [0]), .ZN(\dp/n221 ) );
  OAI22_X1 \dp/U585  ( .A1(\dp/n65 ), .A2(\dp/n451 ), .B1(\dp/n49 ), .B2(
        \dp/n221 ), .ZN(\dp/n781 ) );
  INV_X1 \dp/U584  ( .A(\dp/rf_out2_id_o [1]), .ZN(\dp/n219 ) );
  OAI22_X1 \dp/U583  ( .A1(\dp/n65 ), .A2(\dp/n452 ), .B1(\dp/n49 ), .B2(
        \dp/n219 ), .ZN(\dp/n782 ) );
  INV_X1 \dp/U582  ( .A(\dp/rf_out2_id_o [2]), .ZN(\dp/n217 ) );
  OAI22_X1 \dp/U581  ( .A1(\dp/n64 ), .A2(\dp/n453 ), .B1(\dp/n49 ), .B2(
        \dp/n217 ), .ZN(\dp/n783 ) );
  INV_X1 \dp/U580  ( .A(\dp/rf_out2_id_o [3]), .ZN(\dp/n215 ) );
  OAI22_X1 \dp/U579  ( .A1(\dp/n64 ), .A2(\dp/n454 ), .B1(\dp/n49 ), .B2(
        \dp/n215 ), .ZN(\dp/n784 ) );
  INV_X1 \dp/U578  ( .A(\dp/rf_out2_id_o [4]), .ZN(\dp/n213 ) );
  OAI22_X1 \dp/U577  ( .A1(\dp/n64 ), .A2(\dp/n455 ), .B1(\dp/n49 ), .B2(
        \dp/n213 ), .ZN(\dp/n785 ) );
  INV_X1 \dp/U576  ( .A(\dp/rf_out2_id_o [5]), .ZN(\dp/n211 ) );
  OAI22_X1 \dp/U575  ( .A1(\dp/n64 ), .A2(\dp/n456 ), .B1(\dp/n49 ), .B2(
        \dp/n211 ), .ZN(\dp/n786 ) );
  INV_X1 \dp/U574  ( .A(\dp/rf_out2_id_o [6]), .ZN(\dp/n209 ) );
  OAI22_X1 \dp/U573  ( .A1(\dp/n64 ), .A2(\dp/n457 ), .B1(\dp/n49 ), .B2(
        \dp/n209 ), .ZN(\dp/n787 ) );
  INV_X1 \dp/U572  ( .A(\dp/rf_out2_id_o [7]), .ZN(\dp/n207 ) );
  OAI22_X1 \dp/U571  ( .A1(\dp/n64 ), .A2(\dp/n458 ), .B1(\dp/n49 ), .B2(
        \dp/n207 ), .ZN(\dp/n788 ) );
  INV_X1 \dp/U570  ( .A(\dp/rf_out2_id_o [8]), .ZN(\dp/n205 ) );
  OAI22_X1 \dp/U569  ( .A1(\dp/n64 ), .A2(\dp/n459 ), .B1(\dp/n50 ), .B2(
        \dp/n205 ), .ZN(\dp/n789 ) );
  INV_X1 \dp/U568  ( .A(\dp/rf_out2_id_o [9]), .ZN(\dp/n203 ) );
  OAI22_X1 \dp/U567  ( .A1(\dp/n64 ), .A2(\dp/n460 ), .B1(\dp/n50 ), .B2(
        \dp/n203 ), .ZN(\dp/n790 ) );
  INV_X1 \dp/U566  ( .A(\dp/rf_out2_id_o [10]), .ZN(\dp/n201 ) );
  OAI22_X1 \dp/U565  ( .A1(\dp/n64 ), .A2(\dp/n461 ), .B1(\dp/n50 ), .B2(
        \dp/n201 ), .ZN(\dp/n791 ) );
  INV_X1 \dp/U564  ( .A(\dp/rf_out2_id_o [11]), .ZN(\dp/n199 ) );
  OAI22_X1 \dp/U563  ( .A1(\dp/n64 ), .A2(\dp/n462 ), .B1(\dp/n50 ), .B2(
        \dp/n199 ), .ZN(\dp/n792 ) );
  INV_X1 \dp/U562  ( .A(\dp/rf_out2_id_o [12]), .ZN(\dp/n197 ) );
  OAI22_X1 \dp/U561  ( .A1(\dp/n64 ), .A2(\dp/n463 ), .B1(\dp/n50 ), .B2(
        \dp/n197 ), .ZN(\dp/n793 ) );
  INV_X1 \dp/U560  ( .A(\dp/rf_out2_id_o [13]), .ZN(\dp/n195 ) );
  OAI22_X1 \dp/U559  ( .A1(\dp/n64 ), .A2(\dp/n464 ), .B1(\dp/n50 ), .B2(
        \dp/n195 ), .ZN(\dp/n794 ) );
  INV_X1 \dp/U558  ( .A(\dp/rf_out2_id_o [14]), .ZN(\dp/n193 ) );
  OAI22_X1 \dp/U557  ( .A1(\dp/n63 ), .A2(\dp/n465 ), .B1(\dp/n50 ), .B2(
        \dp/n193 ), .ZN(\dp/n795 ) );
  INV_X1 \dp/U556  ( .A(\dp/rf_out2_id_o [15]), .ZN(\dp/n191 ) );
  OAI22_X1 \dp/U555  ( .A1(\dp/n63 ), .A2(\dp/n466 ), .B1(\dp/n50 ), .B2(
        \dp/n191 ), .ZN(\dp/n796 ) );
  INV_X1 \dp/U554  ( .A(\dp/rf_out2_id_o [16]), .ZN(\dp/n189 ) );
  OAI22_X1 \dp/U553  ( .A1(\dp/n63 ), .A2(\dp/n467 ), .B1(\dp/n50 ), .B2(
        \dp/n189 ), .ZN(\dp/n797 ) );
  INV_X1 \dp/U552  ( .A(\dp/rf_out2_id_o [17]), .ZN(\dp/n187 ) );
  OAI22_X1 \dp/U551  ( .A1(\dp/n63 ), .A2(\dp/n468 ), .B1(\dp/n50 ), .B2(
        \dp/n187 ), .ZN(\dp/n798 ) );
  INV_X1 \dp/U550  ( .A(\dp/rf_out2_id_o [18]), .ZN(\dp/n185 ) );
  OAI22_X1 \dp/U549  ( .A1(\dp/n63 ), .A2(\dp/n469 ), .B1(\dp/n50 ), .B2(
        \dp/n185 ), .ZN(\dp/n799 ) );
  INV_X1 \dp/U548  ( .A(\dp/rf_out2_id_o [19]), .ZN(\dp/n183 ) );
  OAI22_X1 \dp/U547  ( .A1(\dp/n63 ), .A2(\dp/n470 ), .B1(\dp/n51 ), .B2(
        \dp/n183 ), .ZN(\dp/n800 ) );
  INV_X1 \dp/U546  ( .A(\dp/rf_out2_id_o [20]), .ZN(\dp/n181 ) );
  OAI22_X1 \dp/U545  ( .A1(\dp/n63 ), .A2(\dp/n471 ), .B1(\dp/n51 ), .B2(
        \dp/n181 ), .ZN(\dp/n801 ) );
  INV_X1 \dp/U544  ( .A(\dp/rf_out2_id_o [21]), .ZN(\dp/n179 ) );
  OAI22_X1 \dp/U543  ( .A1(\dp/n63 ), .A2(\dp/n472 ), .B1(\dp/n51 ), .B2(
        \dp/n179 ), .ZN(\dp/n802 ) );
  INV_X1 \dp/U542  ( .A(\dp/rf_out2_id_o [22]), .ZN(\dp/n177 ) );
  OAI22_X1 \dp/U541  ( .A1(\dp/n63 ), .A2(\dp/n473 ), .B1(\dp/n51 ), .B2(
        \dp/n177 ), .ZN(\dp/n803 ) );
  INV_X1 \dp/U540  ( .A(\dp/rf_out2_id_o [23]), .ZN(\dp/n175 ) );
  OAI22_X1 \dp/U539  ( .A1(\dp/n63 ), .A2(\dp/n474 ), .B1(\dp/n51 ), .B2(
        \dp/n175 ), .ZN(\dp/n804 ) );
  INV_X1 \dp/U538  ( .A(\dp/rf_out2_id_o [24]), .ZN(\dp/n173 ) );
  OAI22_X1 \dp/U537  ( .A1(\dp/n63 ), .A2(\dp/n475 ), .B1(\dp/n51 ), .B2(
        \dp/n173 ), .ZN(\dp/n805 ) );
  INV_X1 \dp/U536  ( .A(\dp/rf_out2_id_o [25]), .ZN(\dp/n171 ) );
  OAI22_X1 \dp/U535  ( .A1(\dp/n62 ), .A2(\dp/n476 ), .B1(\dp/n51 ), .B2(
        \dp/n171 ), .ZN(\dp/n806 ) );
  INV_X1 \dp/U534  ( .A(\dp/rf_out2_id_o [26]), .ZN(\dp/n169 ) );
  OAI22_X1 \dp/U533  ( .A1(\dp/n62 ), .A2(\dp/n477 ), .B1(\dp/n51 ), .B2(
        \dp/n169 ), .ZN(\dp/n807 ) );
  INV_X1 \dp/U532  ( .A(\dp/rf_out2_id_o [27]), .ZN(\dp/n167 ) );
  OAI22_X1 \dp/U531  ( .A1(\dp/n62 ), .A2(\dp/n478 ), .B1(\dp/n51 ), .B2(
        \dp/n167 ), .ZN(\dp/n808 ) );
  INV_X1 \dp/U530  ( .A(\dp/rf_out2_id_o [28]), .ZN(\dp/n165 ) );
  OAI22_X1 \dp/U529  ( .A1(\dp/n61 ), .A2(\dp/n479 ), .B1(\dp/n51 ), .B2(
        \dp/n165 ), .ZN(\dp/n809 ) );
  INV_X1 \dp/U528  ( .A(\dp/rf_out2_id_o [29]), .ZN(\dp/n163 ) );
  OAI22_X1 \dp/U527  ( .A1(\dp/n61 ), .A2(\dp/n480 ), .B1(\dp/n51 ), .B2(
        \dp/n163 ), .ZN(\dp/n810 ) );
  INV_X1 \dp/U526  ( .A(\dp/rf_out2_id_o [30]), .ZN(\dp/n161 ) );
  OAI22_X1 \dp/U525  ( .A1(\dp/n62 ), .A2(\dp/n481 ), .B1(\dp/n52 ), .B2(
        \dp/n161 ), .ZN(\dp/n811 ) );
  INV_X1 \dp/U524  ( .A(\dp/rf_out2_id_o [31]), .ZN(\dp/n159 ) );
  OAI22_X1 \dp/U523  ( .A1(\dp/n62 ), .A2(\dp/n482 ), .B1(\dp/n52 ), .B2(
        \dp/n159 ), .ZN(\dp/n812 ) );
  INV_X1 \dp/U522  ( .A(\dp/rf_out1_id_o [0]), .ZN(\dp/n222 ) );
  OAI22_X1 \dp/U521  ( .A1(\dp/n63 ), .A2(\dp/n483 ), .B1(\dp/n52 ), .B2(
        \dp/n222 ), .ZN(\dp/n813 ) );
  INV_X1 \dp/U520  ( .A(\dp/rf_out1_id_o [1]), .ZN(\dp/n220 ) );
  OAI22_X1 \dp/U519  ( .A1(\dp/n62 ), .A2(\dp/n484 ), .B1(\dp/n52 ), .B2(
        \dp/n220 ), .ZN(\dp/n814 ) );
  INV_X1 \dp/U518  ( .A(\dp/rf_out1_id_o [2]), .ZN(\dp/n218 ) );
  OAI22_X1 \dp/U517  ( .A1(\dp/n60 ), .A2(\dp/n485 ), .B1(\dp/n52 ), .B2(
        \dp/n218 ), .ZN(\dp/n815 ) );
  INV_X1 \dp/U516  ( .A(\dp/rf_out1_id_o [3]), .ZN(\dp/n216 ) );
  OAI22_X1 \dp/U515  ( .A1(\dp/n60 ), .A2(\dp/n486 ), .B1(\dp/n52 ), .B2(
        \dp/n216 ), .ZN(\dp/n816 ) );
  INV_X1 \dp/U514  ( .A(\dp/rf_out1_id_o [4]), .ZN(\dp/n214 ) );
  OAI22_X1 \dp/U513  ( .A1(\dp/n62 ), .A2(\dp/n487 ), .B1(\dp/n52 ), .B2(
        \dp/n214 ), .ZN(\dp/n817 ) );
  INV_X1 \dp/U512  ( .A(\dp/rf_out1_id_o [5]), .ZN(\dp/n212 ) );
  OAI22_X1 \dp/U511  ( .A1(\dp/n60 ), .A2(\dp/n488 ), .B1(\dp/n52 ), .B2(
        \dp/n212 ), .ZN(\dp/n818 ) );
  INV_X1 \dp/U510  ( .A(\dp/rf_out1_id_o [6]), .ZN(\dp/n210 ) );
  OAI22_X1 \dp/U509  ( .A1(\dp/n62 ), .A2(\dp/n489 ), .B1(\dp/n52 ), .B2(
        \dp/n210 ), .ZN(\dp/n819 ) );
  INV_X1 \dp/U508  ( .A(\dp/rf_out1_id_o [7]), .ZN(\dp/n208 ) );
  OAI22_X1 \dp/U507  ( .A1(\dp/n62 ), .A2(\dp/n490 ), .B1(\dp/n52 ), .B2(
        \dp/n208 ), .ZN(\dp/n820 ) );
  INV_X1 \dp/U506  ( .A(\dp/rf_out1_id_o [8]), .ZN(\dp/n206 ) );
  OAI22_X1 \dp/U505  ( .A1(\dp/n60 ), .A2(\dp/n491 ), .B1(\dp/n52 ), .B2(
        \dp/n206 ), .ZN(\dp/n821 ) );
  INV_X1 \dp/U504  ( .A(\dp/rf_out1_id_o [9]), .ZN(\dp/n204 ) );
  OAI22_X1 \dp/U503  ( .A1(\dp/n60 ), .A2(\dp/n492 ), .B1(\dp/n53 ), .B2(
        \dp/n204 ), .ZN(\dp/n822 ) );
  INV_X1 \dp/U502  ( .A(\dp/rf_out1_id_o [10]), .ZN(\dp/n202 ) );
  OAI22_X1 \dp/U501  ( .A1(\dp/n61 ), .A2(\dp/n493 ), .B1(\dp/n53 ), .B2(
        \dp/n202 ), .ZN(\dp/n823 ) );
  INV_X1 \dp/U500  ( .A(\dp/rf_out1_id_o [11]), .ZN(\dp/n200 ) );
  OAI22_X1 \dp/U499  ( .A1(\dp/n60 ), .A2(\dp/n494 ), .B1(\dp/n53 ), .B2(
        \dp/n200 ), .ZN(\dp/n824 ) );
  INV_X1 \dp/U498  ( .A(\dp/rf_out1_id_o [12]), .ZN(\dp/n198 ) );
  OAI22_X1 \dp/U497  ( .A1(\dp/n60 ), .A2(\dp/n495 ), .B1(\dp/n53 ), .B2(
        \dp/n198 ), .ZN(\dp/n825 ) );
  INV_X1 \dp/U496  ( .A(\dp/rf_out1_id_o [13]), .ZN(\dp/n196 ) );
  OAI22_X1 \dp/U495  ( .A1(\dp/n62 ), .A2(\dp/n496 ), .B1(\dp/n53 ), .B2(
        \dp/n196 ), .ZN(\dp/n826 ) );
  INV_X1 \dp/U494  ( .A(\dp/rf_out1_id_o [14]), .ZN(\dp/n194 ) );
  OAI22_X1 \dp/U493  ( .A1(\dp/n61 ), .A2(\dp/n497 ), .B1(\dp/n53 ), .B2(
        \dp/n194 ), .ZN(\dp/n827 ) );
  INV_X1 \dp/U492  ( .A(\dp/rf_out1_id_o [15]), .ZN(\dp/n192 ) );
  OAI22_X1 \dp/U491  ( .A1(\dp/n60 ), .A2(\dp/n498 ), .B1(\dp/n53 ), .B2(
        \dp/n192 ), .ZN(\dp/n828 ) );
  INV_X1 \dp/U490  ( .A(\dp/rf_out1_id_o [16]), .ZN(\dp/n190 ) );
  OAI22_X1 \dp/U489  ( .A1(\dp/n61 ), .A2(\dp/n499 ), .B1(\dp/n53 ), .B2(
        \dp/n190 ), .ZN(\dp/n829 ) );
  INV_X1 \dp/U488  ( .A(\dp/rf_out1_id_o [17]), .ZN(\dp/n188 ) );
  OAI22_X1 \dp/U487  ( .A1(\dp/n60 ), .A2(\dp/n500 ), .B1(\dp/n53 ), .B2(
        \dp/n188 ), .ZN(\dp/n830 ) );
  INV_X1 \dp/U486  ( .A(\dp/rf_out1_id_o [18]), .ZN(\dp/n186 ) );
  OAI22_X1 \dp/U485  ( .A1(\dp/n60 ), .A2(\dp/n501 ), .B1(\dp/n53 ), .B2(
        \dp/n186 ), .ZN(\dp/n831 ) );
  INV_X1 \dp/U484  ( .A(\dp/rf_out1_id_o [19]), .ZN(\dp/n184 ) );
  OAI22_X1 \dp/U483  ( .A1(\dp/n61 ), .A2(\dp/n502 ), .B1(\dp/n53 ), .B2(
        \dp/n184 ), .ZN(\dp/n832 ) );
  INV_X1 \dp/U482  ( .A(\dp/rf_out1_id_o [20]), .ZN(\dp/n182 ) );
  OAI22_X1 \dp/U481  ( .A1(\dp/n61 ), .A2(\dp/n503 ), .B1(\dp/n54 ), .B2(
        \dp/n182 ), .ZN(\dp/n833 ) );
  INV_X1 \dp/U480  ( .A(\dp/rf_out1_id_o [21]), .ZN(\dp/n180 ) );
  OAI22_X1 \dp/U479  ( .A1(\dp/n60 ), .A2(\dp/n504 ), .B1(\dp/n54 ), .B2(
        \dp/n180 ), .ZN(\dp/n834 ) );
  INV_X1 \dp/U478  ( .A(\dp/rf_out1_id_o [22]), .ZN(\dp/n178 ) );
  OAI22_X1 \dp/U477  ( .A1(\dp/n61 ), .A2(\dp/n505 ), .B1(\dp/n54 ), .B2(
        \dp/n178 ), .ZN(\dp/n835 ) );
  INV_X1 \dp/U476  ( .A(\dp/rf_out1_id_o [23]), .ZN(\dp/n176 ) );
  OAI22_X1 \dp/U475  ( .A1(\dp/n60 ), .A2(\dp/n506 ), .B1(\dp/n54 ), .B2(
        \dp/n176 ), .ZN(\dp/n836 ) );
  INV_X1 \dp/U474  ( .A(\dp/rf_out1_id_o [24]), .ZN(\dp/n174 ) );
  OAI22_X1 \dp/U473  ( .A1(\dp/n61 ), .A2(\dp/n507 ), .B1(\dp/n54 ), .B2(
        \dp/n174 ), .ZN(\dp/n837 ) );
  INV_X1 \dp/U472  ( .A(\dp/rf_out1_id_o [25]), .ZN(\dp/n172 ) );
  OAI22_X1 \dp/U471  ( .A1(\dp/n61 ), .A2(\dp/n508 ), .B1(\dp/n54 ), .B2(
        \dp/n172 ), .ZN(\dp/n838 ) );
  INV_X1 \dp/U470  ( .A(\dp/rf_out1_id_o [26]), .ZN(\dp/n170 ) );
  OAI22_X1 \dp/U469  ( .A1(\dp/n59 ), .A2(\dp/n509 ), .B1(\dp/n54 ), .B2(
        \dp/n170 ), .ZN(\dp/n839 ) );
  INV_X1 \dp/U468  ( .A(\dp/rf_out1_id_o [27]), .ZN(\dp/n168 ) );
  OAI22_X1 \dp/U467  ( .A1(\dp/n62 ), .A2(\dp/n510 ), .B1(\dp/n54 ), .B2(
        \dp/n168 ), .ZN(\dp/n840 ) );
  INV_X1 \dp/U466  ( .A(\dp/rf_out1_id_o [28]), .ZN(\dp/n166 ) );
  OAI22_X1 \dp/U465  ( .A1(\dp/n61 ), .A2(\dp/n511 ), .B1(\dp/n54 ), .B2(
        \dp/n166 ), .ZN(\dp/n841 ) );
  INV_X1 \dp/U464  ( .A(\dp/rf_out1_id_o [29]), .ZN(\dp/n164 ) );
  OAI22_X1 \dp/U463  ( .A1(\dp/n59 ), .A2(\dp/n512 ), .B1(\dp/n54 ), .B2(
        \dp/n164 ), .ZN(\dp/n842 ) );
  INV_X1 \dp/U462  ( .A(\dp/rf_out1_id_o [30]), .ZN(\dp/n162 ) );
  OAI22_X1 \dp/U461  ( .A1(\dp/n62 ), .A2(\dp/n513 ), .B1(\dp/n54 ), .B2(
        \dp/n162 ), .ZN(\dp/n843 ) );
  INV_X1 \dp/U460  ( .A(\dp/rf_out1_id_o [31]), .ZN(\dp/n160 ) );
  OAI22_X1 \dp/U459  ( .A1(\dp/n61 ), .A2(\dp/n514 ), .B1(\dp/n48 ), .B2(
        \dp/n160 ), .ZN(\dp/n844 ) );
  INV_X1 \dp/U458  ( .A(reg31_sel_i), .ZN(\dp/n631 ) );
  INV_X1 \dp/U457  ( .A(regrd_sel_i), .ZN(\dp/n633 ) );
  INV_X1 \dp/U456  ( .A(\dp/rd_fwd_ex_o [0]), .ZN(\dp/n225 ) );
  OAI22_X1 \dp/U455  ( .A1(\dp/n35 ), .A2(\dp/n264 ), .B1(\dp/n31 ), .B2(
        \dp/n225 ), .ZN(\dp/n1014 ) );
  INV_X1 \dp/U454  ( .A(\dp/branch_t_ex_o ), .ZN(\dp/n262 ) );
  OAI22_X1 \dp/U453  ( .A1(\dp/n515 ), .A2(\dp/n33 ), .B1(\dp/n31 ), .B2(
        \dp/n262 ), .ZN(\dp/n845 ) );
  INV_X1 \dp/U452  ( .A(\dp/rd_fwd_ex_o [1]), .ZN(\dp/n226 ) );
  OAI22_X1 \dp/U451  ( .A1(\dp/n35 ), .A2(\dp/n265 ), .B1(\dp/n31 ), .B2(
        \dp/n226 ), .ZN(\dp/n1013 ) );
  INV_X1 \dp/U450  ( .A(\dp/rd_fwd_ex_o [2]), .ZN(\dp/n227 ) );
  OAI22_X1 \dp/U449  ( .A1(\dp/n36 ), .A2(\dp/n266 ), .B1(\dp/n31 ), .B2(
        \dp/n227 ), .ZN(\dp/n1012 ) );
  INV_X1 \dp/U448  ( .A(\dp/rd_fwd_ex_o [3]), .ZN(\dp/n228 ) );
  OAI22_X1 \dp/U447  ( .A1(\dp/n36 ), .A2(\dp/n267 ), .B1(\dp/n31 ), .B2(
        \dp/n228 ), .ZN(\dp/n1011 ) );
  INV_X1 \dp/U446  ( .A(\dp/rd_fwd_ex_o [4]), .ZN(\dp/n229 ) );
  OAI22_X1 \dp/U445  ( .A1(\dp/n36 ), .A2(\dp/n268 ), .B1(\dp/n31 ), .B2(
        \dp/n229 ), .ZN(\dp/n1010 ) );
  OAI22_X1 \dp/U444  ( .A1(\dp/n30 ), .A2(\dp/n516 ), .B1(\dp/n24 ), .B2(
        \dp/n264 ), .ZN(\dp/n1009 ) );
  OAI22_X1 \dp/U443  ( .A1(\dp/n30 ), .A2(\dp/n518 ), .B1(\dp/n24 ), .B2(
        \dp/n265 ), .ZN(\dp/n1008 ) );
  OAI22_X1 \dp/U442  ( .A1(\dp/n30 ), .A2(\dp/n520 ), .B1(\dp/n24 ), .B2(
        \dp/n266 ), .ZN(\dp/n1007 ) );
  OAI22_X1 \dp/U441  ( .A1(\dp/n30 ), .A2(\dp/n522 ), .B1(\dp/n24 ), .B2(
        \dp/n267 ), .ZN(\dp/n1006 ) );
  OAI22_X1 \dp/U440  ( .A1(\dp/n30 ), .A2(\dp/n524 ), .B1(\dp/n24 ), .B2(
        \dp/n268 ), .ZN(\dp/n1005 ) );
  OAI22_X1 \dp/U439  ( .A1(\dp/n303 ), .A2(\dp/n27 ), .B1(\dp/n877 ), .B2(
        \dp/n21 ), .ZN(\dp/n909 ) );
  OAI22_X1 \dp/U438  ( .A1(\dp/n304 ), .A2(\dp/n27 ), .B1(\dp/n876 ), .B2(
        \dp/n21 ), .ZN(\dp/n908 ) );
  OAI22_X1 \dp/U437  ( .A1(\dp/n305 ), .A2(\dp/n28 ), .B1(\dp/n875 ), .B2(
        \dp/n21 ), .ZN(\dp/n907 ) );
  OAI22_X1 \dp/U436  ( .A1(\dp/n306 ), .A2(\dp/n28 ), .B1(\dp/n874 ), .B2(
        \dp/n21 ), .ZN(\dp/n906 ) );
  OAI22_X1 \dp/U435  ( .A1(\dp/n307 ), .A2(\dp/n28 ), .B1(\dp/n873 ), .B2(
        \dp/n21 ), .ZN(\dp/n905 ) );
  OAI22_X1 \dp/U434  ( .A1(\dp/n308 ), .A2(\dp/n28 ), .B1(\dp/n872 ), .B2(
        \dp/n21 ), .ZN(\dp/n904 ) );
  OAI22_X1 \dp/U433  ( .A1(\dp/n309 ), .A2(\dp/n28 ), .B1(\dp/n871 ), .B2(
        \dp/n21 ), .ZN(\dp/n903 ) );
  OAI22_X1 \dp/U432  ( .A1(\dp/n310 ), .A2(\dp/n28 ), .B1(\dp/n870 ), .B2(
        \dp/n21 ), .ZN(\dp/n902 ) );
  OAI22_X1 \dp/U431  ( .A1(\dp/n311 ), .A2(\dp/n28 ), .B1(\dp/n869 ), .B2(
        \dp/n20 ), .ZN(\dp/n901 ) );
  OAI22_X1 \dp/U430  ( .A1(\dp/n312 ), .A2(\dp/n28 ), .B1(\dp/n868 ), .B2(
        \dp/n20 ), .ZN(\dp/n900 ) );
  OAI22_X1 \dp/U429  ( .A1(\dp/n313 ), .A2(\dp/n28 ), .B1(\dp/n867 ), .B2(
        \dp/n20 ), .ZN(\dp/n899 ) );
  OAI22_X1 \dp/U428  ( .A1(\dp/n314 ), .A2(\dp/n28 ), .B1(\dp/n866 ), .B2(
        \dp/n20 ), .ZN(\dp/n898 ) );
  OAI22_X1 \dp/U427  ( .A1(\dp/n315 ), .A2(\dp/n28 ), .B1(\dp/n865 ), .B2(
        \dp/n20 ), .ZN(\dp/n897 ) );
  OAI22_X1 \dp/U426  ( .A1(\dp/n316 ), .A2(\dp/n28 ), .B1(\dp/n864 ), .B2(
        \dp/n20 ), .ZN(\dp/n896 ) );
  OAI22_X1 \dp/U425  ( .A1(\dp/n317 ), .A2(\dp/n29 ), .B1(\dp/n863 ), .B2(
        \dp/n20 ), .ZN(\dp/n895 ) );
  OAI22_X1 \dp/U424  ( .A1(\dp/n318 ), .A2(\dp/n29 ), .B1(\dp/n862 ), .B2(
        \dp/n20 ), .ZN(\dp/n894 ) );
  OAI22_X1 \dp/U423  ( .A1(\dp/n319 ), .A2(\dp/n29 ), .B1(\dp/n861 ), .B2(
        \dp/n20 ), .ZN(\dp/n893 ) );
  OAI22_X1 \dp/U422  ( .A1(\dp/n320 ), .A2(\dp/n29 ), .B1(\dp/n860 ), .B2(
        \dp/n20 ), .ZN(\dp/n892 ) );
  OAI22_X1 \dp/U421  ( .A1(\dp/n321 ), .A2(\dp/n29 ), .B1(\dp/n859 ), .B2(
        \dp/n20 ), .ZN(\dp/n891 ) );
  OAI22_X1 \dp/U420  ( .A1(\dp/n322 ), .A2(\dp/n29 ), .B1(\dp/n858 ), .B2(
        \dp/n20 ), .ZN(\dp/n890 ) );
  OAI22_X1 \dp/U419  ( .A1(\dp/n323 ), .A2(\dp/n29 ), .B1(\dp/n857 ), .B2(
        \dp/n19 ), .ZN(\dp/n889 ) );
  OAI22_X1 \dp/U418  ( .A1(\dp/n324 ), .A2(\dp/n29 ), .B1(\dp/n856 ), .B2(
        \dp/n19 ), .ZN(\dp/n888 ) );
  OAI22_X1 \dp/U417  ( .A1(\dp/n325 ), .A2(\dp/n29 ), .B1(\dp/n855 ), .B2(
        \dp/n19 ), .ZN(\dp/n887 ) );
  OAI22_X1 \dp/U416  ( .A1(\dp/n326 ), .A2(\dp/n29 ), .B1(\dp/n854 ), .B2(
        \dp/n19 ), .ZN(\dp/n886 ) );
  OAI22_X1 \dp/U415  ( .A1(\dp/n327 ), .A2(\dp/n29 ), .B1(\dp/n853 ), .B2(
        \dp/n19 ), .ZN(\dp/n885 ) );
  OAI22_X1 \dp/U414  ( .A1(\dp/n328 ), .A2(\dp/n29 ), .B1(\dp/n852 ), .B2(
        \dp/n19 ), .ZN(\dp/n884 ) );
  OAI22_X1 \dp/U413  ( .A1(\dp/n329 ), .A2(\dp/n30 ), .B1(\dp/n851 ), .B2(
        \dp/n19 ), .ZN(\dp/n883 ) );
  OAI22_X1 \dp/U412  ( .A1(\dp/n330 ), .A2(\dp/n30 ), .B1(\dp/n850 ), .B2(
        \dp/n19 ), .ZN(\dp/n882 ) );
  OAI22_X1 \dp/U411  ( .A1(\dp/n331 ), .A2(\dp/n30 ), .B1(\dp/n849 ), .B2(
        \dp/n19 ), .ZN(\dp/n881 ) );
  OAI22_X1 \dp/U410  ( .A1(\dp/n332 ), .A2(\dp/n30 ), .B1(\dp/n848 ), .B2(
        \dp/n19 ), .ZN(\dp/n880 ) );
  OAI22_X1 \dp/U409  ( .A1(\dp/n333 ), .A2(\dp/n30 ), .B1(\dp/n847 ), .B2(
        \dp/n19 ), .ZN(\dp/n879 ) );
  OAI22_X1 \dp/U408  ( .A1(\dp/n630 ), .A2(\dp/n25 ), .B1(\dp/n846 ), .B2(
        \dp/n19 ), .ZN(\dp/n878 ) );
  INV_X1 \dp/U407  ( .A(instr_i[0]), .ZN(\dp/n1027 ) );
  OAI22_X1 \dp/U406  ( .A1(\dp/n526 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1027 ), .ZN(\dp/n649 ) );
  INV_X1 \dp/U405  ( .A(instr_i[1]), .ZN(\dp/n1026 ) );
  OAI22_X1 \dp/U404  ( .A1(\dp/n527 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1026 ), .ZN(\dp/n650 ) );
  INV_X1 \dp/U403  ( .A(instr_i[2]), .ZN(\dp/n1025 ) );
  OAI22_X1 \dp/U402  ( .A1(\dp/n528 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1025 ), .ZN(\dp/n651 ) );
  INV_X1 \dp/U401  ( .A(instr_i[3]), .ZN(\dp/n1024 ) );
  OAI22_X1 \dp/U400  ( .A1(\dp/n529 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1024 ), .ZN(\dp/n652 ) );
  INV_X1 \dp/U399  ( .A(instr_i[4]), .ZN(\dp/n1023 ) );
  OAI22_X1 \dp/U398  ( .A1(\dp/n530 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1023 ), .ZN(\dp/n653 ) );
  INV_X1 \dp/U397  ( .A(instr_i[5]), .ZN(\dp/n1022 ) );
  OAI22_X1 \dp/U396  ( .A1(\dp/n531 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1022 ), .ZN(\dp/n654 ) );
  INV_X1 \dp/U395  ( .A(instr_i[6]), .ZN(\dp/n1021 ) );
  OAI22_X1 \dp/U394  ( .A1(\dp/n532 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1021 ), .ZN(\dp/n655 ) );
  INV_X1 \dp/U393  ( .A(instr_i[7]), .ZN(\dp/n1020 ) );
  OAI22_X1 \dp/U392  ( .A1(\dp/n533 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1020 ), .ZN(\dp/n656 ) );
  INV_X1 \dp/U391  ( .A(instr_i[8]), .ZN(\dp/n1019 ) );
  OAI22_X1 \dp/U390  ( .A1(\dp/n534 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1019 ), .ZN(\dp/n657 ) );
  INV_X1 \dp/U389  ( .A(instr_i[9]), .ZN(\dp/n1018 ) );
  OAI22_X1 \dp/U388  ( .A1(\dp/n535 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1018 ), .ZN(\dp/n658 ) );
  INV_X1 \dp/U387  ( .A(instr_i[10]), .ZN(\dp/n1017 ) );
  OAI22_X1 \dp/U386  ( .A1(\dp/n536 ), .A2(\dp/n79 ), .B1(\dp/n71 ), .B2(
        \dp/n1017 ), .ZN(\dp/n659 ) );
  INV_X1 \dp/U385  ( .A(instr_i[11]), .ZN(\dp/n1016 ) );
  OAI22_X1 \dp/U384  ( .A1(\dp/n575 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n1016 ), .ZN(\dp/n660 ) );
  INV_X1 \dp/U383  ( .A(instr_i[12]), .ZN(\dp/n648 ) );
  OAI22_X1 \dp/U382  ( .A1(\dp/n577 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n648 ), .ZN(\dp/n661 ) );
  INV_X1 \dp/U381  ( .A(instr_i[13]), .ZN(\dp/n647 ) );
  OAI22_X1 \dp/U380  ( .A1(\dp/n579 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n647 ), .ZN(\dp/n662 ) );
  INV_X1 \dp/U379  ( .A(instr_i[14]), .ZN(\dp/n646 ) );
  OAI22_X1 \dp/U378  ( .A1(\dp/n581 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n646 ), .ZN(\dp/n663 ) );
  INV_X1 \dp/U377  ( .A(instr_i[15]), .ZN(\dp/n645 ) );
  OAI22_X1 \dp/U376  ( .A1(\dp/n583 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n645 ), .ZN(\dp/n664 ) );
  INV_X1 \dp/U375  ( .A(instr_i[16]), .ZN(\dp/n644 ) );
  OAI22_X1 \dp/U374  ( .A1(\dp/n574 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n644 ), .ZN(\dp/n665 ) );
  INV_X1 \dp/U373  ( .A(instr_i[17]), .ZN(\dp/n643 ) );
  OAI22_X1 \dp/U372  ( .A1(\dp/n576 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n643 ), .ZN(\dp/n666 ) );
  INV_X1 \dp/U371  ( .A(instr_i[18]), .ZN(\dp/n642 ) );
  OAI22_X1 \dp/U370  ( .A1(\dp/n578 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n642 ), .ZN(\dp/n667 ) );
  INV_X1 \dp/U369  ( .A(instr_i[19]), .ZN(\dp/n641 ) );
  OAI22_X1 \dp/U368  ( .A1(\dp/n580 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n641 ), .ZN(\dp/n668 ) );
  INV_X1 \dp/U367  ( .A(instr_i[20]), .ZN(\dp/n640 ) );
  OAI22_X1 \dp/U366  ( .A1(\dp/n582 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n640 ), .ZN(\dp/n669 ) );
  INV_X1 \dp/U365  ( .A(instr_i[21]), .ZN(\dp/n639 ) );
  OAI22_X1 \dp/U364  ( .A1(\dp/n537 ), .A2(\dp/n80 ), .B1(\dp/n72 ), .B2(
        \dp/n639 ), .ZN(\dp/n670 ) );
  INV_X1 \dp/U363  ( .A(instr_i[22]), .ZN(\dp/n638 ) );
  OAI22_X1 \dp/U362  ( .A1(\dp/n538 ), .A2(\dp/n80 ), .B1(\dp/n73 ), .B2(
        \dp/n638 ), .ZN(\dp/n671 ) );
  INV_X1 \dp/U361  ( .A(instr_i[23]), .ZN(\dp/n637 ) );
  OAI22_X1 \dp/U360  ( .A1(\dp/n539 ), .A2(\dp/n81 ), .B1(\dp/n73 ), .B2(
        \dp/n637 ), .ZN(\dp/n672 ) );
  INV_X1 \dp/U359  ( .A(instr_i[24]), .ZN(\dp/n636 ) );
  OAI22_X1 \dp/U358  ( .A1(\dp/n540 ), .A2(\dp/n81 ), .B1(\dp/n73 ), .B2(
        \dp/n636 ), .ZN(\dp/n673 ) );
  INV_X1 \dp/U357  ( .A(instr_i[25]), .ZN(\dp/n635 ) );
  OAI22_X1 \dp/U356  ( .A1(\dp/n541 ), .A2(\dp/n81 ), .B1(\dp/n73 ), .B2(
        \dp/n635 ), .ZN(\dp/n674 ) );
  INV_X1 \dp/U355  ( .A(\dp/npc_if_o [0]), .ZN(\dp/n223 ) );
  OAI22_X1 \dp/U354  ( .A1(\dp/n81 ), .A2(\dp/n542 ), .B1(\dp/n73 ), .B2(
        \dp/n223 ), .ZN(\dp/n675 ) );
  INV_X1 \dp/U353  ( .A(\dp/npc_if_o [1]), .ZN(\dp/n124 ) );
  OAI22_X1 \dp/U352  ( .A1(\dp/n83 ), .A2(\dp/n543 ), .B1(\dp/n73 ), .B2(
        \dp/n124 ), .ZN(\dp/n676 ) );
  INV_X1 \dp/U351  ( .A(\dp/npc_if_o [2]), .ZN(\dp/n123 ) );
  OAI22_X1 \dp/U350  ( .A1(\dp/n83 ), .A2(\dp/n544 ), .B1(\dp/n73 ), .B2(
        \dp/n123 ), .ZN(\dp/n677 ) );
  INV_X1 \dp/U349  ( .A(\dp/npc_if_o [3]), .ZN(\dp/n122 ) );
  OAI22_X1 \dp/U348  ( .A1(\dp/n83 ), .A2(\dp/n545 ), .B1(\dp/n73 ), .B2(
        \dp/n122 ), .ZN(\dp/n678 ) );
  INV_X1 \dp/U347  ( .A(\dp/npc_if_o [4]), .ZN(\dp/n121 ) );
  OAI22_X1 \dp/U346  ( .A1(\dp/n83 ), .A2(\dp/n546 ), .B1(\dp/n73 ), .B2(
        \dp/n121 ), .ZN(\dp/n679 ) );
  INV_X1 \dp/U345  ( .A(\dp/npc_if_o [5]), .ZN(\dp/n120 ) );
  OAI22_X1 \dp/U344  ( .A1(\dp/n83 ), .A2(\dp/n547 ), .B1(\dp/n73 ), .B2(
        \dp/n120 ), .ZN(\dp/n680 ) );
  INV_X1 \dp/U343  ( .A(\dp/npc_if_o [6]), .ZN(\dp/n119 ) );
  OAI22_X1 \dp/U342  ( .A1(\dp/n83 ), .A2(\dp/n548 ), .B1(\dp/n73 ), .B2(
        \dp/n119 ), .ZN(\dp/n681 ) );
  INV_X1 \dp/U341  ( .A(\dp/npc_if_o [7]), .ZN(\dp/n118 ) );
  OAI22_X1 \dp/U340  ( .A1(\dp/n83 ), .A2(\dp/n549 ), .B1(\dp/n74 ), .B2(
        \dp/n118 ), .ZN(\dp/n682 ) );
  INV_X1 \dp/U339  ( .A(\dp/npc_if_o [8]), .ZN(\dp/n117 ) );
  OAI22_X1 \dp/U338  ( .A1(\dp/n83 ), .A2(\dp/n550 ), .B1(\dp/n74 ), .B2(
        \dp/n117 ), .ZN(\dp/n683 ) );
  INV_X1 \dp/U337  ( .A(\dp/alu_out_ex_o [28]), .ZN(\dp/n128 ) );
  OAI22_X1 \dp/U336  ( .A1(\dp/n849 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n128 ), .ZN(\dp/n913 ) );
  INV_X1 \dp/U335  ( .A(\dp/alu_out_ex_o [29]), .ZN(\dp/n127 ) );
  OAI22_X1 \dp/U334  ( .A1(\dp/n848 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n127 ), .ZN(\dp/n912 ) );
  INV_X1 \dp/U333  ( .A(\dp/alu_out_ex_o [30]), .ZN(\dp/n126 ) );
  OAI22_X1 \dp/U332  ( .A1(\dp/n847 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n126 ), .ZN(\dp/n911 ) );
  INV_X1 \dp/U331  ( .A(\dp/alu_out_ex_o [31]), .ZN(\dp/n125 ) );
  OAI22_X1 \dp/U330  ( .A1(\dp/n846 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n125 ), .ZN(\dp/n910 ) );
  INV_X1 \dp/U329  ( .A(\dp/alu_out_ex_o [5]), .ZN(\dp/n153 ) );
  OAI22_X1 \dp/U328  ( .A1(\dp/n872 ), .A2(\dp/n35 ), .B1(\dp/n31 ), .B2(
        \dp/n153 ), .ZN(\dp/n936 ) );
  INV_X1 \dp/U327  ( .A(\dp/alu_out_ex_o [6]), .ZN(\dp/n152 ) );
  OAI22_X1 \dp/U326  ( .A1(\dp/n871 ), .A2(\dp/n35 ), .B1(\dp/n31 ), .B2(
        \dp/n152 ), .ZN(\dp/n935 ) );
  INV_X1 \dp/U325  ( .A(\dp/alu_out_ex_o [7]), .ZN(\dp/n151 ) );
  OAI22_X1 \dp/U324  ( .A1(\dp/n870 ), .A2(\dp/n35 ), .B1(\dp/n31 ), .B2(
        \dp/n151 ), .ZN(\dp/n934 ) );
  INV_X1 \dp/U323  ( .A(\dp/alu_out_ex_o [8]), .ZN(\dp/n150 ) );
  OAI22_X1 \dp/U322  ( .A1(\dp/n869 ), .A2(\dp/n35 ), .B1(\dp/n32 ), .B2(
        \dp/n150 ), .ZN(\dp/n933 ) );
  INV_X1 \dp/U321  ( .A(\dp/alu_out_ex_o [9]), .ZN(\dp/n149 ) );
  OAI22_X1 \dp/U320  ( .A1(\dp/n868 ), .A2(\dp/n35 ), .B1(\dp/n32 ), .B2(
        \dp/n149 ), .ZN(\dp/n932 ) );
  INV_X1 \dp/U319  ( .A(\dp/alu_out_ex_o [12]), .ZN(\dp/n146 ) );
  OAI22_X1 \dp/U318  ( .A1(\dp/n865 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n146 ), .ZN(\dp/n929 ) );
  INV_X1 \dp/U317  ( .A(\dp/alu_out_ex_o [17]), .ZN(\dp/n141 ) );
  OAI22_X1 \dp/U316  ( .A1(\dp/n860 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n141 ), .ZN(\dp/n924 ) );
  INV_X1 \dp/U315  ( .A(\dp/alu_out_ex_o [18]), .ZN(\dp/n140 ) );
  OAI22_X1 \dp/U314  ( .A1(\dp/n859 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n140 ), .ZN(\dp/n923 ) );
  INV_X1 \dp/U313  ( .A(\dp/alu_out_ex_o [19]), .ZN(\dp/n139 ) );
  OAI22_X1 \dp/U312  ( .A1(\dp/n858 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n139 ), .ZN(\dp/n922 ) );
  INV_X1 \dp/U311  ( .A(\dp/alu_out_ex_o [20]), .ZN(\dp/n138 ) );
  OAI22_X1 \dp/U310  ( .A1(\dp/n857 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n138 ), .ZN(\dp/n921 ) );
  INV_X1 \dp/U309  ( .A(\dp/alu_out_ex_o [21]), .ZN(\dp/n137 ) );
  OAI22_X1 \dp/U308  ( .A1(\dp/n856 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n137 ), .ZN(\dp/n920 ) );
  INV_X1 \dp/U307  ( .A(\dp/alu_out_ex_o [22]), .ZN(\dp/n136 ) );
  OAI22_X1 \dp/U306  ( .A1(\dp/n855 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n136 ), .ZN(\dp/n919 ) );
  INV_X1 \dp/U305  ( .A(\dp/alu_out_ex_o [23]), .ZN(\dp/n135 ) );
  OAI22_X1 \dp/U304  ( .A1(\dp/n854 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n135 ), .ZN(\dp/n918 ) );
  INV_X1 \dp/U303  ( .A(\dp/alu_out_ex_o [24]), .ZN(\dp/n134 ) );
  OAI22_X1 \dp/U302  ( .A1(\dp/n853 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n134 ), .ZN(\dp/n917 ) );
  INV_X1 \dp/U301  ( .A(\dp/alu_out_ex_o [25]), .ZN(\dp/n133 ) );
  OAI22_X1 \dp/U300  ( .A1(\dp/n852 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n133 ), .ZN(\dp/n916 ) );
  INV_X1 \dp/U299  ( .A(\dp/alu_out_ex_o [26]), .ZN(\dp/n130 ) );
  OAI22_X1 \dp/U298  ( .A1(\dp/n851 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n130 ), .ZN(\dp/n915 ) );
  INV_X1 \dp/U297  ( .A(\dp/alu_out_ex_o [27]), .ZN(\dp/n129 ) );
  OAI22_X1 \dp/U296  ( .A1(\dp/n850 ), .A2(\dp/n33 ), .B1(\dp/n32 ), .B2(
        \dp/n129 ), .ZN(\dp/n914 ) );
  INV_X1 \dp/U295  ( .A(\dp/alu_out_ex_o [1]), .ZN(\dp/n157 ) );
  OAI22_X1 \dp/U294  ( .A1(\dp/n876 ), .A2(\dp/n35 ), .B1(\dp/n31 ), .B2(
        \dp/n157 ), .ZN(\dp/n940 ) );
  INV_X1 \dp/U293  ( .A(\dp/alu_out_ex_o [2]), .ZN(\dp/n156 ) );
  OAI22_X1 \dp/U292  ( .A1(\dp/n875 ), .A2(\dp/n35 ), .B1(\dp/n31 ), .B2(
        \dp/n156 ), .ZN(\dp/n939 ) );
  INV_X1 \dp/U291  ( .A(\dp/alu_out_ex_o [3]), .ZN(\dp/n155 ) );
  OAI22_X1 \dp/U290  ( .A1(\dp/n874 ), .A2(\dp/n35 ), .B1(\dp/n31 ), .B2(
        \dp/n155 ), .ZN(\dp/n938 ) );
  INV_X1 \dp/U289  ( .A(\dp/alu_out_ex_o [4]), .ZN(\dp/n154 ) );
  OAI22_X1 \dp/U288  ( .A1(\dp/n873 ), .A2(\dp/n35 ), .B1(\dp/n31 ), .B2(
        \dp/n154 ), .ZN(\dp/n937 ) );
  INV_X1 \dp/U287  ( .A(\dp/npc_if_o [9]), .ZN(\dp/n116 ) );
  OAI22_X1 \dp/U286  ( .A1(\dp/n83 ), .A2(\dp/n551 ), .B1(\dp/n74 ), .B2(
        \dp/n116 ), .ZN(\dp/n684 ) );
  INV_X1 \dp/U285  ( .A(\dp/npc_if_o [10]), .ZN(\dp/n115 ) );
  OAI22_X1 \dp/U284  ( .A1(\dp/n83 ), .A2(\dp/n552 ), .B1(\dp/n74 ), .B2(
        \dp/n115 ), .ZN(\dp/n685 ) );
  INV_X1 \dp/U283  ( .A(\dp/npc_if_o [11]), .ZN(\dp/n114 ) );
  OAI22_X1 \dp/U282  ( .A1(\dp/n83 ), .A2(\dp/n553 ), .B1(\dp/n74 ), .B2(
        \dp/n114 ), .ZN(\dp/n686 ) );
  INV_X1 \dp/U281  ( .A(\dp/npc_if_o [12]), .ZN(\dp/n113 ) );
  OAI22_X1 \dp/U280  ( .A1(\dp/n82 ), .A2(\dp/n554 ), .B1(\dp/n74 ), .B2(
        \dp/n113 ), .ZN(\dp/n687 ) );
  INV_X1 \dp/U279  ( .A(\dp/npc_if_o [13]), .ZN(\dp/n112 ) );
  OAI22_X1 \dp/U278  ( .A1(\dp/n82 ), .A2(\dp/n555 ), .B1(\dp/n74 ), .B2(
        \dp/n112 ), .ZN(\dp/n688 ) );
  INV_X1 \dp/U277  ( .A(\dp/npc_if_o [14]), .ZN(\dp/n111 ) );
  OAI22_X1 \dp/U276  ( .A1(\dp/n82 ), .A2(\dp/n556 ), .B1(\dp/n74 ), .B2(
        \dp/n111 ), .ZN(\dp/n689 ) );
  INV_X1 \dp/U275  ( .A(\dp/npc_if_o [15]), .ZN(\dp/n110 ) );
  OAI22_X1 \dp/U274  ( .A1(\dp/n82 ), .A2(\dp/n557 ), .B1(\dp/n74 ), .B2(
        \dp/n110 ), .ZN(\dp/n690 ) );
  INV_X1 \dp/U273  ( .A(\dp/npc_if_o [16]), .ZN(\dp/n109 ) );
  OAI22_X1 \dp/U272  ( .A1(\dp/n82 ), .A2(\dp/n558 ), .B1(\dp/n74 ), .B2(
        \dp/n109 ), .ZN(\dp/n691 ) );
  INV_X1 \dp/U271  ( .A(\dp/npc_if_o [17]), .ZN(\dp/n108 ) );
  OAI22_X1 \dp/U270  ( .A1(\dp/n82 ), .A2(\dp/n559 ), .B1(\dp/n74 ), .B2(
        \dp/n108 ), .ZN(\dp/n692 ) );
  INV_X1 \dp/U269  ( .A(\dp/npc_if_o [18]), .ZN(\dp/n107 ) );
  OAI22_X1 \dp/U268  ( .A1(\dp/n82 ), .A2(\dp/n560 ), .B1(\dp/n75 ), .B2(
        \dp/n107 ), .ZN(\dp/n693 ) );
  INV_X1 \dp/U267  ( .A(\dp/npc_if_o [19]), .ZN(\dp/n106 ) );
  OAI22_X1 \dp/U266  ( .A1(\dp/n82 ), .A2(\dp/n561 ), .B1(\dp/n75 ), .B2(
        \dp/n106 ), .ZN(\dp/n694 ) );
  AOI22_X1 \dp/U265  ( .A1(\dp/data_mem_ex_o [8]), .A2(\dp/n14 ), .B1(
        \dp/z_word [8]), .B2(\dp/n11 ), .ZN(\dp/n392 ) );
  OAI221_X1 \dp/U264  ( .B1(\dp/n238 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n358 ), .A(\dp/n392 ), .ZN(\dp/n996 ) );
  AOI22_X1 \dp/U263  ( .A1(\dp/data_mem_ex_o [9]), .A2(\dp/n14 ), .B1(
        \dp/z_word [9]), .B2(\dp/n11 ), .ZN(\dp/n391 ) );
  OAI221_X1 \dp/U262  ( .B1(\dp/n239 ), .B2(\dp/n18 ), .C1(\dp/n37 ), .C2(
        \dp/n357 ), .A(\dp/n391 ), .ZN(\dp/n995 ) );
  AOI22_X1 \dp/U261  ( .A1(\dp/data_mem_ex_o [10]), .A2(\dp/n14 ), .B1(
        \dp/z_word [10]), .B2(\dp/n11 ), .ZN(\dp/n390 ) );
  OAI221_X1 \dp/U260  ( .B1(\dp/n240 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n356 ), .A(\dp/n390 ), .ZN(\dp/n994 ) );
  AOI22_X1 \dp/U259  ( .A1(\dp/data_mem_ex_o [11]), .A2(\dp/n14 ), .B1(
        \dp/z_word [11]), .B2(\dp/n11 ), .ZN(\dp/n389 ) );
  OAI221_X1 \dp/U258  ( .B1(\dp/n241 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n355 ), .A(\dp/n389 ), .ZN(\dp/n993 ) );
  AOI22_X1 \dp/U257  ( .A1(\dp/data_mem_ex_o [12]), .A2(\dp/n14 ), .B1(
        \dp/z_word [12]), .B2(\dp/n11 ), .ZN(\dp/n388 ) );
  OAI221_X1 \dp/U256  ( .B1(\dp/n242 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n354 ), .A(\dp/n388 ), .ZN(\dp/n992 ) );
  AOI22_X1 \dp/U255  ( .A1(\dp/data_mem_ex_o [13]), .A2(\dp/n14 ), .B1(
        \dp/z_word [13]), .B2(\dp/n11 ), .ZN(\dp/n387 ) );
  OAI221_X1 \dp/U254  ( .B1(\dp/n243 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n353 ), .A(\dp/n387 ), .ZN(\dp/n991 ) );
  AOI22_X1 \dp/U253  ( .A1(\dp/data_mem_ex_o [14]), .A2(\dp/n14 ), .B1(
        \dp/z_word [14]), .B2(\dp/n11 ), .ZN(\dp/n386 ) );
  OAI221_X1 \dp/U252  ( .B1(\dp/n244 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n352 ), .A(\dp/n386 ), .ZN(\dp/n990 ) );
  AOI22_X1 \dp/U251  ( .A1(\dp/data_mem_ex_o [15]), .A2(\dp/n14 ), .B1(
        \dp/z_word [15]), .B2(\dp/n11 ), .ZN(\dp/n385 ) );
  OAI221_X1 \dp/U250  ( .B1(\dp/n245 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n351 ), .A(\dp/n385 ), .ZN(\dp/n989 ) );
  AOI22_X1 \dp/U249  ( .A1(\dp/data_mem_ex_o [16]), .A2(\dp/n14 ), .B1(
        \dp/z_word [16]), .B2(\dp/n11 ), .ZN(\dp/n384 ) );
  OAI221_X1 \dp/U248  ( .B1(\dp/n246 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n350 ), .A(\dp/n384 ), .ZN(\dp/n988 ) );
  AOI22_X1 \dp/U247  ( .A1(\dp/data_mem_ex_o [17]), .A2(\dp/n14 ), .B1(
        \dp/z_word [17]), .B2(\dp/n11 ), .ZN(\dp/n383 ) );
  OAI221_X1 \dp/U246  ( .B1(\dp/n247 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n349 ), .A(\dp/n383 ), .ZN(\dp/n987 ) );
  AOI22_X1 \dp/U245  ( .A1(\dp/data_mem_ex_o [18]), .A2(\dp/n14 ), .B1(
        \dp/z_word [18]), .B2(\dp/n11 ), .ZN(\dp/n382 ) );
  OAI221_X1 \dp/U244  ( .B1(\dp/n248 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n348 ), .A(\dp/n382 ), .ZN(\dp/n986 ) );
  AOI22_X1 \dp/U243  ( .A1(\dp/data_mem_ex_o [19]), .A2(\dp/n14 ), .B1(
        \dp/z_word [19]), .B2(\dp/n11 ), .ZN(\dp/n381 ) );
  OAI221_X1 \dp/U242  ( .B1(\dp/n249 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n347 ), .A(\dp/n381 ), .ZN(\dp/n985 ) );
  AOI22_X1 \dp/U241  ( .A1(\dp/data_mem_ex_o [20]), .A2(\dp/n13 ), .B1(
        \dp/z_word [20]), .B2(\dp/n10 ), .ZN(\dp/n380 ) );
  OAI221_X1 \dp/U240  ( .B1(\dp/n250 ), .B2(\dp/n17 ), .C1(\dp/n37 ), .C2(
        \dp/n346 ), .A(\dp/n380 ), .ZN(\dp/n984 ) );
  AOI22_X1 \dp/U239  ( .A1(\dp/data_mem_ex_o [21]), .A2(\dp/n13 ), .B1(
        \dp/z_word [21]), .B2(\dp/n10 ), .ZN(\dp/n379 ) );
  OAI221_X1 \dp/U238  ( .B1(\dp/n251 ), .B2(\dp/n16 ), .C1(\dp/n37 ), .C2(
        \dp/n345 ), .A(\dp/n379 ), .ZN(\dp/n983 ) );
  AOI22_X1 \dp/U237  ( .A1(\dp/data_mem_ex_o [22]), .A2(\dp/n13 ), .B1(
        \dp/z_word [22]), .B2(\dp/n10 ), .ZN(\dp/n378 ) );
  OAI221_X1 \dp/U236  ( .B1(\dp/n252 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n344 ), .A(\dp/n378 ), .ZN(\dp/n982 ) );
  AOI22_X1 \dp/U235  ( .A1(\dp/data_mem_ex_o [23]), .A2(\dp/n13 ), .B1(
        \dp/z_word [23]), .B2(\dp/n10 ), .ZN(\dp/n377 ) );
  OAI221_X1 \dp/U234  ( .B1(\dp/n253 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n343 ), .A(\dp/n377 ), .ZN(\dp/n981 ) );
  AOI22_X1 \dp/U233  ( .A1(\dp/data_mem_ex_o [24]), .A2(\dp/n13 ), .B1(
        \dp/z_word [24]), .B2(\dp/n10 ), .ZN(\dp/n376 ) );
  OAI221_X1 \dp/U232  ( .B1(\dp/n254 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n342 ), .A(\dp/n376 ), .ZN(\dp/n980 ) );
  AOI22_X1 \dp/U231  ( .A1(\dp/data_mem_ex_o [25]), .A2(\dp/n13 ), .B1(
        \dp/z_word [25]), .B2(\dp/n10 ), .ZN(\dp/n375 ) );
  OAI221_X1 \dp/U230  ( .B1(\dp/n255 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n341 ), .A(\dp/n375 ), .ZN(\dp/n979 ) );
  AOI22_X1 \dp/U229  ( .A1(\dp/data_mem_ex_o [26]), .A2(\dp/n13 ), .B1(
        \dp/z_word [26]), .B2(\dp/n10 ), .ZN(\dp/n374 ) );
  OAI221_X1 \dp/U228  ( .B1(\dp/n256 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n340 ), .A(\dp/n374 ), .ZN(\dp/n978 ) );
  AOI22_X1 \dp/U227  ( .A1(\dp/data_mem_ex_o [27]), .A2(\dp/n13 ), .B1(
        \dp/z_word [27]), .B2(\dp/n10 ), .ZN(\dp/n373 ) );
  OAI221_X1 \dp/U226  ( .B1(\dp/n257 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n339 ), .A(\dp/n373 ), .ZN(\dp/n977 ) );
  AOI22_X1 \dp/U225  ( .A1(\dp/data_mem_ex_o [28]), .A2(\dp/n13 ), .B1(
        \dp/z_word [28]), .B2(\dp/n10 ), .ZN(\dp/n372 ) );
  OAI221_X1 \dp/U224  ( .B1(\dp/n258 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n338 ), .A(\dp/n372 ), .ZN(\dp/n976 ) );
  AOI22_X1 \dp/U223  ( .A1(\dp/data_mem_ex_o [29]), .A2(\dp/n13 ), .B1(
        \dp/z_word [29]), .B2(\dp/n10 ), .ZN(\dp/n371 ) );
  OAI221_X1 \dp/U222  ( .B1(\dp/n259 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n337 ), .A(\dp/n371 ), .ZN(\dp/n975 ) );
  AOI22_X1 \dp/U221  ( .A1(\dp/data_mem_ex_o [30]), .A2(\dp/n13 ), .B1(
        \dp/z_word [30]), .B2(\dp/n10 ), .ZN(\dp/n370 ) );
  OAI221_X1 \dp/U220  ( .B1(\dp/n260 ), .B2(\dp/n16 ), .C1(\dp/n38 ), .C2(
        \dp/n336 ), .A(\dp/n370 ), .ZN(\dp/n974 ) );
  AOI22_X1 \dp/U219  ( .A1(\dp/data_mem_ex_o [31]), .A2(\dp/n13 ), .B1(
        \dp/z_word [31]), .B2(\dp/n10 ), .ZN(\dp/n367 ) );
  OAI221_X1 \dp/U218  ( .B1(\dp/n261 ), .B2(\dp/n16 ), .C1(\dp/n36 ), .C2(
        \dp/n335 ), .A(\dp/n367 ), .ZN(\dp/n973 ) );
  AOI22_X1 \dp/U217  ( .A1(\dp/data_mem_ex_o [0]), .A2(\dp/n15 ), .B1(
        \dp/z_word [0]), .B2(\dp/n12 ), .ZN(\dp/n401 ) );
  OAI221_X1 \dp/U216  ( .B1(\dp/n230 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n400 ), .A(\dp/n401 ), .ZN(\dp/n1004 ) );
  AOI22_X1 \dp/U215  ( .A1(\dp/data_mem_ex_o [1]), .A2(\dp/n15 ), .B1(
        \dp/z_word [1]), .B2(\dp/n12 ), .ZN(\dp/n399 ) );
  OAI221_X1 \dp/U214  ( .B1(\dp/n231 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n365 ), .A(\dp/n399 ), .ZN(\dp/n1003 ) );
  AOI22_X1 \dp/U213  ( .A1(\dp/data_mem_ex_o [2]), .A2(\dp/n15 ), .B1(
        \dp/z_word [2]), .B2(\dp/n12 ), .ZN(\dp/n398 ) );
  OAI221_X1 \dp/U212  ( .B1(\dp/n232 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n364 ), .A(\dp/n398 ), .ZN(\dp/n1002 ) );
  AOI22_X1 \dp/U211  ( .A1(\dp/data_mem_ex_o [3]), .A2(\dp/n15 ), .B1(
        \dp/z_word [3]), .B2(\dp/n12 ), .ZN(\dp/n397 ) );
  OAI221_X1 \dp/U210  ( .B1(\dp/n233 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n363 ), .A(\dp/n397 ), .ZN(\dp/n1001 ) );
  AOI22_X1 \dp/U209  ( .A1(\dp/data_mem_ex_o [4]), .A2(\dp/n15 ), .B1(
        \dp/z_word [4]), .B2(\dp/n12 ), .ZN(\dp/n396 ) );
  OAI221_X1 \dp/U208  ( .B1(\dp/n234 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n362 ), .A(\dp/n396 ), .ZN(\dp/n1000 ) );
  AOI22_X1 \dp/U207  ( .A1(\dp/data_mem_ex_o [5]), .A2(\dp/n15 ), .B1(
        \dp/z_word [5]), .B2(\dp/n12 ), .ZN(\dp/n395 ) );
  OAI221_X1 \dp/U206  ( .B1(\dp/n235 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n361 ), .A(\dp/n395 ), .ZN(\dp/n999 ) );
  AOI22_X1 \dp/U205  ( .A1(\dp/data_mem_ex_o [6]), .A2(\dp/n15 ), .B1(
        \dp/z_word [6]), .B2(\dp/n12 ), .ZN(\dp/n394 ) );
  OAI221_X1 \dp/U204  ( .B1(\dp/n236 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n360 ), .A(\dp/n394 ), .ZN(\dp/n998 ) );
  AOI22_X1 \dp/U203  ( .A1(\dp/data_mem_ex_o [7]), .A2(\dp/n15 ), .B1(
        \dp/z_word [7]), .B2(\dp/n12 ), .ZN(\dp/n393 ) );
  OAI221_X1 \dp/U202  ( .B1(\dp/n237 ), .B2(\dp/n18 ), .C1(\dp/n36 ), .C2(
        \dp/n359 ), .A(\dp/n393 ), .ZN(\dp/n997 ) );
  NOR3_X1 \dp/U201  ( .A1(mem_in_en_i), .A2(npc_wb_en_i), .A3(\dp/n31 ), .ZN(
        \dp/n368 ) );
  INV_X1 \dp/U200  ( .A(\dp/alu_out_ex_o [13]), .ZN(\dp/n145 ) );
  OAI22_X1 \dp/U199  ( .A1(\dp/n864 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n145 ), .ZN(\dp/n928 ) );
  INV_X1 \dp/U198  ( .A(\dp/alu_out_ex_o [14]), .ZN(\dp/n144 ) );
  OAI22_X1 \dp/U197  ( .A1(\dp/n863 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n144 ), .ZN(\dp/n927 ) );
  INV_X1 \dp/U196  ( .A(\dp/alu_out_ex_o [15]), .ZN(\dp/n143 ) );
  OAI22_X1 \dp/U195  ( .A1(\dp/n862 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n143 ), .ZN(\dp/n926 ) );
  INV_X1 \dp/U194  ( .A(\dp/alu_out_ex_o [16]), .ZN(\dp/n142 ) );
  OAI22_X1 \dp/U193  ( .A1(\dp/n861 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n142 ), .ZN(\dp/n925 ) );
  INV_X1 \dp/U192  ( .A(\dp/alu_out_ex_o [10]), .ZN(\dp/n148 ) );
  OAI22_X1 \dp/U191  ( .A1(\dp/n867 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n148 ), .ZN(\dp/n931 ) );
  INV_X1 \dp/U190  ( .A(\dp/alu_out_ex_o [11]), .ZN(\dp/n147 ) );
  OAI22_X1 \dp/U189  ( .A1(\dp/n866 ), .A2(\dp/n34 ), .B1(\dp/n32 ), .B2(
        \dp/n147 ), .ZN(\dp/n930 ) );
  INV_X1 \dp/U188  ( .A(\dp/alu_out_ex_o [0]), .ZN(\dp/n158 ) );
  OAI22_X1 \dp/U187  ( .A1(\dp/n877 ), .A2(\dp/n35 ), .B1(\dp/n31 ), .B2(
        \dp/n158 ), .ZN(\dp/n941 ) );
  INV_X1 \dp/U186  ( .A(\dp/npc_if_o [29]), .ZN(\dp/n96 ) );
  OAI22_X1 \dp/U185  ( .A1(\dp/n81 ), .A2(\dp/n571 ), .B1(\dp/n76 ), .B2(
        \dp/n96 ), .ZN(\dp/n704 ) );
  INV_X1 \dp/U184  ( .A(\dp/npc_if_o [30]), .ZN(\dp/n95 ) );
  OAI22_X1 \dp/U183  ( .A1(\dp/n81 ), .A2(\dp/n572 ), .B1(\dp/n76 ), .B2(
        \dp/n95 ), .ZN(\dp/n705 ) );
  INV_X1 \dp/U182  ( .A(\dp/npc_if_o [20]), .ZN(\dp/n105 ) );
  OAI22_X1 \dp/U181  ( .A1(\dp/n82 ), .A2(\dp/n562 ), .B1(\dp/n75 ), .B2(
        \dp/n105 ), .ZN(\dp/n695 ) );
  INV_X1 \dp/U180  ( .A(\dp/npc_if_o [21]), .ZN(\dp/n104 ) );
  OAI22_X1 \dp/U179  ( .A1(\dp/n82 ), .A2(\dp/n563 ), .B1(\dp/n75 ), .B2(
        \dp/n104 ), .ZN(\dp/n696 ) );
  INV_X1 \dp/U178  ( .A(\dp/npc_if_o [22]), .ZN(\dp/n103 ) );
  OAI22_X1 \dp/U177  ( .A1(\dp/n82 ), .A2(\dp/n564 ), .B1(\dp/n75 ), .B2(
        \dp/n103 ), .ZN(\dp/n697 ) );
  INV_X1 \dp/U176  ( .A(\dp/npc_if_o [23]), .ZN(\dp/n102 ) );
  OAI22_X1 \dp/U175  ( .A1(\dp/n82 ), .A2(\dp/n565 ), .B1(\dp/n75 ), .B2(
        \dp/n102 ), .ZN(\dp/n698 ) );
  INV_X1 \dp/U174  ( .A(\dp/npc_if_o [24]), .ZN(\dp/n101 ) );
  OAI22_X1 \dp/U173  ( .A1(\dp/n81 ), .A2(\dp/n566 ), .B1(\dp/n75 ), .B2(
        \dp/n101 ), .ZN(\dp/n699 ) );
  INV_X1 \dp/U172  ( .A(\dp/npc_if_o [25]), .ZN(\dp/n100 ) );
  OAI22_X1 \dp/U171  ( .A1(\dp/n81 ), .A2(\dp/n567 ), .B1(\dp/n75 ), .B2(
        \dp/n100 ), .ZN(\dp/n700 ) );
  INV_X1 \dp/U170  ( .A(\dp/npc_if_o [26]), .ZN(\dp/n99 ) );
  OAI22_X1 \dp/U169  ( .A1(\dp/n81 ), .A2(\dp/n568 ), .B1(\dp/n75 ), .B2(
        \dp/n99 ), .ZN(\dp/n701 ) );
  INV_X1 \dp/U168  ( .A(\dp/npc_if_o [27]), .ZN(\dp/n98 ) );
  OAI22_X1 \dp/U167  ( .A1(\dp/n81 ), .A2(\dp/n569 ), .B1(\dp/n75 ), .B2(
        \dp/n98 ), .ZN(\dp/n702 ) );
  INV_X1 \dp/U166  ( .A(\dp/npc_if_o [28]), .ZN(\dp/n97 ) );
  OAI22_X1 \dp/U165  ( .A1(\dp/n81 ), .A2(\dp/n570 ), .B1(\dp/n75 ), .B2(
        \dp/n97 ), .ZN(\dp/n703 ) );
  INV_X1 \dp/U164  ( .A(\dp/npc_if_o [31]), .ZN(\dp/n94 ) );
  OAI22_X1 \dp/U163  ( .A1(\dp/n81 ), .A2(\dp/n573 ), .B1(\dp/n76 ), .B2(
        \dp/n94 ), .ZN(\dp/n706 ) );
  NAND2_X1 \dp/U162  ( .A1(pipe_clear_n_i), .A2(\dp/n57 ), .ZN(\dp/n132 ) );
  OAI22_X1 \dp/U161  ( .A1(\dp/n224 ), .A2(\dp/n25 ), .B1(\dp/n24 ), .B2(
        \dp/n400 ), .ZN(\dp/n1015 ) );
  OAI22_X1 \dp/U160  ( .A1(\dp/n269 ), .A2(\dp/n25 ), .B1(\dp/n24 ), .B2(
        \dp/n365 ), .ZN(\dp/n972 ) );
  OAI22_X1 \dp/U159  ( .A1(\dp/n270 ), .A2(\dp/n25 ), .B1(\dp/n24 ), .B2(
        \dp/n364 ), .ZN(\dp/n971 ) );
  OAI22_X1 \dp/U158  ( .A1(\dp/n271 ), .A2(\dp/n25 ), .B1(\dp/n24 ), .B2(
        \dp/n363 ), .ZN(\dp/n970 ) );
  NAND2_X1 \dp/U157  ( .A1(pipe_clear_n_i), .A2(\dp/n79 ), .ZN(\dp/n69 ) );
  OAI22_X1 \dp/U156  ( .A1(\dp/n272 ), .A2(\dp/n25 ), .B1(\dp/n23 ), .B2(
        \dp/n362 ), .ZN(\dp/n969 ) );
  OAI22_X1 \dp/U155  ( .A1(\dp/n273 ), .A2(\dp/n25 ), .B1(\dp/n23 ), .B2(
        \dp/n361 ), .ZN(\dp/n968 ) );
  OAI22_X1 \dp/U154  ( .A1(\dp/n274 ), .A2(\dp/n25 ), .B1(\dp/n23 ), .B2(
        \dp/n360 ), .ZN(\dp/n967 ) );
  OAI22_X1 \dp/U153  ( .A1(\dp/n275 ), .A2(\dp/n25 ), .B1(\dp/n23 ), .B2(
        \dp/n359 ), .ZN(\dp/n966 ) );
  OAI22_X1 \dp/U152  ( .A1(\dp/n276 ), .A2(\dp/n25 ), .B1(\dp/n23 ), .B2(
        \dp/n358 ), .ZN(\dp/n965 ) );
  OAI22_X1 \dp/U151  ( .A1(\dp/n277 ), .A2(\dp/n25 ), .B1(\dp/n23 ), .B2(
        \dp/n357 ), .ZN(\dp/n964 ) );
  OAI22_X1 \dp/U150  ( .A1(\dp/n278 ), .A2(\dp/n27 ), .B1(\dp/n23 ), .B2(
        \dp/n356 ), .ZN(\dp/n963 ) );
  OAI22_X1 \dp/U149  ( .A1(\dp/n279 ), .A2(\dp/n26 ), .B1(\dp/n23 ), .B2(
        \dp/n355 ), .ZN(\dp/n962 ) );
  OAI22_X1 \dp/U148  ( .A1(\dp/n280 ), .A2(\dp/n26 ), .B1(\dp/n23 ), .B2(
        \dp/n354 ), .ZN(\dp/n961 ) );
  OAI22_X1 \dp/U147  ( .A1(\dp/n281 ), .A2(\dp/n26 ), .B1(\dp/n23 ), .B2(
        \dp/n353 ), .ZN(\dp/n960 ) );
  OAI22_X1 \dp/U146  ( .A1(\dp/n282 ), .A2(\dp/n26 ), .B1(\dp/n23 ), .B2(
        \dp/n352 ), .ZN(\dp/n959 ) );
  OAI22_X1 \dp/U145  ( .A1(\dp/n283 ), .A2(\dp/n26 ), .B1(\dp/n23 ), .B2(
        \dp/n351 ), .ZN(\dp/n958 ) );
  OAI22_X1 \dp/U144  ( .A1(\dp/n284 ), .A2(\dp/n26 ), .B1(\dp/n22 ), .B2(
        \dp/n350 ), .ZN(\dp/n957 ) );
  OAI22_X1 \dp/U143  ( .A1(\dp/n285 ), .A2(\dp/n26 ), .B1(\dp/n22 ), .B2(
        \dp/n349 ), .ZN(\dp/n956 ) );
  OAI22_X1 \dp/U142  ( .A1(\dp/n286 ), .A2(\dp/n26 ), .B1(\dp/n22 ), .B2(
        \dp/n348 ), .ZN(\dp/n955 ) );
  OAI22_X1 \dp/U141  ( .A1(\dp/n287 ), .A2(\dp/n26 ), .B1(\dp/n22 ), .B2(
        \dp/n347 ), .ZN(\dp/n954 ) );
  OAI22_X1 \dp/U140  ( .A1(\dp/n288 ), .A2(\dp/n26 ), .B1(\dp/n22 ), .B2(
        \dp/n346 ), .ZN(\dp/n953 ) );
  OAI22_X1 \dp/U139  ( .A1(\dp/n289 ), .A2(\dp/n26 ), .B1(\dp/n22 ), .B2(
        \dp/n345 ), .ZN(\dp/n952 ) );
  OAI22_X1 \dp/U138  ( .A1(\dp/n290 ), .A2(\dp/n26 ), .B1(\dp/n22 ), .B2(
        \dp/n344 ), .ZN(\dp/n951 ) );
  OAI22_X1 \dp/U137  ( .A1(\dp/n291 ), .A2(\dp/n27 ), .B1(\dp/n22 ), .B2(
        \dp/n343 ), .ZN(\dp/n950 ) );
  OAI22_X1 \dp/U136  ( .A1(\dp/n292 ), .A2(\dp/n27 ), .B1(\dp/n22 ), .B2(
        \dp/n342 ), .ZN(\dp/n949 ) );
  OAI22_X1 \dp/U135  ( .A1(\dp/n293 ), .A2(\dp/n27 ), .B1(\dp/n22 ), .B2(
        \dp/n341 ), .ZN(\dp/n948 ) );
  OAI22_X1 \dp/U134  ( .A1(\dp/n294 ), .A2(\dp/n27 ), .B1(\dp/n22 ), .B2(
        \dp/n340 ), .ZN(\dp/n947 ) );
  OAI22_X1 \dp/U133  ( .A1(\dp/n295 ), .A2(\dp/n27 ), .B1(\dp/n22 ), .B2(
        \dp/n339 ), .ZN(\dp/n946 ) );
  NAND2_X1 \dp/U132  ( .A1(pipe_clear_n_i), .A2(\dp/n25 ), .ZN(\dp/n302 ) );
  OAI22_X1 \dp/U131  ( .A1(\dp/n296 ), .A2(\dp/n27 ), .B1(\dp/n21 ), .B2(
        \dp/n338 ), .ZN(\dp/n945 ) );
  OAI22_X1 \dp/U130  ( .A1(\dp/n297 ), .A2(\dp/n27 ), .B1(\dp/n21 ), .B2(
        \dp/n337 ), .ZN(\dp/n944 ) );
  OAI22_X1 \dp/U129  ( .A1(\dp/n299 ), .A2(\dp/n27 ), .B1(\dp/n21 ), .B2(
        \dp/n336 ), .ZN(\dp/n943 ) );
  OAI22_X1 \dp/U128  ( .A1(\dp/n300 ), .A2(\dp/n27 ), .B1(\dp/n21 ), .B2(
        \dp/n335 ), .ZN(\dp/n942 ) );
  INV_X1 \dp/U127  ( .A(wb_mux_sel_i), .ZN(\dp/n93 ) );
  INV_X1 \dp/U126  ( .A(pipe_clear_n_i), .ZN(\dp/n263 ) );
  AND2_X1 \dp/U125  ( .A1(pipe_clear_n_i), .A2(\dp/n33 ), .ZN(\dp/n9 ) );
  NOR2_X1 \dp/U124  ( .A1(\dp/n632 ), .A2(\dp/n31 ), .ZN(\dp/n369 ) );
  BUF_X1 \dp/U123  ( .A(\dp/n366 ), .Z(\dp/n18 ) );
  BUF_X1 \dp/U122  ( .A(\dp/n366 ), .Z(\dp/n17 ) );
  BUF_X1 \dp/U121  ( .A(\dp/n366 ), .Z(\dp/n16 ) );
  BUF_X1 \dp/U120  ( .A(\dp/n368 ), .Z(\dp/n15 ) );
  BUF_X1 \dp/U119  ( .A(\dp/n368 ), .Z(\dp/n14 ) );
  BUF_X1 \dp/U118  ( .A(\dp/n368 ), .Z(\dp/n13 ) );
  OR2_X1 \dp/U117  ( .A1(pipe_if_id_en_i), .A2(\dp/n263 ), .ZN(\dp/n131 ) );
  OR2_X1 \dp/U116  ( .A1(pipe_if_id_en_i), .A2(\dp/n263 ), .ZN(\dp/n68 ) );
  OR2_X1 \dp/U115  ( .A1(pipe_if_id_en_i), .A2(\dp/n263 ), .ZN(\dp/n301 ) );
  BUF_X1 \dp/U114  ( .A(\dp/n302 ), .Z(\dp/n24 ) );
  BUF_X1 \dp/U113  ( .A(\dp/n69 ), .Z(\dp/n71 ) );
  BUF_X1 \dp/U112  ( .A(\dp/n69 ), .Z(\dp/n72 ) );
  BUF_X1 \dp/U111  ( .A(\dp/n69 ), .Z(\dp/n73 ) );
  BUF_X1 \dp/U110  ( .A(\dp/n69 ), .Z(\dp/n74 ) );
  BUF_X1 \dp/U109  ( .A(\dp/n69 ), .Z(\dp/n75 ) );
  BUF_X1 \dp/U108  ( .A(\dp/n302 ), .Z(\dp/n23 ) );
  BUF_X1 \dp/U107  ( .A(\dp/n302 ), .Z(\dp/n22 ) );
  BUF_X1 \dp/U106  ( .A(\dp/n302 ), .Z(\dp/n21 ) );
  BUF_X1 \dp/U105  ( .A(\dp/n302 ), .Z(\dp/n20 ) );
  BUF_X1 \dp/U104  ( .A(\dp/n302 ), .Z(\dp/n19 ) );
  INV_X1 \dp/U103  ( .A(\dp/n9 ), .ZN(\dp/n32 ) );
  BUF_X1 \dp/U102  ( .A(\dp/n93 ), .Z(\dp/n90 ) );
  BUF_X1 \dp/U101  ( .A(\dp/n93 ), .Z(\dp/n89 ) );
  BUF_X1 \dp/U100  ( .A(\dp/n93 ), .Z(\dp/n88 ) );
  BUF_X1 \dp/U99  ( .A(\dp/n93 ), .Z(\dp/n87 ) );
  BUF_X1 \dp/U98  ( .A(\dp/n93 ), .Z(\dp/n86 ) );
  BUF_X1 \dp/U97  ( .A(\dp/n93 ), .Z(\dp/n91 ) );
  BUF_X1 \dp/U96  ( .A(\dp/n93 ), .Z(\dp/n92 ) );
  OR2_X1 \dp/U95  ( .A1(pipe_if_id_en_i), .A2(\dp/n263 ), .ZN(\dp/n298 ) );
  BUF_X1 \dp/U94  ( .A(\dp/n369 ), .Z(\dp/n12 ) );
  BUF_X1 \dp/U93  ( .A(\dp/n369 ), .Z(\dp/n11 ) );
  BUF_X1 \dp/U92  ( .A(\dp/n369 ), .Z(\dp/n10 ) );
  INV_X1 \dp/U91  ( .A(\dp/n9 ), .ZN(\dp/n31 ) );
  BUF_X1 \dp/U90  ( .A(\dp/n68 ), .Z(\dp/n78 ) );
  BUF_X1 \dp/U89  ( .A(\dp/n68 ), .Z(\dp/n77 ) );
  BUF_X1 \dp/U88  ( .A(\dp/n131 ), .Z(\dp/n56 ) );
  BUF_X1 \dp/U87  ( .A(\dp/n131 ), .Z(\dp/n55 ) );
  BUF_X1 \dp/U86  ( .A(\dp/n39 ), .Z(\dp/n43 ) );
  BUF_X1 \dp/U85  ( .A(\dp/n39 ), .Z(\dp/n44 ) );
  BUF_X1 \dp/U84  ( .A(\dp/n39 ), .Z(\dp/n45 ) );
  BUF_X1 \dp/U83  ( .A(\dp/n40 ), .Z(\dp/n46 ) );
  BUF_X1 \dp/U82  ( .A(\dp/n40 ), .Z(\dp/n47 ) );
  BUF_X1 \dp/U81  ( .A(\dp/n40 ), .Z(\dp/n48 ) );
  BUF_X1 \dp/U80  ( .A(\dp/n41 ), .Z(\dp/n49 ) );
  BUF_X1 \dp/U79  ( .A(\dp/n41 ), .Z(\dp/n50 ) );
  BUF_X1 \dp/U78  ( .A(\dp/n41 ), .Z(\dp/n51 ) );
  BUF_X1 \dp/U77  ( .A(\dp/n42 ), .Z(\dp/n52 ) );
  BUF_X1 \dp/U76  ( .A(\dp/n42 ), .Z(\dp/n53 ) );
  BUF_X1 \dp/U75  ( .A(\dp/n42 ), .Z(\dp/n54 ) );
  BUF_X1 \dp/U74  ( .A(\dp/n298 ), .Z(\dp/n38 ) );
  BUF_X1 \dp/U73  ( .A(\dp/n301 ), .Z(\dp/n30 ) );
  BUF_X1 \dp/U72  ( .A(\dp/n298 ), .Z(\dp/n37 ) );
  BUF_X1 \dp/U71  ( .A(\dp/n298 ), .Z(\dp/n35 ) );
  BUF_X1 \dp/U70  ( .A(\dp/n298 ), .Z(\dp/n36 ) );
  BUF_X1 \dp/U69  ( .A(\dp/n301 ), .Z(\dp/n27 ) );
  BUF_X1 \dp/U68  ( .A(\dp/n301 ), .Z(\dp/n26 ) );
  BUF_X1 \dp/U67  ( .A(\dp/n301 ), .Z(\dp/n28 ) );
  BUF_X1 \dp/U66  ( .A(\dp/n298 ), .Z(\dp/n34 ) );
  BUF_X1 \dp/U65  ( .A(\dp/n301 ), .Z(\dp/n29 ) );
  BUF_X1 \dp/U64  ( .A(\dp/n301 ), .Z(\dp/n25 ) );
  BUF_X1 \dp/U63  ( .A(\dp/n298 ), .Z(\dp/n33 ) );
  BUF_X1 \dp/U62  ( .A(\dp/n78 ), .Z(\dp/n83 ) );
  BUF_X1 \dp/U61  ( .A(\dp/n78 ), .Z(\dp/n82 ) );
  BUF_X1 \dp/U60  ( .A(\dp/n56 ), .Z(\dp/n67 ) );
  BUF_X1 \dp/U59  ( .A(\dp/n56 ), .Z(\dp/n66 ) );
  BUF_X1 \dp/U58  ( .A(\dp/n56 ), .Z(\dp/n65 ) );
  BUF_X1 \dp/U57  ( .A(\dp/n56 ), .Z(\dp/n64 ) );
  BUF_X1 \dp/U56  ( .A(\dp/n56 ), .Z(\dp/n63 ) );
  BUF_X1 \dp/U55  ( .A(\dp/n55 ), .Z(\dp/n62 ) );
  BUF_X1 \dp/U54  ( .A(\dp/n55 ), .Z(\dp/n61 ) );
  BUF_X1 \dp/U53  ( .A(\dp/n55 ), .Z(\dp/n60 ) );
  BUF_X1 \dp/U52  ( .A(\dp/n77 ), .Z(\dp/n81 ) );
  BUF_X1 \dp/U51  ( .A(\dp/n55 ), .Z(\dp/n59 ) );
  BUF_X1 \dp/U50  ( .A(\dp/n77 ), .Z(\dp/n80 ) );
  BUF_X1 \dp/U49  ( .A(\dp/n55 ), .Z(\dp/n58 ) );
  BUF_X1 \dp/U48  ( .A(\dp/n77 ), .Z(\dp/n79 ) );
  BUF_X1 \dp/U47  ( .A(\dp/n55 ), .Z(\dp/n57 ) );
  OAI22_X4 \dp/U46  ( .A1(\dp/n86 ), .A2(\dp/n303 ), .B1(\dp/n85 ), .B2(
        \dp/n224 ), .ZN(\dp/wr_data_id_i [0]) );
  OAI22_X4 \dp/U45  ( .A1(\dp/n88 ), .A2(\dp/n304 ), .B1(\dp/n85 ), .B2(
        \dp/n269 ), .ZN(\dp/wr_data_id_i [1]) );
  OAI22_X4 \dp/U44  ( .A1(\dp/n90 ), .A2(\dp/n305 ), .B1(\dp/n84 ), .B2(
        \dp/n270 ), .ZN(\dp/wr_data_id_i [2]) );
  OAI22_X4 \dp/U43  ( .A1(\dp/n91 ), .A2(\dp/n306 ), .B1(\dp/n84 ), .B2(
        \dp/n271 ), .ZN(\dp/wr_data_id_i [3]) );
  OAI22_X4 \dp/U42  ( .A1(\dp/n86 ), .A2(\dp/n313 ), .B1(\dp/n84 ), .B2(
        \dp/n278 ), .ZN(\dp/wr_data_id_i [10]) );
  OAI22_X4 \dp/U41  ( .A1(\dp/n88 ), .A2(\dp/n322 ), .B1(\dp/n85 ), .B2(
        \dp/n287 ), .ZN(\dp/wr_data_id_i [19]) );
  OAI22_X4 \dp/U40  ( .A1(\dp/n91 ), .A2(\dp/n307 ), .B1(\dp/n84 ), .B2(
        \dp/n272 ), .ZN(\dp/wr_data_id_i [4]) );
  OAI22_X4 \dp/U39  ( .A1(\dp/n86 ), .A2(\dp/n314 ), .B1(\dp/n85 ), .B2(
        \dp/n279 ), .ZN(\dp/wr_data_id_i [11]) );
  OAI22_X4 \dp/U38  ( .A1(\dp/n88 ), .A2(\dp/n323 ), .B1(\dp/n85 ), .B2(
        \dp/n288 ), .ZN(\dp/wr_data_id_i [20]) );
  OAI22_X4 \dp/U37  ( .A1(\dp/n91 ), .A2(\dp/n308 ), .B1(\dp/n84 ), .B2(
        \dp/n273 ), .ZN(\dp/wr_data_id_i [5]) );
  OAI22_X4 \dp/U36  ( .A1(\dp/n86 ), .A2(\dp/n315 ), .B1(\dp/n84 ), .B2(
        \dp/n280 ), .ZN(\dp/wr_data_id_i [12]) );
  OAI22_X4 \dp/U35  ( .A1(\dp/n88 ), .A2(\dp/n324 ), .B1(\dp/n85 ), .B2(
        \dp/n289 ), .ZN(\dp/wr_data_id_i [21]) );
  OAI22_X4 \dp/U34  ( .A1(\dp/n91 ), .A2(\dp/n309 ), .B1(\dp/n84 ), .B2(
        \dp/n274 ), .ZN(\dp/wr_data_id_i [6]) );
  OAI22_X4 \dp/U33  ( .A1(\dp/n86 ), .A2(\dp/n316 ), .B1(\dp/n85 ), .B2(
        \dp/n281 ), .ZN(\dp/wr_data_id_i [13]) );
  OAI22_X4 \dp/U32  ( .A1(\dp/n88 ), .A2(\dp/n325 ), .B1(\dp/n85 ), .B2(
        \dp/n290 ), .ZN(\dp/wr_data_id_i [22]) );
  INV_X2 \dp/U31  ( .A(\dp/n92 ), .ZN(\dp/n84 ) );
  OAI22_X4 \dp/U30  ( .A1(\dp/n91 ), .A2(\dp/n310 ), .B1(\dp/n84 ), .B2(
        \dp/n275 ), .ZN(\dp/wr_data_id_i [7]) );
  OAI22_X4 \dp/U29  ( .A1(\dp/n92 ), .A2(\dp/n311 ), .B1(\dp/n84 ), .B2(
        \dp/n276 ), .ZN(\dp/wr_data_id_i [8]) );
  OAI22_X4 \dp/U28  ( .A1(\dp/n87 ), .A2(\dp/n317 ), .B1(\dp/n84 ), .B2(
        \dp/n282 ), .ZN(\dp/wr_data_id_i [14]) );
  INV_X2 \dp/U27  ( .A(\dp/n92 ), .ZN(\dp/n85 ) );
  OAI22_X4 \dp/U26  ( .A1(\dp/n89 ), .A2(\dp/n326 ), .B1(\dp/n85 ), .B2(
        \dp/n291 ), .ZN(\dp/wr_data_id_i [23]) );
  OAI22_X4 \dp/U25  ( .A1(\dp/n90 ), .A2(\dp/n331 ), .B1(\dp/n85 ), .B2(
        \dp/n296 ), .ZN(\dp/wr_data_id_i [28]) );
  OAI22_X4 \dp/U24  ( .A1(\dp/n92 ), .A2(\dp/n312 ), .B1(\dp/n84 ), .B2(
        \dp/n277 ), .ZN(\dp/wr_data_id_i [9]) );
  OAI22_X4 \dp/U23  ( .A1(\dp/n87 ), .A2(\dp/n318 ), .B1(\dp/n84 ), .B2(
        \dp/n283 ), .ZN(\dp/wr_data_id_i [15]) );
  OAI22_X4 \dp/U22  ( .A1(\dp/n89 ), .A2(\dp/n327 ), .B1(\dp/n85 ), .B2(
        \dp/n292 ), .ZN(\dp/wr_data_id_i [24]) );
  OAI22_X4 \dp/U21  ( .A1(\dp/n87 ), .A2(\dp/n319 ), .B1(\dp/n85 ), .B2(
        \dp/n284 ), .ZN(\dp/wr_data_id_i [16]) );
  OAI22_X4 \dp/U20  ( .A1(\dp/n89 ), .A2(\dp/n328 ), .B1(\dp/n85 ), .B2(
        \dp/n293 ), .ZN(\dp/wr_data_id_i [25]) );
  OAI22_X4 \dp/U19  ( .A1(\dp/n90 ), .A2(\dp/n332 ), .B1(\dp/n84 ), .B2(
        \dp/n297 ), .ZN(\dp/wr_data_id_i [29]) );
  OAI22_X4 \dp/U18  ( .A1(\dp/n87 ), .A2(\dp/n320 ), .B1(\dp/n84 ), .B2(
        \dp/n285 ), .ZN(\dp/wr_data_id_i [17]) );
  OAI22_X4 \dp/U17  ( .A1(\dp/n89 ), .A2(\dp/n329 ), .B1(\dp/n85 ), .B2(
        \dp/n294 ), .ZN(\dp/wr_data_id_i [26]) );
  OAI22_X4 \dp/U16  ( .A1(\dp/n90 ), .A2(\dp/n333 ), .B1(\dp/n84 ), .B2(
        \dp/n299 ), .ZN(\dp/wr_data_id_i [30]) );
  INV_X16 \dp/U15  ( .A(RST), .ZN(\dp/n634 ) );
  OAI22_X1 \dp/U14  ( .A1(\dp/n90 ), .A2(\dp/n630 ), .B1(\dp/n84 ), .B2(
        \dp/n300 ), .ZN(\dp/wr_data_id_i [31]) );
  INV_X1 \dp/U13  ( .A(\dp/n7 ), .ZN(\dp/n8 ) );
  INV_X1 \dp/U12  ( .A(\dp/wr_data_id_i [31]), .ZN(\dp/n7 ) );
  OAI22_X1 \dp/U11  ( .A1(\dp/n89 ), .A2(\dp/n330 ), .B1(\dp/n85 ), .B2(
        \dp/n295 ), .ZN(\dp/wr_data_id_i [27]) );
  INV_X1 \dp/U10  ( .A(\dp/n5 ), .ZN(\dp/n6 ) );
  INV_X1 \dp/U9  ( .A(\dp/wr_data_id_i [27]), .ZN(\dp/n5 ) );
  OAI22_X1 \dp/U8  ( .A1(\dp/n87 ), .A2(\dp/n321 ), .B1(\dp/n85 ), .B2(
        \dp/n286 ), .ZN(\dp/wr_data_id_i [18]) );
  INV_X1 \dp/U7  ( .A(\dp/n3 ), .ZN(\dp/n4 ) );
  INV_X1 \dp/U6  ( .A(\dp/wr_data_id_i [18]), .ZN(\dp/n3 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[0]  ( .D(\dp/n941 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[0]), .QN(\dp/n877 ) );
  DFFR_X1 \dp/npc_id_i_reg[31]  ( .D(\dp/n706 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [31]), .QN(\dp/n573 ) );
  DFFR_X1 \dp/npc_id_i_reg[30]  ( .D(\dp/n705 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [30]), .QN(\dp/n572 ) );
  DFFR_X1 \dp/npc_id_i_reg[29]  ( .D(\dp/n704 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [29]), .QN(\dp/n571 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[4]  ( .D(\dp/n937 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[4]), .QN(\dp/n873 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[6]  ( .D(\dp/n935 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[6]), .QN(\dp/n871 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[5]  ( .D(\dp/n936 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[5]), .QN(\dp/n872 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[1]  ( .D(\dp/n940 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[1]), .QN(\dp/n876 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[2]  ( .D(\dp/n939 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[2]), .QN(\dp/n875 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[17]  ( .D(\dp/n924 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[17]), .QN(\dp/n860 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[16]  ( .D(\dp/n925 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[16]), .QN(\dp/n861 ) );
  DFFR_X1 \dp/npc_id_i_reg[28]  ( .D(\dp/n703 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [28]), .QN(\dp/n570 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[3]  ( .D(\dp/n938 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[3]), .QN(\dp/n874 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[18]  ( .D(\dp/n923 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[18]), .QN(\dp/n859 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[8]  ( .D(\dp/n933 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[8]), .QN(\dp/n869 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[9]  ( .D(\dp/n932 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[9]), .QN(\dp/n868 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[10]  ( .D(\dp/n931 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[10]), .QN(\dp/n867 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[20]  ( .D(\dp/n921 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[20]), .QN(\dp/n857 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[19]  ( .D(\dp/n922 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[19]), .QN(\dp/n858 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[21]  ( .D(\dp/n920 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[21]), .QN(\dp/n856 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[22]  ( .D(\dp/n919 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[22]), .QN(\dp/n855 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[23]  ( .D(\dp/n918 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[23]), .QN(\dp/n854 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[24]  ( .D(\dp/n917 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[24]), .QN(\dp/n853 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[25]  ( .D(\dp/n916 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[25]), .QN(\dp/n852 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[26]  ( .D(\dp/n915 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[26]), .QN(\dp/n851 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[27]  ( .D(\dp/n914 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[27]), .QN(\dp/n850 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[28]  ( .D(\dp/n913 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[28]), .QN(\dp/n849 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[29]  ( .D(\dp/n912 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[29]), .QN(\dp/n848 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[30]  ( .D(\dp/n911 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[30]), .QN(\dp/n847 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[31]  ( .D(\dp/n910 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[31]), .QN(\dp/n846 ) );
  DFFR_X1 \dp/npc_id_i_reg[27]  ( .D(\dp/n702 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [27]), .QN(\dp/n569 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[11]  ( .D(\dp/n930 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[11]), .QN(\dp/n866 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[14]  ( .D(\dp/n927 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[14]), .QN(\dp/n863 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[12]  ( .D(\dp/n929 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[12]), .QN(\dp/n865 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[13]  ( .D(\dp/n928 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[13]), .QN(\dp/n864 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[7]  ( .D(\dp/n934 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[7]), .QN(\dp/n870 ) );
  DFFR_X1 \dp/alu_out_mem_i_reg[15]  ( .D(\dp/n926 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_ADDRESS[15]), .QN(\dp/n862 ) );
  DFFR_X1 \dp/npc_id_i_reg[26]  ( .D(\dp/n701 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [26]), .QN(\dp/n568 ) );
  DFFR_X1 \dp/npc_id_i_reg[25]  ( .D(\dp/n700 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [25]), .QN(\dp/n567 ) );
  DFFR_X1 \dp/npc_id_i_reg[24]  ( .D(\dp/n699 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [24]), .QN(\dp/n566 ) );
  DFFR_X1 \dp/npc_id_i_reg[23]  ( .D(\dp/n698 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [23]), .QN(\dp/n565 ) );
  DFFR_X1 \dp/npc_id_i_reg[22]  ( .D(\dp/n697 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [22]), .QN(\dp/n564 ) );
  DFFR_X1 \dp/npc_id_i_reg[21]  ( .D(\dp/n696 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [21]), .QN(\dp/n563 ) );
  DFFR_X1 \dp/npc_id_i_reg[20]  ( .D(\dp/n695 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [20]), .QN(\dp/n562 ) );
  DFFR_X1 \dp/npc_id_i_reg[19]  ( .D(\dp/n694 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [19]), .QN(\dp/n561 ) );
  DFFR_X1 \dp/npc_id_i_reg[18]  ( .D(\dp/n693 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [18]), .QN(\dp/n560 ) );
  DFFR_X1 \dp/npc_id_i_reg[17]  ( .D(\dp/n692 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [17]), .QN(\dp/n559 ) );
  DFFR_X1 \dp/npc_id_i_reg[16]  ( .D(\dp/n691 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [16]), .QN(\dp/n558 ) );
  DFFR_X1 \dp/npc_id_i_reg[15]  ( .D(\dp/n690 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [15]), .QN(\dp/n557 ) );
  DFFR_X1 \dp/npc_id_i_reg[14]  ( .D(\dp/n689 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [14]), .QN(\dp/n556 ) );
  DFFR_X1 \dp/npc_id_i_reg[13]  ( .D(\dp/n688 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [13]), .QN(\dp/n555 ) );
  DFFR_X1 \dp/imm_ex_i_reg[0]  ( .D(\dp/n749 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [0]), .QN(\dp/n419 ) );
  DFFR_X1 \dp/imm_ex_i_reg[1]  ( .D(\dp/n750 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [1]), .QN(\dp/n420 ) );
  DFFR_X1 \dp/imm_ex_i_reg[2]  ( .D(\dp/n751 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [2]), .QN(\dp/n421 ) );
  DFFR_X1 \dp/imm_ex_i_reg[3]  ( .D(\dp/n752 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [3]), .QN(\dp/n422 ) );
  DFFR_X1 \dp/imm_ex_i_reg[4]  ( .D(\dp/n753 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [4]), .QN(\dp/n423 ) );
  DFFR_X1 \dp/imm_ex_i_reg[5]  ( .D(\dp/n754 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [5]), .QN(\dp/n424 ) );
  DFFR_X1 \dp/imm_ex_i_reg[6]  ( .D(\dp/n755 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [6]), .QN(\dp/n425 ) );
  DFFR_X1 \dp/imm_ex_i_reg[7]  ( .D(\dp/n756 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [7]), .QN(\dp/n426 ) );
  DFFR_X1 \dp/imm_ex_i_reg[8]  ( .D(\dp/n757 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [8]), .QN(\dp/n427 ) );
  DFFR_X1 \dp/imm_ex_i_reg[9]  ( .D(\dp/n758 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [9]), .QN(\dp/n428 ) );
  DFFR_X1 \dp/imm_ex_i_reg[10]  ( .D(\dp/n759 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [10]), .QN(\dp/n429 ) );
  DFFR_X1 \dp/imm_ex_i_reg[11]  ( .D(\dp/n760 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [11]), .QN(\dp/n430 ) );
  DFFR_X1 \dp/imm_ex_i_reg[12]  ( .D(\dp/n761 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [12]), .QN(\dp/n431 ) );
  DFFR_X1 \dp/imm_ex_i_reg[13]  ( .D(\dp/n762 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [13]), .QN(\dp/n432 ) );
  DFFR_X1 \dp/imm_ex_i_reg[14]  ( .D(\dp/n763 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [14]), .QN(\dp/n433 ) );
  DFFR_X1 \dp/imm_ex_i_reg[15]  ( .D(\dp/n764 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [15]), .QN(\dp/n434 ) );
  DFFR_X1 \dp/imm_ex_i_reg[16]  ( .D(\dp/n765 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [16]), .QN(\dp/n435 ) );
  DFFR_X1 \dp/imm_ex_i_reg[17]  ( .D(\dp/n766 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [17]), .QN(\dp/n436 ) );
  DFFR_X1 \dp/imm_ex_i_reg[18]  ( .D(\dp/n767 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [18]), .QN(\dp/n437 ) );
  DFFR_X1 \dp/imm_ex_i_reg[19]  ( .D(\dp/n768 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [19]), .QN(\dp/n438 ) );
  DFFR_X1 \dp/imm_ex_i_reg[20]  ( .D(\dp/n769 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [20]), .QN(\dp/n439 ) );
  DFFR_X1 \dp/imm_ex_i_reg[21]  ( .D(\dp/n770 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [21]), .QN(\dp/n440 ) );
  DFFR_X1 \dp/imm_ex_i_reg[22]  ( .D(\dp/n771 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [22]), .QN(\dp/n441 ) );
  DFFR_X1 \dp/imm_ex_i_reg[23]  ( .D(\dp/n772 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [23]), .QN(\dp/n442 ) );
  DFFR_X1 \dp/imm_ex_i_reg[24]  ( .D(\dp/n773 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [24]), .QN(\dp/n443 ) );
  DFFR_X1 \dp/imm_ex_i_reg[25]  ( .D(\dp/n774 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [25]), .QN(\dp/n444 ) );
  DFFR_X1 \dp/imm_ex_i_reg[26]  ( .D(\dp/n775 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [26]), .QN(\dp/n445 ) );
  DFFR_X1 \dp/imm_ex_i_reg[27]  ( .D(\dp/n776 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [27]), .QN(\dp/n446 ) );
  DFFR_X1 \dp/imm_ex_i_reg[28]  ( .D(\dp/n777 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [28]), .QN(\dp/n447 ) );
  DFFR_X1 \dp/imm_ex_i_reg[29]  ( .D(\dp/n778 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [29]), .QN(\dp/n448 ) );
  DFFR_X1 \dp/imm_ex_i_reg[30]  ( .D(\dp/n779 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [30]), .QN(\dp/n449 ) );
  DFFR_X1 \dp/imm_ex_i_reg[31]  ( .D(\dp/n780 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/imm_ex_i [31]), .QN(\dp/n450 ) );
  DFFR_X1 \dp/rd_fwd_ex_i_reg[0]  ( .D(\dp/n712 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_ex_o [0]), .QN(\dp/n414 ) );
  DFFR_X1 \dp/rd_fwd_ex_i_reg[1]  ( .D(\dp/n713 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_ex_o [1]), .QN(\dp/n415 ) );
  DFFR_X1 \dp/rd_fwd_ex_i_reg[2]  ( .D(\dp/n714 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_ex_o [2]), .QN(\dp/n416 ) );
  DFFR_X1 \dp/rd_fwd_ex_i_reg[3]  ( .D(\dp/n715 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_ex_o [3]), .QN(\dp/n417 ) );
  DFFR_X1 \dp/rd_fwd_ex_i_reg[4]  ( .D(\dp/n716 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_ex_o [4]), .QN(\dp/n418 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[0]  ( .D(\dp/n813 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [0]), .QN(\dp/n483 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[1]  ( .D(\dp/n814 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [1]), .QN(\dp/n484 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[2]  ( .D(\dp/n815 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [2]), .QN(\dp/n485 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[3]  ( .D(\dp/n816 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [3]), .QN(\dp/n486 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[4]  ( .D(\dp/n817 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [4]), .QN(\dp/n487 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[5]  ( .D(\dp/n818 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [5]), .QN(\dp/n488 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[6]  ( .D(\dp/n819 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [6]), .QN(\dp/n489 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[7]  ( .D(\dp/n820 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [7]), .QN(\dp/n490 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[8]  ( .D(\dp/n821 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [8]), .QN(\dp/n491 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[9]  ( .D(\dp/n822 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [9]), .QN(\dp/n492 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[10]  ( .D(\dp/n823 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [10]), .QN(\dp/n493 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[11]  ( .D(\dp/n824 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [11]), .QN(\dp/n494 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[12]  ( .D(\dp/n825 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [12]), .QN(\dp/n495 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[13]  ( .D(\dp/n826 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [13]), .QN(\dp/n496 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[14]  ( .D(\dp/n827 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [14]), .QN(\dp/n497 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[15]  ( .D(\dp/n828 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [15]), .QN(\dp/n498 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[16]  ( .D(\dp/n829 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [16]), .QN(\dp/n499 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[17]  ( .D(\dp/n830 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [17]), .QN(\dp/n500 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[18]  ( .D(\dp/n831 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [18]), .QN(\dp/n501 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[19]  ( .D(\dp/n832 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [19]), .QN(\dp/n502 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[20]  ( .D(\dp/n833 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [20]), .QN(\dp/n503 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[21]  ( .D(\dp/n834 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [21]), .QN(\dp/n504 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[22]  ( .D(\dp/n835 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [22]), .QN(\dp/n505 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[23]  ( .D(\dp/n836 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [23]), .QN(\dp/n506 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[24]  ( .D(\dp/n837 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [24]), .QN(\dp/n507 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[25]  ( .D(\dp/n838 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [25]), .QN(\dp/n508 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[26]  ( .D(\dp/n839 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [26]), .QN(\dp/n509 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[27]  ( .D(\dp/n840 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [27]), .QN(\dp/n510 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[28]  ( .D(\dp/n841 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [28]), .QN(\dp/n511 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[29]  ( .D(\dp/n842 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [29]), .QN(\dp/n512 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[30]  ( .D(\dp/n843 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [30]), .QN(\dp/n513 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[0]  ( .D(\dp/n781 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [0]), .QN(\dp/n451 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[1]  ( .D(\dp/n782 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [1]), .QN(\dp/n452 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[2]  ( .D(\dp/n783 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [2]), .QN(\dp/n453 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[3]  ( .D(\dp/n784 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [3]), .QN(\dp/n454 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[4]  ( .D(\dp/n785 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [4]), .QN(\dp/n455 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[5]  ( .D(\dp/n786 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [5]), .QN(\dp/n456 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[6]  ( .D(\dp/n787 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [6]), .QN(\dp/n457 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[7]  ( .D(\dp/n788 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [7]), .QN(\dp/n458 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[8]  ( .D(\dp/n789 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [8]), .QN(\dp/n459 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[9]  ( .D(\dp/n790 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [9]), .QN(\dp/n460 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[10]  ( .D(\dp/n791 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [10]), .QN(\dp/n461 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[11]  ( .D(\dp/n792 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [11]), .QN(\dp/n462 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[12]  ( .D(\dp/n793 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [12]), .QN(\dp/n463 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[13]  ( .D(\dp/n794 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [13]), .QN(\dp/n464 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[14]  ( .D(\dp/n795 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [14]), .QN(\dp/n465 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[15]  ( .D(\dp/n796 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [15]), .QN(\dp/n466 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[16]  ( .D(\dp/n797 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [16]), .QN(\dp/n467 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[17]  ( .D(\dp/n798 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [17]), .QN(\dp/n468 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[18]  ( .D(\dp/n799 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [18]), .QN(\dp/n469 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[19]  ( .D(\dp/n800 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [19]), .QN(\dp/n470 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[20]  ( .D(\dp/n801 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [20]), .QN(\dp/n471 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[21]  ( .D(\dp/n802 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [21]), .QN(\dp/n472 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[22]  ( .D(\dp/n803 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [22]), .QN(\dp/n473 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[23]  ( .D(\dp/n804 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [23]), .QN(\dp/n474 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[24]  ( .D(\dp/n805 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [24]), .QN(\dp/n475 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[25]  ( .D(\dp/n806 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [25]), .QN(\dp/n476 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[26]  ( .D(\dp/n807 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [26]), .QN(\dp/n477 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[27]  ( .D(\dp/n808 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [27]), .QN(\dp/n478 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[28]  ( .D(\dp/n809 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [28]), .QN(\dp/n479 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[29]  ( .D(\dp/n810 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [29]), .QN(\dp/n480 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[30]  ( .D(\dp/n811 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [30]), .QN(\dp/n481 ) );
  DFFR_X1 \dp/rf_out2_ex_i_reg[31]  ( .D(\dp/n812 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/data_mem_ex_o [31]), .QN(\dp/n482 ) );
  DFFR_X1 \dp/npc_id_i_reg[12]  ( .D(\dp/n687 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [12]), .QN(\dp/n554 ) );
  DFFR_X1 \dp/ir_reg[0]  ( .D(\dp/n649 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[0] ), .QN(\dp/n526 ) );
  DFFR_X1 \dp/ir_reg[1]  ( .D(\dp/n650 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[1] ), .QN(\dp/n527 ) );
  DFFR_X1 \dp/ir_reg[2]  ( .D(\dp/n651 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[2] ), .QN(\dp/n528 ) );
  DFFR_X1 \dp/ir_reg[3]  ( .D(\dp/n652 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[3] ), .QN(\dp/n529 ) );
  DFFR_X1 \dp/ir_reg[4]  ( .D(\dp/n653 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[4] ), .QN(\dp/n530 ) );
  DFFR_X1 \dp/ir_reg[5]  ( .D(\dp/n654 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[5] ), .QN(\dp/n531 ) );
  DFFR_X1 \dp/ir_reg[6]  ( .D(\dp/n655 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[6] ), .QN(\dp/n532 ) );
  DFFR_X1 \dp/ir_reg[7]  ( .D(\dp/n656 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[7] ), .QN(\dp/n533 ) );
  DFFR_X1 \dp/ir_reg[8]  ( .D(\dp/n657 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[8] ), .QN(\dp/n534 ) );
  DFFR_X1 \dp/ir_reg[9]  ( .D(\dp/n658 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[9] ), .QN(\dp/n535 ) );
  DFFR_X1 \dp/ir_reg[10]  ( .D(\dp/n659 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[10] ), .QN(\dp/n536 ) );
  DFFR_X1 \dp/ir_reg[11]  ( .D(\dp/n660 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[11] ), .QN(\dp/n575 ) );
  DFFR_X1 \dp/ir_reg[12]  ( .D(\dp/n661 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[12] ), .QN(\dp/n577 ) );
  DFFR_X1 \dp/ir_reg[13]  ( .D(\dp/n662 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[13] ), .QN(\dp/n579 ) );
  DFFR_X1 \dp/ir_reg[14]  ( .D(\dp/n663 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[14] ), .QN(\dp/n581 ) );
  DFFR_X1 \dp/ir_reg[15]  ( .D(\dp/n664 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[15] ), .QN(\dp/n583 ) );
  DFFR_X1 \dp/ir_reg[16]  ( .D(\dp/n665 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[16] ), .QN(\dp/n574 ) );
  DFFR_X1 \dp/ir_reg[17]  ( .D(\dp/n666 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[17] ), .QN(\dp/n576 ) );
  DFFR_X1 \dp/ir_reg[18]  ( .D(\dp/n667 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[18] ), .QN(\dp/n578 ) );
  DFFR_X1 \dp/ir_reg[19]  ( .D(\dp/n668 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[19] ), .QN(\dp/n580 ) );
  DFFR_X1 \dp/ir_reg[20]  ( .D(\dp/n669 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[20] ), .QN(\dp/n582 ) );
  DFFR_X1 \dp/ir_reg[21]  ( .D(\dp/n670 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[21] ), .QN(\dp/n537 ) );
  DFFR_X1 \dp/ir_reg[22]  ( .D(\dp/n671 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[22] ), .QN(\dp/n538 ) );
  DFFR_X1 \dp/ir_reg[23]  ( .D(\dp/n672 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[23] ), .QN(\dp/n539 ) );
  DFFR_X1 \dp/ir_reg[24]  ( .D(\dp/n673 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[24] ), .QN(\dp/n540 ) );
  DFFR_X1 \dp/ir_reg[25]  ( .D(\dp/n674 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/ir[25] ), .QN(\dp/n541 ) );
  DFFR_X1 \dp/npc_id_i_reg[0]  ( .D(\dp/n675 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [0]), .QN(\dp/n542 ) );
  DFFR_X1 \dp/npc_id_i_reg[1]  ( .D(\dp/n676 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [1]), .QN(\dp/n543 ) );
  DFFR_X1 \dp/npc_id_i_reg[2]  ( .D(\dp/n677 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [2]), .QN(\dp/n544 ) );
  DFFR_X1 \dp/npc_id_i_reg[3]  ( .D(\dp/n678 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [3]), .QN(\dp/n545 ) );
  DFFR_X1 \dp/npc_id_i_reg[4]  ( .D(\dp/n679 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [4]), .QN(\dp/n546 ) );
  DFFR_X1 \dp/npc_id_i_reg[5]  ( .D(\dp/n680 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [5]), .QN(\dp/n547 ) );
  DFFR_X1 \dp/npc_id_i_reg[6]  ( .D(\dp/n681 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [6]), .QN(\dp/n548 ) );
  DFFR_X1 \dp/npc_id_i_reg[7]  ( .D(\dp/n682 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [7]), .QN(\dp/n549 ) );
  DFFR_X1 \dp/npc_id_i_reg[8]  ( .D(\dp/n683 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [8]), .QN(\dp/n550 ) );
  DFFR_X1 \dp/npc_id_i_reg[9]  ( .D(\dp/n684 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [9]), .QN(\dp/n551 ) );
  DFFR_X1 \dp/npc_id_i_reg[10]  ( .D(\dp/n685 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [10]), .QN(\dp/n552 ) );
  DFFR_X1 \dp/npc_id_i_reg[11]  ( .D(\dp/n686 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_id_o [11]), .QN(\dp/n553 ) );
  DFFR_X1 \dp/rf_out1_ex_i_reg[31]  ( .D(\dp/n844 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rf_out1_ex_i [31]), .QN(\dp/n514 ) );
  DFFR_X1 \dp/branch_t_mem_i_reg  ( .D(\dp/n845 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(is_zero_i), .QN(\dp/n515 ) );
  DFFR_X1 \dp/rd_fwd_wb_i_reg[0]  ( .D(\dp/n1009 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_wb_i [0]), .QN(\dp/n516 ) );
  DFFR_X1 \dp/rd_fwd_wb_i_reg[1]  ( .D(\dp/n1008 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_wb_i [1]), .QN(\dp/n518 ) );
  DFFR_X1 \dp/rd_fwd_wb_i_reg[2]  ( .D(\dp/n1007 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_wb_i [2]), .QN(\dp/n520 ) );
  DFFR_X1 \dp/rd_fwd_wb_i_reg[3]  ( .D(\dp/n1006 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_wb_i [3]), .QN(\dp/n522 ) );
  DFFR_X1 \dp/rd_fwd_wb_i_reg[4]  ( .D(\dp/n1005 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(\dp/rd_fwd_wb_i [4]), .QN(\dp/n524 ) );
  DFFR_X1 \dp/data_mem_mem_i_reg[10]  ( .D(\dp/n994 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[10]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[11]  ( .D(\dp/n993 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[11]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[12]  ( .D(\dp/n992 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[12]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[13]  ( .D(\dp/n991 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[13]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[14]  ( .D(\dp/n990 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[14]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[15]  ( .D(\dp/n989 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[15]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[16]  ( .D(\dp/n988 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[16]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[17]  ( .D(\dp/n987 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[17]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[18]  ( .D(\dp/n986 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[18]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[19]  ( .D(\dp/n985 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[19]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[20]  ( .D(\dp/n984 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[20]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[21]  ( .D(\dp/n983 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[21]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[22]  ( .D(\dp/n982 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[22]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[23]  ( .D(\dp/n981 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[23]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[24]  ( .D(\dp/n980 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[24]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[25]  ( .D(\dp/n979 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[25]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[26]  ( .D(\dp/n978 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[26]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[27]  ( .D(\dp/n977 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[27]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[28]  ( .D(\dp/n976 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[28]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[29]  ( .D(\dp/n975 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[29]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[30]  ( .D(\dp/n974 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[30]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[31]  ( .D(\dp/n973 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[31]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[8]  ( .D(\dp/n996 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_DATA[8]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[9]  ( .D(\dp/n995 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_DATA[9]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[0]  ( .D(\dp/n1004 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[0]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[1]  ( .D(\dp/n1003 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[1]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[2]  ( .D(\dp/n1002 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[2]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[3]  ( .D(\dp/n1001 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[3]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[4]  ( .D(\dp/n1000 ), .CK(CLK), .RN(\dp/n634 ), .Q(DRAM_DATA[4]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[5]  ( .D(\dp/n999 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_DATA[5]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[6]  ( .D(\dp/n998 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_DATA[6]) );
  DFFR_X1 \dp/data_mem_mem_i_reg[7]  ( .D(\dp/n997 ), .CK(CLK), .RN(\dp/n634 ), 
        .Q(DRAM_DATA[7]) );
  DFFR_X1 \dp/npc_ex_i_reg[0]  ( .D(\dp/n717 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [0]), .QN(\dp/n230 ) );
  DFFR_X1 \dp/npc_ex_i_reg[1]  ( .D(\dp/n718 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [1]), .QN(\dp/n231 ) );
  DFFR_X1 \dp/npc_ex_i_reg[2]  ( .D(\dp/n719 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [2]), .QN(\dp/n232 ) );
  DFFR_X1 \dp/npc_ex_i_reg[3]  ( .D(\dp/n720 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [3]), .QN(\dp/n233 ) );
  DFFR_X1 \dp/npc_ex_i_reg[4]  ( .D(\dp/n721 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [4]), .QN(\dp/n234 ) );
  DFFR_X1 \dp/npc_ex_i_reg[5]  ( .D(\dp/n722 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [5]), .QN(\dp/n235 ) );
  DFFR_X1 \dp/npc_ex_i_reg[6]  ( .D(\dp/n723 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [6]), .QN(\dp/n236 ) );
  DFFR_X1 \dp/npc_ex_i_reg[7]  ( .D(\dp/n724 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [7]), .QN(\dp/n237 ) );
  DFFR_X1 \dp/npc_ex_i_reg[8]  ( .D(\dp/n725 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [8]), .QN(\dp/n238 ) );
  DFFR_X1 \dp/npc_ex_i_reg[9]  ( .D(\dp/n726 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [9]), .QN(\dp/n239 ) );
  DFFR_X1 \dp/npc_ex_i_reg[10]  ( .D(\dp/n727 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [10]), .QN(\dp/n240 ) );
  DFFR_X1 \dp/npc_ex_i_reg[11]  ( .D(\dp/n728 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [11]), .QN(\dp/n241 ) );
  DFFR_X1 \dp/npc_ex_i_reg[12]  ( .D(\dp/n729 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [12]), .QN(\dp/n242 ) );
  DFFR_X1 \dp/npc_ex_i_reg[13]  ( .D(\dp/n730 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [13]), .QN(\dp/n243 ) );
  DFFR_X1 \dp/npc_ex_i_reg[14]  ( .D(\dp/n731 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [14]), .QN(\dp/n244 ) );
  DFFR_X1 \dp/npc_ex_i_reg[15]  ( .D(\dp/n732 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [15]), .QN(\dp/n245 ) );
  DFFR_X1 \dp/npc_ex_i_reg[16]  ( .D(\dp/n733 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [16]), .QN(\dp/n246 ) );
  DFFR_X1 \dp/npc_ex_i_reg[17]  ( .D(\dp/n734 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [17]), .QN(\dp/n247 ) );
  DFFR_X1 \dp/npc_ex_i_reg[18]  ( .D(\dp/n735 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [18]), .QN(\dp/n248 ) );
  DFFR_X1 \dp/npc_ex_i_reg[19]  ( .D(\dp/n736 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [19]), .QN(\dp/n249 ) );
  DFFR_X1 \dp/npc_ex_i_reg[20]  ( .D(\dp/n737 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [20]), .QN(\dp/n250 ) );
  DFFR_X1 \dp/npc_ex_i_reg[21]  ( .D(\dp/n738 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [21]), .QN(\dp/n251 ) );
  DFFR_X1 \dp/npc_ex_i_reg[22]  ( .D(\dp/n739 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [22]), .QN(\dp/n252 ) );
  DFFR_X1 \dp/npc_ex_i_reg[23]  ( .D(\dp/n740 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [23]), .QN(\dp/n253 ) );
  DFFR_X1 \dp/npc_ex_i_reg[24]  ( .D(\dp/n741 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [24]), .QN(\dp/n254 ) );
  DFFR_X1 \dp/npc_ex_i_reg[25]  ( .D(\dp/n742 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [25]), .QN(\dp/n255 ) );
  DFFR_X1 \dp/npc_ex_i_reg[26]  ( .D(\dp/n743 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [26]), .QN(\dp/n256 ) );
  DFFR_X1 \dp/npc_ex_i_reg[27]  ( .D(\dp/n744 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [27]), .QN(\dp/n257 ) );
  DFFR_X1 \dp/npc_ex_i_reg[28]  ( .D(\dp/n745 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [28]), .QN(\dp/n258 ) );
  DFFR_X1 \dp/npc_ex_i_reg[29]  ( .D(\dp/n746 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [29]), .QN(\dp/n259 ) );
  DFFR_X1 \dp/npc_ex_i_reg[30]  ( .D(\dp/n747 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [30]), .QN(\dp/n260 ) );
  DFFR_X1 \dp/npc_ex_i_reg[31]  ( .D(\dp/n748 ), .CK(CLK), .RN(\dp/n634 ), .Q(
        \dp/npc_ex_i [31]), .QN(\dp/n261 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[0]  ( .D(\dp/n909 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n303 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[1]  ( .D(\dp/n908 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n304 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[2]  ( .D(\dp/n907 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n305 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[3]  ( .D(\dp/n906 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n306 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[4]  ( .D(\dp/n905 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n307 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[5]  ( .D(\dp/n904 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n308 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[6]  ( .D(\dp/n903 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n309 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[7]  ( .D(\dp/n902 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n310 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[8]  ( .D(\dp/n901 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n311 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[9]  ( .D(\dp/n900 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n312 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[10]  ( .D(\dp/n899 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n313 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[11]  ( .D(\dp/n898 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n314 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[12]  ( .D(\dp/n897 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n315 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[13]  ( .D(\dp/n896 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n316 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[14]  ( .D(\dp/n895 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n317 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[15]  ( .D(\dp/n894 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n318 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[16]  ( .D(\dp/n893 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n319 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[17]  ( .D(\dp/n892 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n320 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[18]  ( .D(\dp/n891 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n321 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[19]  ( .D(\dp/n890 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n322 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[20]  ( .D(\dp/n889 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n323 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[21]  ( .D(\dp/n888 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n324 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[22]  ( .D(\dp/n887 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n325 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[23]  ( .D(\dp/n886 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n326 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[24]  ( .D(\dp/n885 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n327 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[25]  ( .D(\dp/n884 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n328 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[26]  ( .D(\dp/n883 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n329 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[27]  ( .D(\dp/n882 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n330 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[28]  ( .D(\dp/n881 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n331 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[29]  ( .D(\dp/n880 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n332 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[30]  ( .D(\dp/n879 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n333 ) );
  DFFR_X1 \dp/alu_out_wb_i_reg[31]  ( .D(\dp/n878 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n630 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[4]  ( .D(\dp/n969 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n272 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[5]  ( .D(\dp/n968 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n273 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[6]  ( .D(\dp/n967 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n274 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[7]  ( .D(\dp/n966 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n275 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[8]  ( .D(\dp/n965 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n276 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[9]  ( .D(\dp/n964 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n277 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[10]  ( .D(\dp/n963 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n278 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[11]  ( .D(\dp/n962 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n279 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[12]  ( .D(\dp/n961 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n280 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[13]  ( .D(\dp/n960 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n281 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[14]  ( .D(\dp/n959 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n282 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[15]  ( .D(\dp/n958 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n283 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[16]  ( .D(\dp/n957 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n284 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[17]  ( .D(\dp/n956 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n285 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[18]  ( .D(\dp/n955 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n286 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[19]  ( .D(\dp/n954 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n287 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[20]  ( .D(\dp/n953 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n288 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[21]  ( .D(\dp/n952 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n289 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[22]  ( .D(\dp/n951 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n290 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[23]  ( .D(\dp/n950 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n291 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[24]  ( .D(\dp/n949 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n292 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[25]  ( .D(\dp/n948 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n293 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[26]  ( .D(\dp/n947 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n294 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[27]  ( .D(\dp/n946 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n295 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[28]  ( .D(\dp/n945 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n296 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[29]  ( .D(\dp/n944 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n297 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[30]  ( .D(\dp/n943 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n299 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[31]  ( .D(\dp/n942 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n300 ) );
  DFFR_X1 \dp/rd_fwd_mem_i_reg[0]  ( .D(\dp/n1014 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n264 ) );
  DFFR_X1 \dp/rd_fwd_mem_i_reg[1]  ( .D(\dp/n1013 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n265 ) );
  DFFR_X1 \dp/rd_fwd_mem_i_reg[2]  ( .D(\dp/n1012 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n266 ) );
  DFFR_X1 \dp/rd_fwd_mem_i_reg[3]  ( .D(\dp/n1011 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n267 ) );
  DFFR_X1 \dp/rd_fwd_mem_i_reg[4]  ( .D(\dp/n1010 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n268 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[0]  ( .D(\dp/n1015 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n224 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[1]  ( .D(\dp/n972 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n269 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[2]  ( .D(\dp/n971 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n270 ) );
  DFFR_X1 \dp/data_mem_wb_i_reg[3]  ( .D(\dp/n970 ), .CK(CLK), .RN(\dp/n634 ), 
        .QN(\dp/n271 ) );
  TBUF_X1 \dp/z_word_tri[31]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [31]) );
  TBUF_X1 \dp/z_word_tri[30]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [30]) );
  TBUF_X1 \dp/z_word_tri[29]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [29]) );
  TBUF_X1 \dp/z_word_tri[28]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [28]) );
  TBUF_X1 \dp/z_word_tri[27]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [27]) );
  TBUF_X1 \dp/z_word_tri[26]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [26]) );
  TBUF_X1 \dp/z_word_tri[25]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [25]) );
  TBUF_X1 \dp/z_word_tri[24]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [24]) );
  TBUF_X1 \dp/z_word_tri[23]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [23]) );
  TBUF_X1 \dp/z_word_tri[22]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [22]) );
  TBUF_X1 \dp/z_word_tri[21]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [21]) );
  TBUF_X1 \dp/z_word_tri[20]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [20]) );
  TBUF_X1 \dp/z_word_tri[19]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [19]) );
  TBUF_X1 \dp/z_word_tri[18]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [18]) );
  TBUF_X1 \dp/z_word_tri[17]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [17]) );
  TBUF_X1 \dp/z_word_tri[16]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [16]) );
  TBUF_X1 \dp/z_word_tri[15]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [15]) );
  TBUF_X1 \dp/z_word_tri[14]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [14]) );
  TBUF_X1 \dp/z_word_tri[13]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [13]) );
  TBUF_X1 \dp/z_word_tri[12]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [12]) );
  TBUF_X1 \dp/z_word_tri[11]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [11]) );
  TBUF_X1 \dp/z_word_tri[10]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [10]) );
  TBUF_X1 \dp/z_word_tri[9]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [9]) );
  TBUF_X1 \dp/z_word_tri[8]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [8]) );
  TBUF_X1 \dp/z_word_tri[7]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [7]) );
  TBUF_X1 \dp/z_word_tri[6]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [6]) );
  TBUF_X1 \dp/z_word_tri[5]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [5]) );
  TBUF_X1 \dp/z_word_tri[4]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [4]) );
  TBUF_X1 \dp/z_word_tri[3]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [3]) );
  TBUF_X1 \dp/z_word_tri[2]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [2]) );
  TBUF_X1 \dp/z_word_tri[1]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [1]) );
  TBUF_X1 \dp/z_word_tri[0]  ( .A(1'b0), .EN(1'b1), .Z(\dp/z_word [0]) );
  NAND3_X1 \dp/U753  ( .A1(\dp/n9 ), .A2(\dp/n632 ), .A3(npc_wb_en_i), .ZN(
        \dp/n366 ) );
  CLKBUF_X1 \dp/if_stage/U74  ( .A(pc_latch_en_i), .Z(\dp/if_stage/n103 ) );
  CLKBUF_X1 \dp/if_stage/U73  ( .A(pc_latch_en_i), .Z(\dp/if_stage/n102 ) );
  CLKBUF_X1 \dp/if_stage/U72  ( .A(pc_latch_en_i), .Z(\dp/if_stage/n101 ) );
  CLKBUF_X1 \dp/if_stage/U71  ( .A(pc_latch_en_i), .Z(\dp/if_stage/n100 ) );
  CLKBUF_X1 \dp/if_stage/U70  ( .A(pc_latch_en_i), .Z(\dp/if_stage/n99 ) );
  CLKBUF_X1 \dp/if_stage/U69  ( .A(pc_latch_en_i), .Z(\dp/if_stage/n96 ) );
  NAND2_X1 \dp/if_stage/U67  ( .A1(\dp/npc_if_o [0]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n32 ) );
  OAI21_X1 \dp/if_stage/U66  ( .B1(\dp/if_stage/n64 ), .B2(\dp/if_stage/n103 ), 
        .A(\dp/if_stage/n32 ), .ZN(\dp/if_stage/n97 ) );
  NAND2_X1 \dp/if_stage/U65  ( .A1(\dp/npc_if_o [1]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n31 ) );
  OAI21_X1 \dp/if_stage/U64  ( .B1(\dp/if_stage/n63 ), .B2(\dp/if_stage/n103 ), 
        .A(\dp/if_stage/n31 ), .ZN(\dp/if_stage/n95 ) );
  NAND2_X1 \dp/if_stage/U63  ( .A1(\dp/npc_if_o [2]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n30 ) );
  OAI21_X1 \dp/if_stage/U62  ( .B1(\dp/if_stage/n62 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n30 ), .ZN(\dp/if_stage/n94 ) );
  NAND2_X1 \dp/if_stage/U61  ( .A1(\dp/npc_if_o [3]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n29 ) );
  OAI21_X1 \dp/if_stage/U60  ( .B1(\dp/if_stage/n61 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n29 ), .ZN(\dp/if_stage/n93 ) );
  NAND2_X1 \dp/if_stage/U59  ( .A1(\dp/npc_if_o [4]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n28 ) );
  OAI21_X1 \dp/if_stage/U58  ( .B1(\dp/if_stage/n60 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n28 ), .ZN(\dp/if_stage/n92 ) );
  NAND2_X1 \dp/if_stage/U57  ( .A1(\dp/npc_if_o [5]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n27 ) );
  OAI21_X1 \dp/if_stage/U56  ( .B1(\dp/if_stage/n59 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n27 ), .ZN(\dp/if_stage/n91 ) );
  NAND2_X1 \dp/if_stage/U55  ( .A1(\dp/npc_if_o [6]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n26 ) );
  OAI21_X1 \dp/if_stage/U54  ( .B1(\dp/if_stage/n58 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n26 ), .ZN(\dp/if_stage/n90 ) );
  NAND2_X1 \dp/if_stage/U53  ( .A1(\dp/npc_if_o [7]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n25 ) );
  OAI21_X1 \dp/if_stage/U52  ( .B1(\dp/if_stage/n57 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n25 ), .ZN(\dp/if_stage/n89 ) );
  NAND2_X1 \dp/if_stage/U51  ( .A1(\dp/npc_if_o [8]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n24 ) );
  OAI21_X1 \dp/if_stage/U50  ( .B1(\dp/if_stage/n56 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n24 ), .ZN(\dp/if_stage/n88 ) );
  NAND2_X1 \dp/if_stage/U49  ( .A1(\dp/npc_if_o [9]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n23 ) );
  OAI21_X1 \dp/if_stage/U48  ( .B1(\dp/if_stage/n55 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n23 ), .ZN(\dp/if_stage/n87 ) );
  NAND2_X1 \dp/if_stage/U47  ( .A1(\dp/npc_if_o [10]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n22 ) );
  OAI21_X1 \dp/if_stage/U46  ( .B1(\dp/if_stage/n54 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n22 ), .ZN(\dp/if_stage/n86 ) );
  NAND2_X1 \dp/if_stage/U45  ( .A1(\dp/npc_if_o [11]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n21 ) );
  OAI21_X1 \dp/if_stage/U44  ( .B1(\dp/if_stage/n53 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n21 ), .ZN(\dp/if_stage/n85 ) );
  NAND2_X1 \dp/if_stage/U43  ( .A1(\dp/npc_if_o [12]), .A2(\dp/if_stage/n96 ), 
        .ZN(\dp/if_stage/n20 ) );
  OAI21_X1 \dp/if_stage/U42  ( .B1(\dp/if_stage/n52 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n20 ), .ZN(\dp/if_stage/n84 ) );
  NAND2_X1 \dp/if_stage/U41  ( .A1(\dp/npc_if_o [13]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n19 ) );
  OAI21_X1 \dp/if_stage/U40  ( .B1(\dp/if_stage/n51 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n19 ), .ZN(\dp/if_stage/n83 ) );
  NAND2_X1 \dp/if_stage/U39  ( .A1(\dp/npc_if_o [14]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n18 ) );
  OAI21_X1 \dp/if_stage/U38  ( .B1(\dp/if_stage/n50 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n18 ), .ZN(\dp/if_stage/n82 ) );
  NAND2_X1 \dp/if_stage/U37  ( .A1(\dp/npc_if_o [15]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n17 ) );
  OAI21_X1 \dp/if_stage/U36  ( .B1(\dp/if_stage/n49 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n17 ), .ZN(\dp/if_stage/n81 ) );
  NAND2_X1 \dp/if_stage/U35  ( .A1(\dp/npc_if_o [16]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n16 ) );
  OAI21_X1 \dp/if_stage/U34  ( .B1(\dp/if_stage/n48 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n16 ), .ZN(\dp/if_stage/n80 ) );
  NAND2_X1 \dp/if_stage/U33  ( .A1(\dp/npc_if_o [17]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n15 ) );
  OAI21_X1 \dp/if_stage/U32  ( .B1(\dp/if_stage/n47 ), .B2(\dp/if_stage/n100 ), 
        .A(\dp/if_stage/n15 ), .ZN(\dp/if_stage/n79 ) );
  NAND2_X1 \dp/if_stage/U31  ( .A1(\dp/npc_if_o [18]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n14 ) );
  OAI21_X1 \dp/if_stage/U30  ( .B1(\dp/if_stage/n46 ), .B2(\dp/if_stage/n100 ), 
        .A(\dp/if_stage/n14 ), .ZN(\dp/if_stage/n78 ) );
  NAND2_X1 \dp/if_stage/U29  ( .A1(\dp/npc_if_o [19]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n13 ) );
  OAI21_X1 \dp/if_stage/U28  ( .B1(\dp/if_stage/n45 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n13 ), .ZN(\dp/if_stage/n77 ) );
  NAND2_X1 \dp/if_stage/U27  ( .A1(\dp/npc_if_o [23]), .A2(\dp/if_stage/n100 ), 
        .ZN(\dp/if_stage/n9 ) );
  OAI21_X1 \dp/if_stage/U26  ( .B1(\dp/if_stage/n41 ), .B2(\dp/if_stage/n100 ), 
        .A(\dp/if_stage/n9 ), .ZN(\dp/if_stage/n73 ) );
  NAND2_X1 \dp/if_stage/U25  ( .A1(\dp/npc_if_o [25]), .A2(\dp/if_stage/n100 ), 
        .ZN(\dp/if_stage/n7 ) );
  OAI21_X1 \dp/if_stage/U24  ( .B1(\dp/if_stage/n39 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n7 ), .ZN(\dp/if_stage/n71 ) );
  NAND2_X1 \dp/if_stage/U23  ( .A1(\dp/npc_if_o [26]), .A2(\dp/if_stage/n100 ), 
        .ZN(\dp/if_stage/n6 ) );
  OAI21_X1 \dp/if_stage/U22  ( .B1(\dp/if_stage/n38 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n6 ), .ZN(\dp/if_stage/n70 ) );
  NAND2_X1 \dp/if_stage/U21  ( .A1(\dp/npc_if_o [27]), .A2(\dp/if_stage/n100 ), 
        .ZN(\dp/if_stage/n5 ) );
  OAI21_X1 \dp/if_stage/U20  ( .B1(\dp/if_stage/n37 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n5 ), .ZN(\dp/if_stage/n69 ) );
  NAND2_X1 \dp/if_stage/U19  ( .A1(\dp/npc_if_o [28]), .A2(\dp/if_stage/n100 ), 
        .ZN(\dp/if_stage/n4 ) );
  OAI21_X1 \dp/if_stage/U18  ( .B1(\dp/if_stage/n36 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n4 ), .ZN(\dp/if_stage/n68 ) );
  NAND2_X1 \dp/if_stage/U17  ( .A1(\dp/npc_if_o [29]), .A2(\dp/if_stage/n100 ), 
        .ZN(\dp/if_stage/n3 ) );
  OAI21_X1 \dp/if_stage/U16  ( .B1(\dp/if_stage/n35 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n3 ), .ZN(\dp/if_stage/n67 ) );
  NAND2_X1 \dp/if_stage/U15  ( .A1(\dp/npc_if_o [30]), .A2(\dp/if_stage/n100 ), 
        .ZN(\dp/if_stage/n2 ) );
  OAI21_X1 \dp/if_stage/U14  ( .B1(\dp/if_stage/n34 ), .B2(\dp/if_stage/n102 ), 
        .A(\dp/if_stage/n2 ), .ZN(\dp/if_stage/n66 ) );
  NAND2_X1 \dp/if_stage/U13  ( .A1(\dp/npc_if_o [20]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n12 ) );
  OAI21_X1 \dp/if_stage/U12  ( .B1(\dp/if_stage/n44 ), .B2(\dp/if_stage/n100 ), 
        .A(\dp/if_stage/n12 ), .ZN(\dp/if_stage/n76 ) );
  NAND2_X1 \dp/if_stage/U11  ( .A1(\dp/npc_if_o [21]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n11 ) );
  OAI21_X1 \dp/if_stage/U10  ( .B1(\dp/if_stage/n43 ), .B2(\dp/if_stage/n100 ), 
        .A(\dp/if_stage/n11 ), .ZN(\dp/if_stage/n75 ) );
  NAND2_X1 \dp/if_stage/U9  ( .A1(\dp/npc_if_o [22]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n10 ) );
  OAI21_X1 \dp/if_stage/U8  ( .B1(\dp/if_stage/n42 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n10 ), .ZN(\dp/if_stage/n74 ) );
  NAND2_X1 \dp/if_stage/U7  ( .A1(\dp/npc_if_o [24]), .A2(\dp/if_stage/n99 ), 
        .ZN(\dp/if_stage/n8 ) );
  OAI21_X1 \dp/if_stage/U6  ( .B1(\dp/if_stage/n40 ), .B2(\dp/if_stage/n101 ), 
        .A(\dp/if_stage/n8 ), .ZN(\dp/if_stage/n72 ) );
  NAND2_X1 \dp/if_stage/U5  ( .A1(\dp/if_stage/n103 ), .A2(\dp/npc_if_o [31]), 
        .ZN(\dp/if_stage/n1 ) );
  OAI21_X1 \dp/if_stage/U4  ( .B1(\dp/if_stage/n33 ), .B2(\dp/if_stage/n103 ), 
        .A(\dp/if_stage/n1 ), .ZN(\dp/if_stage/n65 ) );
  INV_X2 \dp/if_stage/U3  ( .A(RST), .ZN(\dp/if_stage/n104 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[31]  ( .D(\dp/if_stage/n65 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[31]), .QN(\dp/if_stage/n33 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[30]  ( .D(\dp/if_stage/n66 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[30]), .QN(\dp/if_stage/n34 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[29]  ( .D(\dp/if_stage/n67 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[29]), .QN(\dp/if_stage/n35 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[28]  ( .D(\dp/if_stage/n68 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[28]), .QN(\dp/if_stage/n36 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[27]  ( .D(\dp/if_stage/n69 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[27]), .QN(\dp/if_stage/n37 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[26]  ( .D(\dp/if_stage/n70 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[26]), .QN(\dp/if_stage/n38 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[25]  ( .D(\dp/if_stage/n71 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[25]), .QN(\dp/if_stage/n39 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[24]  ( .D(\dp/if_stage/n72 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[24]), .QN(\dp/if_stage/n40 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[23]  ( .D(\dp/if_stage/n73 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[23]), .QN(\dp/if_stage/n41 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[22]  ( .D(\dp/if_stage/n74 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[22]), .QN(\dp/if_stage/n42 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[21]  ( .D(\dp/if_stage/n75 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[21]), .QN(\dp/if_stage/n43 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[20]  ( .D(\dp/if_stage/n76 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[20]), .QN(\dp/if_stage/n44 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[19]  ( .D(\dp/if_stage/n77 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[19]), .QN(\dp/if_stage/n45 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[18]  ( .D(\dp/if_stage/n78 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[18]), .QN(\dp/if_stage/n46 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[17]  ( .D(\dp/if_stage/n79 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[17]), .QN(\dp/if_stage/n47 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[16]  ( .D(\dp/if_stage/n80 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[16]), .QN(\dp/if_stage/n48 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[15]  ( .D(\dp/if_stage/n81 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[15]), .QN(\dp/if_stage/n49 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[14]  ( .D(\dp/if_stage/n82 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[14]), .QN(\dp/if_stage/n50 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[13]  ( .D(\dp/if_stage/n83 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[13]), .QN(\dp/if_stage/n51 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[12]  ( .D(\dp/if_stage/n84 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[12]), .QN(\dp/if_stage/n52 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[11]  ( .D(\dp/if_stage/n85 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[11]), .QN(\dp/if_stage/n53 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[10]  ( .D(\dp/if_stage/n86 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[10]), .QN(\dp/if_stage/n54 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[2]  ( .D(\dp/if_stage/n94 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[2]), .QN(\dp/if_stage/n62 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[0]  ( .D(\dp/if_stage/n97 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(\dp/if_stage/NPC_4_i [0]), .QN(
        \dp/if_stage/n64 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[1]  ( .D(\dp/if_stage/n95 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(\dp/if_stage/NPC_4_i [1]), .QN(
        \dp/if_stage/n63 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[9]  ( .D(\dp/if_stage/n87 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[9]), .QN(\dp/if_stage/n55 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[3]  ( .D(\dp/if_stage/n93 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[3]), .QN(\dp/if_stage/n61 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[4]  ( .D(\dp/if_stage/n92 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[4]), .QN(\dp/if_stage/n60 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[5]  ( .D(\dp/if_stage/n91 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[5]), .QN(\dp/if_stage/n59 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[6]  ( .D(\dp/if_stage/n90 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[6]), .QN(\dp/if_stage/n58 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[7]  ( .D(\dp/if_stage/n89 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[7]), .QN(\dp/if_stage/n57 ) );
  DFFR_X1 \dp/if_stage/PC_i_reg[8]  ( .D(\dp/if_stage/n88 ), .CK(CLK), .RN(
        \dp/if_stage/n104 ), .Q(IRAM_ADDRESS[8]), .QN(\dp/if_stage/n56 ) );
  INV_X1 \dp/if_stage/mux/U78  ( .A(\dp/if_stage/mux/n14 ), .ZN(
        \dp/if_stage/mux/n5 ) );
  AOI22_X1 \dp/if_stage/mux/U77  ( .A1(\dp/if_stage/NPC_4_i [7]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[7]), .B2(\dp/if_stage/mux/n6 ), 
        .ZN(\dp/if_stage/mux/n36 ) );
  INV_X1 \dp/if_stage/mux/U76  ( .A(\dp/if_stage/mux/n36 ), .ZN(
        \dp/npc_if_o [7]) );
  AOI22_X1 \dp/if_stage/mux/U75  ( .A1(\dp/if_stage/NPC_4_i [8]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[8]), .B2(\dp/if_stage/mux/n6 ), 
        .ZN(\dp/if_stage/mux/n35 ) );
  INV_X1 \dp/if_stage/mux/U74  ( .A(\dp/if_stage/mux/n35 ), .ZN(
        \dp/npc_if_o [8]) );
  AOI22_X1 \dp/if_stage/mux/U73  ( .A1(\dp/if_stage/NPC_4_i [0]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[0]), .B2(\dp/if_stage/mux/n13 ), .ZN(\dp/if_stage/mux/n65 ) );
  INV_X1 \dp/if_stage/mux/U72  ( .A(\dp/if_stage/mux/n65 ), .ZN(
        \dp/npc_if_o [0]) );
  AOI22_X1 \dp/if_stage/mux/U71  ( .A1(\dp/if_stage/NPC_4_i [1]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[1]), .B2(\dp/if_stage/mux/n10 ), .ZN(\dp/if_stage/mux/n54 ) );
  INV_X1 \dp/if_stage/mux/U70  ( .A(\dp/if_stage/mux/n54 ), .ZN(
        \dp/npc_if_o [1]) );
  AOI22_X1 \dp/if_stage/mux/U69  ( .A1(\dp/if_stage/NPC_4_i [2]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[2]), .B2(\dp/if_stage/mux/n7 ), 
        .ZN(\dp/if_stage/mux/n43 ) );
  INV_X1 \dp/if_stage/mux/U68  ( .A(\dp/if_stage/mux/n43 ), .ZN(
        \dp/npc_if_o [2]) );
  AOI22_X1 \dp/if_stage/mux/U67  ( .A1(\dp/if_stage/NPC_4_i [3]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[3]), .B2(\dp/if_stage/mux/n7 ), 
        .ZN(\dp/if_stage/mux/n40 ) );
  INV_X1 \dp/if_stage/mux/U66  ( .A(\dp/if_stage/mux/n40 ), .ZN(
        \dp/npc_if_o [3]) );
  AOI22_X1 \dp/if_stage/mux/U65  ( .A1(\dp/if_stage/NPC_4_i [4]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[4]), .B2(\dp/if_stage/mux/n7 ), 
        .ZN(\dp/if_stage/mux/n39 ) );
  INV_X1 \dp/if_stage/mux/U64  ( .A(\dp/if_stage/mux/n39 ), .ZN(
        \dp/npc_if_o [4]) );
  AOI22_X1 \dp/if_stage/mux/U63  ( .A1(\dp/if_stage/NPC_4_i [5]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[5]), .B2(\dp/if_stage/mux/n6 ), 
        .ZN(\dp/if_stage/mux/n38 ) );
  INV_X1 \dp/if_stage/mux/U62  ( .A(\dp/if_stage/mux/n38 ), .ZN(
        \dp/npc_if_o [5]) );
  AOI22_X1 \dp/if_stage/mux/U61  ( .A1(\dp/if_stage/NPC_4_i [6]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[6]), .B2(\dp/if_stage/mux/n6 ), 
        .ZN(\dp/if_stage/mux/n37 ) );
  INV_X1 \dp/if_stage/mux/U60  ( .A(\dp/if_stage/mux/n37 ), .ZN(
        \dp/npc_if_o [6]) );
  AOI22_X1 \dp/if_stage/mux/U59  ( .A1(\dp/if_stage/NPC_4_i [9]), .A2(
        \dp/if_stage/mux/n5 ), .B1(\dp/if_stage/mux/n13 ), .B2(DRAM_ADDRESS[9]), .ZN(\dp/if_stage/mux/n34 ) );
  INV_X1 \dp/if_stage/mux/U58  ( .A(\dp/if_stage/mux/n34 ), .ZN(
        \dp/npc_if_o [9]) );
  AOI22_X1 \dp/if_stage/mux/U57  ( .A1(\dp/if_stage/NPC_4_i [10]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[10]), .B2(
        \dp/if_stage/mux/n13 ), .ZN(\dp/if_stage/mux/n64 ) );
  INV_X1 \dp/if_stage/mux/U56  ( .A(\dp/if_stage/mux/n64 ), .ZN(
        \dp/npc_if_o [10]) );
  AOI22_X1 \dp/if_stage/mux/U55  ( .A1(\dp/if_stage/NPC_4_i [11]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[11]), .B2(
        \dp/if_stage/mux/n13 ), .ZN(\dp/if_stage/mux/n63 ) );
  INV_X1 \dp/if_stage/mux/U54  ( .A(\dp/if_stage/mux/n63 ), .ZN(
        \dp/npc_if_o [11]) );
  AOI22_X1 \dp/if_stage/mux/U53  ( .A1(\dp/if_stage/NPC_4_i [12]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[12]), .B2(
        \dp/if_stage/mux/n12 ), .ZN(\dp/if_stage/mux/n62 ) );
  INV_X1 \dp/if_stage/mux/U52  ( .A(\dp/if_stage/mux/n62 ), .ZN(
        \dp/npc_if_o [12]) );
  AOI22_X1 \dp/if_stage/mux/U51  ( .A1(\dp/if_stage/NPC_4_i [13]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[13]), .B2(
        \dp/if_stage/mux/n12 ), .ZN(\dp/if_stage/mux/n61 ) );
  INV_X1 \dp/if_stage/mux/U50  ( .A(\dp/if_stage/mux/n61 ), .ZN(
        \dp/npc_if_o [13]) );
  AOI22_X1 \dp/if_stage/mux/U49  ( .A1(\dp/if_stage/NPC_4_i [14]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[14]), .B2(
        \dp/if_stage/mux/n12 ), .ZN(\dp/if_stage/mux/n60 ) );
  INV_X1 \dp/if_stage/mux/U48  ( .A(\dp/if_stage/mux/n60 ), .ZN(
        \dp/npc_if_o [14]) );
  AOI22_X1 \dp/if_stage/mux/U47  ( .A1(\dp/if_stage/NPC_4_i [15]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[15]), .B2(
        \dp/if_stage/mux/n12 ), .ZN(\dp/if_stage/mux/n59 ) );
  INV_X1 \dp/if_stage/mux/U46  ( .A(\dp/if_stage/mux/n59 ), .ZN(
        \dp/npc_if_o [15]) );
  AOI22_X1 \dp/if_stage/mux/U45  ( .A1(\dp/if_stage/NPC_4_i [16]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[16]), .B2(
        \dp/if_stage/mux/n11 ), .ZN(\dp/if_stage/mux/n58 ) );
  INV_X1 \dp/if_stage/mux/U44  ( .A(\dp/if_stage/mux/n58 ), .ZN(
        \dp/npc_if_o [16]) );
  AOI22_X1 \dp/if_stage/mux/U43  ( .A1(\dp/if_stage/NPC_4_i [17]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[17]), .B2(
        \dp/if_stage/mux/n11 ), .ZN(\dp/if_stage/mux/n57 ) );
  INV_X1 \dp/if_stage/mux/U42  ( .A(\dp/if_stage/mux/n57 ), .ZN(
        \dp/npc_if_o [17]) );
  AOI22_X1 \dp/if_stage/mux/U41  ( .A1(\dp/if_stage/NPC_4_i [18]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[18]), .B2(
        \dp/if_stage/mux/n11 ), .ZN(\dp/if_stage/mux/n56 ) );
  INV_X1 \dp/if_stage/mux/U40  ( .A(\dp/if_stage/mux/n56 ), .ZN(
        \dp/npc_if_o [18]) );
  AOI22_X1 \dp/if_stage/mux/U39  ( .A1(\dp/if_stage/NPC_4_i [19]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[19]), .B2(
        \dp/if_stage/mux/n11 ), .ZN(\dp/if_stage/mux/n55 ) );
  INV_X1 \dp/if_stage/mux/U38  ( .A(\dp/if_stage/mux/n55 ), .ZN(
        \dp/npc_if_o [19]) );
  AOI22_X1 \dp/if_stage/mux/U37  ( .A1(\dp/if_stage/NPC_4_i [20]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[20]), .B2(
        \dp/if_stage/mux/n10 ), .ZN(\dp/if_stage/mux/n53 ) );
  INV_X1 \dp/if_stage/mux/U36  ( .A(\dp/if_stage/mux/n53 ), .ZN(
        \dp/npc_if_o [20]) );
  AOI22_X1 \dp/if_stage/mux/U35  ( .A1(\dp/if_stage/NPC_4_i [21]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[21]), .B2(
        \dp/if_stage/mux/n10 ), .ZN(\dp/if_stage/mux/n52 ) );
  INV_X1 \dp/if_stage/mux/U34  ( .A(\dp/if_stage/mux/n52 ), .ZN(
        \dp/npc_if_o [21]) );
  AOI22_X1 \dp/if_stage/mux/U33  ( .A1(\dp/if_stage/NPC_4_i [22]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[22]), .B2(\dp/if_stage/mux/n9 ), .ZN(\dp/if_stage/mux/n51 ) );
  INV_X1 \dp/if_stage/mux/U32  ( .A(\dp/if_stage/mux/n51 ), .ZN(
        \dp/npc_if_o [22]) );
  AOI22_X1 \dp/if_stage/mux/U31  ( .A1(\dp/if_stage/NPC_4_i [23]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[23]), .B2(\dp/if_stage/mux/n9 ), .ZN(\dp/if_stage/mux/n50 ) );
  INV_X1 \dp/if_stage/mux/U30  ( .A(\dp/if_stage/mux/n50 ), .ZN(
        \dp/npc_if_o [23]) );
  AOI22_X1 \dp/if_stage/mux/U29  ( .A1(\dp/if_stage/NPC_4_i [24]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[24]), .B2(\dp/if_stage/mux/n9 ), .ZN(\dp/if_stage/mux/n49 ) );
  INV_X1 \dp/if_stage/mux/U28  ( .A(\dp/if_stage/mux/n49 ), .ZN(
        \dp/npc_if_o [24]) );
  AOI22_X1 \dp/if_stage/mux/U27  ( .A1(\dp/if_stage/NPC_4_i [25]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[25]), .B2(\dp/if_stage/mux/n9 ), .ZN(\dp/if_stage/mux/n48 ) );
  INV_X1 \dp/if_stage/mux/U26  ( .A(\dp/if_stage/mux/n48 ), .ZN(
        \dp/npc_if_o [25]) );
  AOI22_X1 \dp/if_stage/mux/U25  ( .A1(\dp/if_stage/NPC_4_i [26]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[26]), .B2(\dp/if_stage/mux/n8 ), .ZN(\dp/if_stage/mux/n47 ) );
  INV_X1 \dp/if_stage/mux/U24  ( .A(\dp/if_stage/mux/n47 ), .ZN(
        \dp/npc_if_o [26]) );
  AOI22_X1 \dp/if_stage/mux/U23  ( .A1(\dp/if_stage/NPC_4_i [27]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[27]), .B2(\dp/if_stage/mux/n8 ), .ZN(\dp/if_stage/mux/n46 ) );
  INV_X1 \dp/if_stage/mux/U22  ( .A(\dp/if_stage/mux/n46 ), .ZN(
        \dp/npc_if_o [27]) );
  AOI22_X1 \dp/if_stage/mux/U21  ( .A1(\dp/if_stage/NPC_4_i [28]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[28]), .B2(\dp/if_stage/mux/n8 ), .ZN(\dp/if_stage/mux/n45 ) );
  INV_X1 \dp/if_stage/mux/U20  ( .A(\dp/if_stage/mux/n45 ), .ZN(
        \dp/npc_if_o [28]) );
  AOI22_X1 \dp/if_stage/mux/U19  ( .A1(\dp/if_stage/NPC_4_i [29]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[29]), .B2(\dp/if_stage/mux/n8 ), .ZN(\dp/if_stage/mux/n44 ) );
  INV_X1 \dp/if_stage/mux/U18  ( .A(\dp/if_stage/mux/n44 ), .ZN(
        \dp/npc_if_o [29]) );
  AOI22_X1 \dp/if_stage/mux/U17  ( .A1(\dp/if_stage/NPC_4_i [30]), .A2(
        \dp/if_stage/mux/n4 ), .B1(DRAM_ADDRESS[30]), .B2(
        \dp/if_stage/mux/n10 ), .ZN(\dp/if_stage/mux/n42 ) );
  INV_X1 \dp/if_stage/mux/U16  ( .A(\dp/if_stage/mux/n42 ), .ZN(
        \dp/npc_if_o [30]) );
  AOI22_X1 \dp/if_stage/mux/U15  ( .A1(\dp/if_stage/NPC_4_i [31]), .A2(
        \dp/if_stage/mux/n5 ), .B1(DRAM_ADDRESS[31]), .B2(\dp/if_stage/mux/n7 ), .ZN(\dp/if_stage/mux/n41 ) );
  INV_X1 \dp/if_stage/mux/U14  ( .A(\dp/if_stage/mux/n41 ), .ZN(
        \dp/npc_if_o [31]) );
  BUF_X1 \dp/if_stage/mux/U13  ( .A(jump_en_i), .Z(\dp/if_stage/mux/n2 ) );
  BUF_X1 \dp/if_stage/mux/U12  ( .A(jump_en_i), .Z(\dp/if_stage/mux/n1 ) );
  BUF_X1 \dp/if_stage/mux/U11  ( .A(jump_en_i), .Z(\dp/if_stage/mux/n3 ) );
  BUF_X1 \dp/if_stage/mux/U10  ( .A(\dp/if_stage/mux/n3 ), .Z(
        \dp/if_stage/mux/n13 ) );
  BUF_X1 \dp/if_stage/mux/U9  ( .A(\dp/if_stage/mux/n3 ), .Z(
        \dp/if_stage/mux/n14 ) );
  BUF_X1 \dp/if_stage/mux/U8  ( .A(\dp/if_stage/mux/n2 ), .Z(
        \dp/if_stage/mux/n10 ) );
  BUF_X1 \dp/if_stage/mux/U7  ( .A(\dp/if_stage/mux/n1 ), .Z(
        \dp/if_stage/mux/n7 ) );
  BUF_X1 \dp/if_stage/mux/U6  ( .A(\dp/if_stage/mux/n1 ), .Z(
        \dp/if_stage/mux/n6 ) );
  BUF_X1 \dp/if_stage/mux/U5  ( .A(\dp/if_stage/mux/n3 ), .Z(
        \dp/if_stage/mux/n12 ) );
  BUF_X1 \dp/if_stage/mux/U4  ( .A(\dp/if_stage/mux/n2 ), .Z(
        \dp/if_stage/mux/n11 ) );
  BUF_X1 \dp/if_stage/mux/U3  ( .A(\dp/if_stage/mux/n2 ), .Z(
        \dp/if_stage/mux/n9 ) );
  BUF_X1 \dp/if_stage/mux/U2  ( .A(\dp/if_stage/mux/n1 ), .Z(
        \dp/if_stage/mux/n8 ) );
  INV_X1 \dp/if_stage/mux/U1  ( .A(\dp/if_stage/mux/n14 ), .ZN(
        \dp/if_stage/mux/n4 ) );
  INV_X1 \dp/if_stage/add_77/U58  ( .A(IRAM_ADDRESS[2]), .ZN(
        \dp/if_stage/NPC_4_i [2]) );
  AND2_X1 \dp/if_stage/add_77/U57  ( .A1(IRAM_ADDRESS[24]), .A2(
        \dp/if_stage/add_77/n30 ), .ZN(\dp/if_stage/add_77/n57 ) );
  AND2_X1 \dp/if_stage/add_77/U56  ( .A1(IRAM_ADDRESS[25]), .A2(
        \dp/if_stage/add_77/n57 ), .ZN(\dp/if_stage/add_77/n56 ) );
  AND2_X1 \dp/if_stage/add_77/U55  ( .A1(IRAM_ADDRESS[26]), .A2(
        \dp/if_stage/add_77/n56 ), .ZN(\dp/if_stage/add_77/n55 ) );
  AND2_X1 \dp/if_stage/add_77/U54  ( .A1(IRAM_ADDRESS[27]), .A2(
        \dp/if_stage/add_77/n55 ), .ZN(\dp/if_stage/add_77/n54 ) );
  AND2_X1 \dp/if_stage/add_77/U53  ( .A1(IRAM_ADDRESS[28]), .A2(
        \dp/if_stage/add_77/n54 ), .ZN(\dp/if_stage/add_77/n53 ) );
  AND2_X1 \dp/if_stage/add_77/U52  ( .A1(IRAM_ADDRESS[29]), .A2(
        \dp/if_stage/add_77/n53 ), .ZN(\dp/if_stage/add_77/n52 ) );
  AND2_X1 \dp/if_stage/add_77/U51  ( .A1(IRAM_ADDRESS[30]), .A2(
        \dp/if_stage/add_77/n52 ), .ZN(\dp/if_stage/add_77/n51 ) );
  AND2_X1 \dp/if_stage/add_77/U50  ( .A1(IRAM_ADDRESS[3]), .A2(IRAM_ADDRESS[2]), .ZN(\dp/if_stage/add_77/n50 ) );
  AND2_X1 \dp/if_stage/add_77/U49  ( .A1(IRAM_ADDRESS[4]), .A2(
        \dp/if_stage/add_77/n50 ), .ZN(\dp/if_stage/add_77/n49 ) );
  AND2_X1 \dp/if_stage/add_77/U48  ( .A1(IRAM_ADDRESS[5]), .A2(
        \dp/if_stage/add_77/n49 ), .ZN(\dp/if_stage/add_77/n48 ) );
  AND2_X1 \dp/if_stage/add_77/U47  ( .A1(IRAM_ADDRESS[6]), .A2(
        \dp/if_stage/add_77/n48 ), .ZN(\dp/if_stage/add_77/n47 ) );
  AND2_X1 \dp/if_stage/add_77/U46  ( .A1(IRAM_ADDRESS[7]), .A2(
        \dp/if_stage/add_77/n47 ), .ZN(\dp/if_stage/add_77/n46 ) );
  AND2_X1 \dp/if_stage/add_77/U45  ( .A1(IRAM_ADDRESS[8]), .A2(
        \dp/if_stage/add_77/n46 ), .ZN(\dp/if_stage/add_77/n45 ) );
  AND2_X1 \dp/if_stage/add_77/U44  ( .A1(IRAM_ADDRESS[9]), .A2(
        \dp/if_stage/add_77/n45 ), .ZN(\dp/if_stage/add_77/n44 ) );
  AND2_X1 \dp/if_stage/add_77/U43  ( .A1(IRAM_ADDRESS[10]), .A2(
        \dp/if_stage/add_77/n44 ), .ZN(\dp/if_stage/add_77/n43 ) );
  AND2_X1 \dp/if_stage/add_77/U42  ( .A1(IRAM_ADDRESS[11]), .A2(
        \dp/if_stage/add_77/n43 ), .ZN(\dp/if_stage/add_77/n42 ) );
  AND2_X1 \dp/if_stage/add_77/U41  ( .A1(IRAM_ADDRESS[12]), .A2(
        \dp/if_stage/add_77/n42 ), .ZN(\dp/if_stage/add_77/n41 ) );
  AND2_X1 \dp/if_stage/add_77/U40  ( .A1(IRAM_ADDRESS[13]), .A2(
        \dp/if_stage/add_77/n41 ), .ZN(\dp/if_stage/add_77/n40 ) );
  AND2_X1 \dp/if_stage/add_77/U39  ( .A1(IRAM_ADDRESS[14]), .A2(
        \dp/if_stage/add_77/n40 ), .ZN(\dp/if_stage/add_77/n39 ) );
  AND2_X1 \dp/if_stage/add_77/U38  ( .A1(IRAM_ADDRESS[15]), .A2(
        \dp/if_stage/add_77/n39 ), .ZN(\dp/if_stage/add_77/n38 ) );
  AND2_X1 \dp/if_stage/add_77/U37  ( .A1(IRAM_ADDRESS[16]), .A2(
        \dp/if_stage/add_77/n38 ), .ZN(\dp/if_stage/add_77/n37 ) );
  AND2_X1 \dp/if_stage/add_77/U36  ( .A1(IRAM_ADDRESS[17]), .A2(
        \dp/if_stage/add_77/n37 ), .ZN(\dp/if_stage/add_77/n36 ) );
  AND2_X1 \dp/if_stage/add_77/U35  ( .A1(IRAM_ADDRESS[18]), .A2(
        \dp/if_stage/add_77/n36 ), .ZN(\dp/if_stage/add_77/n35 ) );
  AND2_X1 \dp/if_stage/add_77/U34  ( .A1(IRAM_ADDRESS[19]), .A2(
        \dp/if_stage/add_77/n35 ), .ZN(\dp/if_stage/add_77/n34 ) );
  AND2_X1 \dp/if_stage/add_77/U33  ( .A1(IRAM_ADDRESS[20]), .A2(
        \dp/if_stage/add_77/n34 ), .ZN(\dp/if_stage/add_77/n33 ) );
  AND2_X1 \dp/if_stage/add_77/U32  ( .A1(IRAM_ADDRESS[21]), .A2(
        \dp/if_stage/add_77/n33 ), .ZN(\dp/if_stage/add_77/n32 ) );
  AND2_X1 \dp/if_stage/add_77/U31  ( .A1(IRAM_ADDRESS[22]), .A2(
        \dp/if_stage/add_77/n32 ), .ZN(\dp/if_stage/add_77/n31 ) );
  AND2_X1 \dp/if_stage/add_77/U30  ( .A1(IRAM_ADDRESS[23]), .A2(
        \dp/if_stage/add_77/n31 ), .ZN(\dp/if_stage/add_77/n30 ) );
  XOR2_X1 \dp/if_stage/add_77/U29  ( .A(IRAM_ADDRESS[7]), .B(
        \dp/if_stage/add_77/n47 ), .Z(\dp/if_stage/NPC_4_i [7]) );
  XOR2_X1 \dp/if_stage/add_77/U28  ( .A(IRAM_ADDRESS[8]), .B(
        \dp/if_stage/add_77/n46 ), .Z(\dp/if_stage/NPC_4_i [8]) );
  XOR2_X1 \dp/if_stage/add_77/U27  ( .A(IRAM_ADDRESS[4]), .B(
        \dp/if_stage/add_77/n50 ), .Z(\dp/if_stage/NPC_4_i [4]) );
  XOR2_X1 \dp/if_stage/add_77/U26  ( .A(IRAM_ADDRESS[5]), .B(
        \dp/if_stage/add_77/n49 ), .Z(\dp/if_stage/NPC_4_i [5]) );
  XOR2_X1 \dp/if_stage/add_77/U25  ( .A(IRAM_ADDRESS[6]), .B(
        \dp/if_stage/add_77/n48 ), .Z(\dp/if_stage/NPC_4_i [6]) );
  XOR2_X1 \dp/if_stage/add_77/U24  ( .A(IRAM_ADDRESS[9]), .B(
        \dp/if_stage/add_77/n45 ), .Z(\dp/if_stage/NPC_4_i [9]) );
  XOR2_X1 \dp/if_stage/add_77/U23  ( .A(IRAM_ADDRESS[10]), .B(
        \dp/if_stage/add_77/n44 ), .Z(\dp/if_stage/NPC_4_i [10]) );
  XOR2_X1 \dp/if_stage/add_77/U22  ( .A(IRAM_ADDRESS[11]), .B(
        \dp/if_stage/add_77/n43 ), .Z(\dp/if_stage/NPC_4_i [11]) );
  XOR2_X1 \dp/if_stage/add_77/U21  ( .A(IRAM_ADDRESS[12]), .B(
        \dp/if_stage/add_77/n42 ), .Z(\dp/if_stage/NPC_4_i [12]) );
  XOR2_X1 \dp/if_stage/add_77/U20  ( .A(IRAM_ADDRESS[13]), .B(
        \dp/if_stage/add_77/n41 ), .Z(\dp/if_stage/NPC_4_i [13]) );
  XOR2_X1 \dp/if_stage/add_77/U19  ( .A(IRAM_ADDRESS[14]), .B(
        \dp/if_stage/add_77/n40 ), .Z(\dp/if_stage/NPC_4_i [14]) );
  XOR2_X1 \dp/if_stage/add_77/U18  ( .A(IRAM_ADDRESS[3]), .B(IRAM_ADDRESS[2]), 
        .Z(\dp/if_stage/NPC_4_i [3]) );
  XOR2_X1 \dp/if_stage/add_77/U17  ( .A(IRAM_ADDRESS[31]), .B(
        \dp/if_stage/add_77/n51 ), .Z(\dp/if_stage/NPC_4_i [31]) );
  XOR2_X1 \dp/if_stage/add_77/U16  ( .A(IRAM_ADDRESS[15]), .B(
        \dp/if_stage/add_77/n39 ), .Z(\dp/if_stage/NPC_4_i [15]) );
  XOR2_X1 \dp/if_stage/add_77/U15  ( .A(IRAM_ADDRESS[16]), .B(
        \dp/if_stage/add_77/n38 ), .Z(\dp/if_stage/NPC_4_i [16]) );
  XOR2_X1 \dp/if_stage/add_77/U14  ( .A(IRAM_ADDRESS[17]), .B(
        \dp/if_stage/add_77/n37 ), .Z(\dp/if_stage/NPC_4_i [17]) );
  XOR2_X1 \dp/if_stage/add_77/U13  ( .A(IRAM_ADDRESS[18]), .B(
        \dp/if_stage/add_77/n36 ), .Z(\dp/if_stage/NPC_4_i [18]) );
  XOR2_X1 \dp/if_stage/add_77/U12  ( .A(IRAM_ADDRESS[19]), .B(
        \dp/if_stage/add_77/n35 ), .Z(\dp/if_stage/NPC_4_i [19]) );
  XOR2_X1 \dp/if_stage/add_77/U11  ( .A(IRAM_ADDRESS[20]), .B(
        \dp/if_stage/add_77/n34 ), .Z(\dp/if_stage/NPC_4_i [20]) );
  XOR2_X1 \dp/if_stage/add_77/U10  ( .A(IRAM_ADDRESS[21]), .B(
        \dp/if_stage/add_77/n33 ), .Z(\dp/if_stage/NPC_4_i [21]) );
  XOR2_X1 \dp/if_stage/add_77/U9  ( .A(IRAM_ADDRESS[22]), .B(
        \dp/if_stage/add_77/n32 ), .Z(\dp/if_stage/NPC_4_i [22]) );
  XOR2_X1 \dp/if_stage/add_77/U8  ( .A(IRAM_ADDRESS[23]), .B(
        \dp/if_stage/add_77/n31 ), .Z(\dp/if_stage/NPC_4_i [23]) );
  XOR2_X1 \dp/if_stage/add_77/U7  ( .A(IRAM_ADDRESS[24]), .B(
        \dp/if_stage/add_77/n30 ), .Z(\dp/if_stage/NPC_4_i [24]) );
  XOR2_X1 \dp/if_stage/add_77/U6  ( .A(IRAM_ADDRESS[25]), .B(
        \dp/if_stage/add_77/n57 ), .Z(\dp/if_stage/NPC_4_i [25]) );
  XOR2_X1 \dp/if_stage/add_77/U5  ( .A(IRAM_ADDRESS[26]), .B(
        \dp/if_stage/add_77/n56 ), .Z(\dp/if_stage/NPC_4_i [26]) );
  XOR2_X1 \dp/if_stage/add_77/U4  ( .A(IRAM_ADDRESS[27]), .B(
        \dp/if_stage/add_77/n55 ), .Z(\dp/if_stage/NPC_4_i [27]) );
  XOR2_X1 \dp/if_stage/add_77/U3  ( .A(IRAM_ADDRESS[28]), .B(
        \dp/if_stage/add_77/n54 ), .Z(\dp/if_stage/NPC_4_i [28]) );
  XOR2_X1 \dp/if_stage/add_77/U2  ( .A(IRAM_ADDRESS[29]), .B(
        \dp/if_stage/add_77/n53 ), .Z(\dp/if_stage/NPC_4_i [29]) );
  XOR2_X1 \dp/if_stage/add_77/U1  ( .A(IRAM_ADDRESS[30]), .B(
        \dp/if_stage/add_77/n52 ), .Z(\dp/if_stage/NPC_4_i [30]) );
  XOR2_X1 \dp/id_stage/U147  ( .A(\dp/rd_fwd_wb_i [4]), .B(\dp/id_stage/n27 ), 
        .Z(\dp/id_stage/p_addr_wRD [4]) );
  NOR2_X1 \dp/id_stage/U146  ( .A1(\dp/rd_fwd_wb_i [3]), .A2(\dp/id_stage/n26 ), .ZN(\dp/id_stage/n27 ) );
  XNOR2_X1 \dp/id_stage/U145  ( .A(\dp/rd_fwd_wb_i [3]), .B(\dp/id_stage/n26 ), 
        .ZN(\dp/id_stage/p_addr_wRD [3]) );
  OAI21_X1 \dp/id_stage/U144  ( .B1(\dp/id_stage/n25 ), .B2(\dp/id_stage/n28 ), 
        .A(\dp/id_stage/n26 ), .ZN(\dp/id_stage/p_addr_wRD [2]) );
  NAND2_X1 \dp/id_stage/U143  ( .A1(\dp/id_stage/n25 ), .A2(\dp/id_stage/n28 ), 
        .ZN(\dp/id_stage/n26 ) );
  AOI21_X1 \dp/id_stage/U142  ( .B1(\dp/rd_fwd_wb_i [0]), .B2(
        \dp/rd_fwd_wb_i [1]), .A(\dp/id_stage/n25 ), .ZN(\dp/id_stage/n24 ) );
  NOR2_X1 \dp/id_stage/U141  ( .A1(\dp/rd_fwd_wb_i [1]), .A2(
        \dp/rd_fwd_wb_i [0]), .ZN(\dp/id_stage/n25 ) );
  XOR2_X1 \dp/id_stage/U140  ( .A(\dp/ir[20] ), .B(\dp/id_stage/n15 ), .Z(
        \dp/id_stage/p_addr_wRS2 [4]) );
  NOR2_X1 \dp/id_stage/U139  ( .A1(\dp/ir[19] ), .A2(\dp/id_stage/n14 ), .ZN(
        \dp/id_stage/n15 ) );
  XNOR2_X1 \dp/id_stage/U138  ( .A(\dp/ir[19] ), .B(\dp/id_stage/n14 ), .ZN(
        \dp/id_stage/p_addr_wRS2 [3]) );
  OAI21_X1 \dp/id_stage/U137  ( .B1(\dp/id_stage/n13 ), .B2(\dp/id_stage/n16 ), 
        .A(\dp/id_stage/n14 ), .ZN(\dp/id_stage/p_addr_wRS2 [2]) );
  NAND2_X1 \dp/id_stage/U136  ( .A1(\dp/id_stage/n13 ), .A2(\dp/id_stage/n16 ), 
        .ZN(\dp/id_stage/n14 ) );
  AOI21_X1 \dp/id_stage/U135  ( .B1(\dp/ir[16] ), .B2(\dp/ir[17] ), .A(
        \dp/id_stage/n13 ), .ZN(\dp/id_stage/n12 ) );
  NOR2_X1 \dp/id_stage/U134  ( .A1(\dp/ir[17] ), .A2(\dp/ir[16] ), .ZN(
        \dp/id_stage/n13 ) );
  XOR2_X1 \dp/id_stage/U133  ( .A(\dp/ir[25] ), .B(\dp/id_stage/n10 ), .Z(
        \dp/id_stage/p_addr_wRS1 [4]) );
  NOR2_X1 \dp/id_stage/U132  ( .A1(\dp/ir[24] ), .A2(\dp/id_stage/n9 ), .ZN(
        \dp/id_stage/n10 ) );
  XNOR2_X1 \dp/id_stage/U131  ( .A(\dp/ir[24] ), .B(\dp/id_stage/n9 ), .ZN(
        \dp/id_stage/p_addr_wRS1 [3]) );
  OAI21_X1 \dp/id_stage/U130  ( .B1(\dp/id_stage/n8 ), .B2(\dp/id_stage/n11 ), 
        .A(\dp/id_stage/n9 ), .ZN(\dp/id_stage/p_addr_wRS1 [2]) );
  NAND2_X1 \dp/id_stage/U129  ( .A1(\dp/id_stage/n8 ), .A2(\dp/id_stage/n11 ), 
        .ZN(\dp/id_stage/n9 ) );
  AOI21_X1 \dp/id_stage/U128  ( .B1(\dp/ir[21] ), .B2(\dp/ir[22] ), .A(
        \dp/id_stage/n8 ), .ZN(\dp/id_stage/n7 ) );
  NOR2_X1 \dp/id_stage/U127  ( .A1(\dp/ir[22] ), .A2(\dp/ir[21] ), .ZN(
        \dp/id_stage/n8 ) );
  INV_X1 \dp/id_stage/U126  ( .A(\dp/ir[23] ), .ZN(\dp/id_stage/n11 ) );
  INV_X1 \dp/id_stage/U125  ( .A(\dp/ir[18] ), .ZN(\dp/id_stage/n16 ) );
  INV_X1 \dp/id_stage/U124  ( .A(\dp/id_stage/n7 ), .ZN(
        \dp/id_stage/p_addr_wRS1 [1]) );
  INV_X1 \dp/id_stage/U123  ( .A(\dp/ir[21] ), .ZN(
        \dp/id_stage/p_addr_wRS1 [0]) );
  INV_X1 \dp/id_stage/U122  ( .A(\dp/id_stage/n12 ), .ZN(
        \dp/id_stage/p_addr_wRS2 [1]) );
  INV_X1 \dp/id_stage/U121  ( .A(\dp/ir[16] ), .ZN(
        \dp/id_stage/p_addr_wRS2 [0]) );
  INV_X1 \dp/id_stage/U120  ( .A(imm_uns_i), .ZN(\dp/id_stage/n39 ) );
  OR3_X1 \dp/id_stage/U119  ( .A1(\dp/ir[20] ), .A2(\dp/ir[19] ), .A3(
        \dp/ir[18] ), .ZN(\dp/id_stage/n18 ) );
  OR3_X1 \dp/id_stage/U118  ( .A1(\dp/ir[17] ), .A2(\dp/ir[16] ), .A3(
        \dp/id_stage/n18 ), .ZN(\dp/id_stage/n17 ) );
  OR3_X1 \dp/id_stage/U117  ( .A1(\dp/ir[25] ), .A2(\dp/ir[24] ), .A3(
        \dp/ir[23] ), .ZN(\dp/id_stage/n20 ) );
  OR3_X1 \dp/id_stage/U116  ( .A1(\dp/ir[22] ), .A2(\dp/ir[21] ), .A3(
        \dp/id_stage/n20 ), .ZN(\dp/id_stage/n19 ) );
  INV_X1 \dp/id_stage/U115  ( .A(\dp/ir[19] ), .ZN(\dp/id_stage/n32 ) );
  OAI21_X1 \dp/id_stage/U114  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n32 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [19]) );
  AND2_X1 \dp/id_stage/U113  ( .A1(\dp/ir[6] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [6]) );
  AND2_X1 \dp/id_stage/U112  ( .A1(\dp/ir[7] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [7]) );
  AND2_X1 \dp/id_stage/U111  ( .A1(\dp/id_stage/n21 ), .A2(\dp/ir[15] ), .ZN(
        \dp/imm_id_o [15]) );
  INV_X1 \dp/id_stage/U110  ( .A(\dp/ir[16] ), .ZN(\dp/id_stage/n29 ) );
  OAI21_X1 \dp/id_stage/U109  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n29 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [16]) );
  INV_X1 \dp/id_stage/U108  ( .A(\dp/ir[17] ), .ZN(\dp/id_stage/n30 ) );
  OAI21_X1 \dp/id_stage/U107  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n30 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [17]) );
  INV_X1 \dp/id_stage/U106  ( .A(\dp/ir[18] ), .ZN(\dp/id_stage/n31 ) );
  OAI21_X1 \dp/id_stage/U105  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n31 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [18]) );
  INV_X1 \dp/id_stage/U104  ( .A(\dp/ir[20] ), .ZN(\dp/id_stage/n33 ) );
  OAI21_X1 \dp/id_stage/U103  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n33 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [20]) );
  INV_X1 \dp/id_stage/U102  ( .A(\dp/ir[21] ), .ZN(\dp/id_stage/n34 ) );
  OAI21_X1 \dp/id_stage/U101  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n34 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [21]) );
  INV_X1 \dp/id_stage/U100  ( .A(\dp/ir[22] ), .ZN(\dp/id_stage/n35 ) );
  OAI21_X1 \dp/id_stage/U99  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n35 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [22]) );
  INV_X1 \dp/id_stage/U98  ( .A(\dp/ir[23] ), .ZN(\dp/id_stage/n36 ) );
  OAI21_X1 \dp/id_stage/U97  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n36 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [23]) );
  INV_X1 \dp/id_stage/U96  ( .A(\dp/ir[24] ), .ZN(\dp/id_stage/n37 ) );
  OAI21_X1 \dp/id_stage/U95  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n37 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [24]) );
  AND2_X1 \dp/id_stage/U94  ( .A1(\dp/ir[0] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [0]) );
  AND2_X1 \dp/id_stage/U93  ( .A1(\dp/ir[1] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [1]) );
  AND2_X1 \dp/id_stage/U92  ( .A1(\dp/ir[2] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [2]) );
  AND2_X1 \dp/id_stage/U91  ( .A1(\dp/ir[3] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [3]) );
  AND2_X1 \dp/id_stage/U90  ( .A1(\dp/ir[4] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [4]) );
  AND2_X1 \dp/id_stage/U89  ( .A1(\dp/ir[5] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [5]) );
  AND2_X1 \dp/id_stage/U88  ( .A1(\dp/ir[8] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [8]) );
  AND2_X1 \dp/id_stage/U87  ( .A1(\dp/ir[9] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [9]) );
  AND2_X1 \dp/id_stage/U86  ( .A1(\dp/ir[10] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [10]) );
  AND2_X1 \dp/id_stage/U85  ( .A1(\dp/ir[11] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [11]) );
  AND2_X1 \dp/id_stage/U84  ( .A1(\dp/ir[12] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [12]) );
  AND2_X1 \dp/id_stage/U83  ( .A1(\dp/ir[13] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [13]) );
  AND2_X1 \dp/id_stage/U82  ( .A1(\dp/ir[14] ), .A2(\dp/id_stage/n21 ), .ZN(
        \dp/imm_id_o [14]) );
  AND2_X1 \dp/id_stage/U81  ( .A1(\dp/id_stage/out2_i [0]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [0]) );
  AND2_X1 \dp/id_stage/U80  ( .A1(\dp/id_stage/out2_i [1]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [1]) );
  AND2_X1 \dp/id_stage/U79  ( .A1(\dp/id_stage/out2_i [2]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [2]) );
  AND2_X1 \dp/id_stage/U78  ( .A1(\dp/id_stage/out2_i [3]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [3]) );
  AND2_X1 \dp/id_stage/U77  ( .A1(\dp/id_stage/out2_i [4]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [4]) );
  AND2_X1 \dp/id_stage/U76  ( .A1(\dp/id_stage/out2_i [5]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [5]) );
  AND2_X1 \dp/id_stage/U75  ( .A1(\dp/id_stage/out2_i [6]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [6]) );
  AND2_X1 \dp/id_stage/U74  ( .A1(\dp/id_stage/out2_i [7]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [7]) );
  AND2_X1 \dp/id_stage/U73  ( .A1(\dp/id_stage/out2_i [8]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [8]) );
  AND2_X1 \dp/id_stage/U72  ( .A1(\dp/id_stage/out2_i [9]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [9]) );
  AND2_X1 \dp/id_stage/U71  ( .A1(\dp/id_stage/out2_i [10]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [10]) );
  AND2_X1 \dp/id_stage/U70  ( .A1(\dp/id_stage/out2_i [11]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [11]) );
  AND2_X1 \dp/id_stage/U69  ( .A1(\dp/id_stage/out2_i [12]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [12]) );
  AND2_X1 \dp/id_stage/U68  ( .A1(\dp/id_stage/out2_i [13]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [13]) );
  AND2_X1 \dp/id_stage/U67  ( .A1(\dp/id_stage/out2_i [14]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [14]) );
  AND2_X1 \dp/id_stage/U66  ( .A1(\dp/id_stage/out2_i [15]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [15]) );
  AND2_X1 \dp/id_stage/U65  ( .A1(\dp/id_stage/out2_i [16]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [16]) );
  AND2_X1 \dp/id_stage/U64  ( .A1(\dp/id_stage/out2_i [17]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [17]) );
  AND2_X1 \dp/id_stage/U63  ( .A1(\dp/id_stage/out2_i [18]), .A2(
        \dp/id_stage/n6 ), .ZN(\dp/rf_out2_id_o [18]) );
  AND2_X1 \dp/id_stage/U62  ( .A1(\dp/id_stage/out2_i [19]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [19]) );
  AND2_X1 \dp/id_stage/U61  ( .A1(\dp/id_stage/out2_i [20]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [20]) );
  AND2_X1 \dp/id_stage/U60  ( .A1(\dp/id_stage/out2_i [21]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [21]) );
  AND2_X1 \dp/id_stage/U59  ( .A1(\dp/id_stage/out2_i [22]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [22]) );
  AND2_X1 \dp/id_stage/U58  ( .A1(\dp/id_stage/out2_i [23]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [23]) );
  AND2_X1 \dp/id_stage/U57  ( .A1(\dp/id_stage/out2_i [24]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [24]) );
  AND2_X1 \dp/id_stage/U56  ( .A1(\dp/id_stage/out2_i [25]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [25]) );
  AND2_X1 \dp/id_stage/U55  ( .A1(\dp/id_stage/out2_i [26]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [26]) );
  AND2_X1 \dp/id_stage/U54  ( .A1(\dp/id_stage/out2_i [27]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [27]) );
  AND2_X1 \dp/id_stage/U53  ( .A1(\dp/id_stage/out2_i [28]), .A2(
        \dp/id_stage/n5 ), .ZN(\dp/rf_out2_id_o [28]) );
  AND2_X1 \dp/id_stage/U52  ( .A1(\dp/id_stage/out2_i [29]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [29]) );
  AND2_X1 \dp/id_stage/U51  ( .A1(\dp/id_stage/out2_i [30]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [30]) );
  AND2_X1 \dp/id_stage/U50  ( .A1(\dp/id_stage/out2_i [31]), .A2(
        \dp/id_stage/n4 ), .ZN(\dp/rf_out2_id_o [31]) );
  AND2_X1 \dp/id_stage/U49  ( .A1(\dp/id_stage/out1_i [0]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [0]) );
  AND2_X1 \dp/id_stage/U48  ( .A1(\dp/id_stage/out1_i [1]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [1]) );
  AND2_X1 \dp/id_stage/U47  ( .A1(\dp/id_stage/out1_i [2]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [2]) );
  AND2_X1 \dp/id_stage/U46  ( .A1(\dp/id_stage/out1_i [3]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [3]) );
  AND2_X1 \dp/id_stage/U45  ( .A1(\dp/id_stage/out1_i [4]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [4]) );
  AND2_X1 \dp/id_stage/U44  ( .A1(\dp/id_stage/out1_i [5]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [5]) );
  AND2_X1 \dp/id_stage/U43  ( .A1(\dp/id_stage/out1_i [6]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [6]) );
  AND2_X1 \dp/id_stage/U42  ( .A1(\dp/id_stage/out1_i [7]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [7]) );
  AND2_X1 \dp/id_stage/U41  ( .A1(\dp/id_stage/out1_i [8]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [8]) );
  AND2_X1 \dp/id_stage/U40  ( .A1(\dp/id_stage/out1_i [9]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [9]) );
  AND2_X1 \dp/id_stage/U39  ( .A1(\dp/id_stage/out1_i [10]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [10]) );
  AND2_X1 \dp/id_stage/U38  ( .A1(\dp/id_stage/out1_i [11]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [11]) );
  AND2_X1 \dp/id_stage/U37  ( .A1(\dp/id_stage/out1_i [12]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [12]) );
  AND2_X1 \dp/id_stage/U36  ( .A1(\dp/id_stage/out1_i [13]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [13]) );
  AND2_X1 \dp/id_stage/U35  ( .A1(\dp/id_stage/out1_i [14]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [14]) );
  AND2_X1 \dp/id_stage/U34  ( .A1(\dp/id_stage/out1_i [15]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [15]) );
  AND2_X1 \dp/id_stage/U33  ( .A1(\dp/id_stage/out1_i [16]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [16]) );
  AND2_X1 \dp/id_stage/U32  ( .A1(\dp/id_stage/out1_i [17]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [17]) );
  AND2_X1 \dp/id_stage/U31  ( .A1(\dp/id_stage/out1_i [18]), .A2(
        \dp/id_stage/n3 ), .ZN(\dp/rf_out1_id_o [18]) );
  AND2_X1 \dp/id_stage/U30  ( .A1(\dp/id_stage/out1_i [19]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [19]) );
  AND2_X1 \dp/id_stage/U29  ( .A1(\dp/id_stage/out1_i [20]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [20]) );
  AND2_X1 \dp/id_stage/U28  ( .A1(\dp/id_stage/out1_i [21]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [21]) );
  AND2_X1 \dp/id_stage/U27  ( .A1(\dp/id_stage/out1_i [22]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [22]) );
  AND2_X1 \dp/id_stage/U26  ( .A1(\dp/id_stage/out1_i [23]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [23]) );
  AND2_X1 \dp/id_stage/U25  ( .A1(\dp/id_stage/out1_i [24]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [24]) );
  AND2_X1 \dp/id_stage/U24  ( .A1(\dp/id_stage/out1_i [25]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [25]) );
  AND2_X1 \dp/id_stage/U23  ( .A1(\dp/id_stage/out1_i [26]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [26]) );
  AND2_X1 \dp/id_stage/U22  ( .A1(\dp/id_stage/out1_i [27]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [27]) );
  AND2_X1 \dp/id_stage/U21  ( .A1(\dp/id_stage/out1_i [28]), .A2(
        \dp/id_stage/n2 ), .ZN(\dp/rf_out1_id_o [28]) );
  AND2_X1 \dp/id_stage/U20  ( .A1(\dp/id_stage/out1_i [29]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [29]) );
  AND2_X1 \dp/id_stage/U19  ( .A1(\dp/id_stage/out1_i [30]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [30]) );
  AND2_X1 \dp/id_stage/U18  ( .A1(\dp/id_stage/out1_i [31]), .A2(
        \dp/id_stage/n1 ), .ZN(\dp/rf_out1_id_o [31]) );
  NAND2_X1 \dp/id_stage/U17  ( .A1(imm_isoff_i), .A2(\dp/id_stage/n22 ), .ZN(
        \dp/id_stage/n21 ) );
  NAND2_X1 \dp/id_stage/U16  ( .A1(imm_isoff_i), .A2(\dp/id_stage/n39 ), .ZN(
        \dp/id_stage/n22 ) );
  INV_X1 \dp/id_stage/U15  ( .A(imm_isoff_i), .ZN(\dp/id_stage/n40 ) );
  NAND3_X1 \dp/id_stage/U14  ( .A1(\dp/id_stage/n40 ), .A2(\dp/id_stage/n39 ), 
        .A3(\dp/ir[15] ), .ZN(\dp/id_stage/n23 ) );
  INV_X1 \dp/id_stage/U13  ( .A(\dp/ir[25] ), .ZN(\dp/id_stage/n38 ) );
  OAI21_X1 \dp/id_stage/U12  ( .B1(\dp/id_stage/n22 ), .B2(\dp/id_stage/n38 ), 
        .A(\dp/id_stage/n23 ), .ZN(\dp/imm_id_o [31]) );
  INV_X1 \dp/id_stage/U11  ( .A(\dp/rd_fwd_wb_i [2]), .ZN(\dp/id_stage/n28 )
         );
  INV_X1 \dp/id_stage/U10  ( .A(\dp/rd_fwd_wb_i [0]), .ZN(
        \dp/id_stage/p_addr_wRD [0]) );
  INV_X1 \dp/id_stage/U9  ( .A(\dp/id_stage/n24 ), .ZN(
        \dp/id_stage/p_addr_wRD [1]) );
  BUF_X1 \dp/id_stage/U8  ( .A(\dp/id_stage/n17 ), .Z(\dp/id_stage/n5 ) );
  BUF_X1 \dp/id_stage/U7  ( .A(\dp/id_stage/n17 ), .Z(\dp/id_stage/n4 ) );
  BUF_X1 \dp/id_stage/U6  ( .A(\dp/id_stage/n19 ), .Z(\dp/id_stage/n2 ) );
  BUF_X1 \dp/id_stage/U5  ( .A(\dp/id_stage/n19 ), .Z(\dp/id_stage/n1 ) );
  BUF_X1 \dp/id_stage/U4  ( .A(\dp/id_stage/n17 ), .Z(\dp/id_stage/n6 ) );
  BUF_X1 \dp/id_stage/U3  ( .A(\dp/id_stage/n19 ), .Z(\dp/id_stage/n3 ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U46  ( .A(1'b0), .ZN(
        \dp/id_stage/regfile/ControlUnit/n15 ) );
  AND2_X1 \dp/id_stage/regfile/ControlUnit/U45  ( .A1(
        \dp/id_stage/regfile/canrestore ), .A2(1'b0), .ZN(
        \dp/id_stage/regfile/ControlUnit/n24 ) );
  OAI22_X1 \dp/id_stage/regfile/ControlUnit/U44  ( .A1(
        \dp/id_stage/regfile/cansave ), .A2(
        \dp/id_stage/regfile/ControlUnit/n15 ), .B1(1'b0), .B2(
        \dp/id_stage/regfile/ControlUnit/n24 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n23 ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U43  ( .A(
        \dp/id_stage/regfile/end_sf ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n16 ) );
  AND3_X1 \dp/id_stage/regfile/ControlUnit/U42  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n13 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n12 ), .A3(
        \dp/id_stage/regfile/ControlUnit/current_state[3] ), .ZN(
        \dp/id_stage/regfile/cnt_swp ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U41  ( .A1(1'b0), .A2(
        \dp/id_stage/regfile/ControlUnit/n5 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n19 ) );
  AOI21_X1 \dp/id_stage/regfile/ControlUnit/U40  ( .B1(
        \dp/id_stage/regfile/ControlUnit/n17 ), .B2(
        \dp/id_stage/regfile/ControlUnit/n19 ), .A(RST), .ZN(
        \dp/id_stage/regfile/ControlUnit/next_state [1]) );
  AOI21_X1 \dp/id_stage/regfile/ControlUnit/U39  ( .B1(
        \dp/id_stage/regfile/ControlUnit/n17 ), .B2(
        \dp/id_stage/regfile/ControlUnit/n18 ), .A(RST), .ZN(
        \dp/id_stage/regfile/ControlUnit/next_state [2]) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U38  ( .A(
        \dp/id_stage/regfile/ControlUnit/n26 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n11 ) );
  AOI21_X1 \dp/id_stage/regfile/ControlUnit/U37  ( .B1(
        \dp/id_stage/regfile/ControlUnit/n5 ), .B2(
        \dp/id_stage/regfile/ControlUnit/n23 ), .A(\dp/id_stage/regfile/rd_cu ), .ZN(\dp/id_stage/regfile/ControlUnit/n22 ) );
  AOI22_X1 \dp/id_stage/regfile/ControlUnit/U36  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n11 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n12 ), .B1(
        \dp/id_stage/regfile/ControlUnit/n25 ), .B2(
        \dp/id_stage/regfile/ControlUnit/n14 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n21 ) );
  AOI21_X1 \dp/id_stage/regfile/ControlUnit/U35  ( .B1(
        \dp/id_stage/regfile/ControlUnit/n21 ), .B2(
        \dp/id_stage/regfile/ControlUnit/n22 ), .A(RST), .ZN(
        \dp/id_stage/regfile/ControlUnit/next_state [0]) );
  NOR3_X1 \dp/id_stage/regfile/ControlUnit/U34  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n16 ), .A2(RST), .A3(
        \dp/id_stage/regfile/ControlUnit/n8 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/next_state [3]) );
  AOI21_X1 \dp/id_stage/regfile/ControlUnit/U33  ( .B1(
        \dp/id_stage/regfile/ControlUnit/n13 ), .B2(
        \dp/id_stage/regfile/ControlUnit/current_state[3] ), .A(
        \dp/id_stage/regfile/ControlUnit/n27 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n26 ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U32  ( .A(
        \dp/id_stage/regfile/ControlUnit/n29 ), .ZN(
        \dp/id_stage/regfile/wr_cu ) );
  NOR2_X1 \dp/id_stage/regfile/ControlUnit/U31  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n14 ), .A2(
        \dp/id_stage/regfile/ControlUnit/current_state[2] ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n40 ) );
  NOR2_X1 \dp/id_stage/regfile/ControlUnit/U30  ( .A1(
        \dp/id_stage/regfile/ControlUnit/current_state[3] ), .A2(
        \dp/id_stage/regfile/ControlUnit/current_state[1] ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n25 ) );
  NOR2_X1 \dp/id_stage/regfile/ControlUnit/U29  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n13 ), .A2(
        \dp/id_stage/regfile/ControlUnit/current_state[3] ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n27 ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U28  ( .A(
        \dp/id_stage/regfile/up_dwn_cwp ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n4 ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U27  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n35 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n4 ), .ZN(
        \dp/id_stage/regfile/up_dwn_rest ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U26  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n35 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n29 ), .ZN(rf_fill_i) );
  AND3_X1 \dp/id_stage/regfile/ControlUnit/U25  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n38 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n32 ), .A3(
        \dp/id_stage/regfile/ControlUnit/n39 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n34 ) );
  NAND4_X1 \dp/id_stage/regfile/ControlUnit/U24  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n30 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n31 ), .A3(
        \dp/id_stage/regfile/ControlUnit/n32 ), .A4(
        \dp/id_stage/regfile/ControlUnit/n8 ), .ZN(
        \dp/id_stage/regfile/up_dwn_swp ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U23  ( .A(
        \dp/id_stage/regfile/ControlUnit/n28 ), .ZN(
        \dp/id_stage/regfile/rd_cu ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U22  ( .A(
        \dp/id_stage/regfile/ControlUnit/n32 ), .ZN(
        \dp/id_stage/regfile/rst_rf ) );
  NOR2_X1 \dp/id_stage/regfile/ControlUnit/U21  ( .A1(
        \dp/id_stage/regfile/cnt_swp ), .A2(\dp/id_stage/regfile/rf_enable ), 
        .ZN(\dp/id_stage/regfile/ControlUnit/n39 ) );
  AOI21_X1 \dp/id_stage/regfile/ControlUnit/U20  ( .B1(
        \dp/id_stage/regfile/ControlUnit/n16 ), .B2(
        \dp/id_stage/regfile/rf_enable ), .A(
        \dp/id_stage/regfile/ControlUnit/n20 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n17 ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U19  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n37 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n28 ), .ZN(rf_spill_i) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U18  ( .A(rf_spill_i), .ZN(
        \dp/id_stage/regfile/ControlUnit/n3 ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U17  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n30 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n3 ), .ZN(
        \dp/id_stage/regfile/sel_wp ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U16  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n40 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n25 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n38 ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U15  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n36 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n33 ), .ZN(
        \dp/id_stage/regfile/cnt_save ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U14  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n37 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n35 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n20 ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U13  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n40 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n27 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n37 ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U12  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n29 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n28 ), .ZN(
        \dp/id_stage/regfile/rf_enable ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U11  ( .A(
        \dp/id_stage/regfile/rf_enable ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n8 ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U10  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n39 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n31 ), .ZN(
        \dp/id_stage/regfile/rst_swp ) );
  NAND4_X1 \dp/id_stage/regfile/ControlUnit/U9  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n39 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n37 ), .A3(
        \dp/id_stage/regfile/ControlUnit/n38 ), .A4(
        \dp/id_stage/regfile/ControlUnit/n9 ), .ZN(
        \dp/id_stage/regfile/rst_spill_fill ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U8  ( .A(
        \dp/id_stage/regfile/ControlUnit/n20 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n2 ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U7  ( .A(
        \dp/id_stage/regfile/cnt_save ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n9 ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U6  ( .A(
        \dp/id_stage/regfile/ControlUnit/n38 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n5 ) );
  NAND2_X1 \dp/id_stage/regfile/ControlUnit/U5  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n2 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n9 ), .ZN(
        \dp/id_stage/regfile/cnt_cwp ) );
  NOR2_X1 \dp/id_stage/regfile/ControlUnit/U4  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n5 ), .A2(
        \dp/id_stage/regfile/cnt_cwp ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n31 ) );
  INV_X1 \dp/id_stage/regfile/ControlUnit/U3  ( .A(
        \dp/id_stage/regfile/ControlUnit/n31 ), .ZN(
        \dp/id_stage/regfile/cpu_work ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U56  ( .A1(
        \dp/id_stage/regfile/ControlUnit/current_state[2] ), .A2(
        \dp/id_stage/regfile/ControlUnit/current_state[0] ), .A3(
        \dp/id_stage/regfile/ControlUnit/n25 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n35 ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U55  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n14 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n12 ), .A3(
        \dp/id_stage/regfile/ControlUnit/n27 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n36 ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U54  ( .A1(
        \dp/id_stage/regfile/ControlUnit/current_state[2] ), .A2(
        \dp/id_stage/regfile/ControlUnit/n14 ), .A3(
        \dp/id_stage/regfile/ControlUnit/n25 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n33 ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U53  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n27 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n14 ), .A3(
        \dp/id_stage/regfile/ControlUnit/current_state[2] ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n29 ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U52  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n14 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n12 ), .A3(
        \dp/id_stage/regfile/ControlUnit/n25 ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n32 ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U51  ( .A1(
        \dp/id_stage/regfile/ControlUnit/current_state[0] ), .A2(
        \dp/id_stage/regfile/ControlUnit/n27 ), .A3(
        \dp/id_stage/regfile/ControlUnit/current_state[2] ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n28 ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U50  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n40 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n13 ), .A3(
        \dp/id_stage/regfile/ControlUnit/current_state[3] ), .ZN(
        \dp/id_stage/regfile/ControlUnit/n30 ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U49  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n36 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n37 ), .A3(
        \dp/id_stage/regfile/ControlUnit/n34 ), .ZN(
        \dp/id_stage/regfile/up_dwn_cwp ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U48  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n2 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n33 ), .A3(
        \dp/id_stage/regfile/ControlUnit/n34 ), .ZN(
        \dp/id_stage/regfile/up_dwn_save ) );
  NAND3_X1 \dp/id_stage/regfile/ControlUnit/U47  ( .A1(
        \dp/id_stage/regfile/ControlUnit/n5 ), .A2(
        \dp/id_stage/regfile/ControlUnit/n15 ), .A3(1'b0), .ZN(
        \dp/id_stage/regfile/ControlUnit/n18 ) );
  DFF_X1 \dp/id_stage/regfile/ControlUnit/current_state_reg[3]  ( .D(
        \dp/id_stage/regfile/ControlUnit/next_state [3]), .CK(CLK), .Q(
        \dp/id_stage/regfile/ControlUnit/current_state[3] ) );
  DFF_X1 \dp/id_stage/regfile/ControlUnit/current_state_reg[2]  ( .D(
        \dp/id_stage/regfile/ControlUnit/next_state [2]), .CK(CLK), .Q(
        \dp/id_stage/regfile/ControlUnit/current_state[2] ), .QN(
        \dp/id_stage/regfile/ControlUnit/n12 ) );
  DFF_X1 \dp/id_stage/regfile/ControlUnit/current_state_reg[1]  ( .D(
        \dp/id_stage/regfile/ControlUnit/next_state [1]), .CK(CLK), .Q(
        \dp/id_stage/regfile/ControlUnit/current_state[1] ), .QN(
        \dp/id_stage/regfile/ControlUnit/n13 ) );
  DFF_X1 \dp/id_stage/regfile/ControlUnit/current_state_reg[0]  ( .D(
        \dp/id_stage/regfile/ControlUnit/next_state [0]), .CK(CLK), .Q(
        \dp/id_stage/regfile/ControlUnit/current_state[0] ), .QN(
        \dp/id_stage/regfile/ControlUnit/n14 ) );
  AND3_X1 \dp/id_stage/regfile/DataPath/U4  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_sf_in[1] ), .A2(
        \dp/id_stage/regfile/DataPath/addr_sf_in[0] ), .A3(
        \dp/id_stage/regfile/DataPath/addr_sf_in[2] ), .ZN(
        \dp/id_stage/regfile/end_sf ) );
  INV_X1 \dp/id_stage/regfile/DataPath/U3  ( .A(
        \dp/id_stage/regfile/DataPath/CWP[0] ), .ZN(
        \dp/id_stage/regfile/DataPath/cwp_1[0] ) );
  AOI21_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U20  ( .B1(
        \dp/id_stage/p_addr_wRS1 [3]), .B2(\dp/id_stage/p_addr_wRS1 [2]), .A(
        \dp/id_stage/p_addr_wRS1 [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/N1 ) );
  XNOR2_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U19  ( .A(
        \dp/id_stage/p_addr_wRS1 [3]), .B(
        \dp/id_stage/regfile/DataPath/CWP[0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n18 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U18  ( .A(
        \dp/id_stage/p_addr_wRS1 [3]), .B(\dp/id_stage/p_addr_wRS1 [2]), .Z(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n4 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U17  ( .A1(
        \dp/id_stage/p_addr_wRS1 [3]), .A2(\dp/id_stage/p_addr_wRS1 [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n3 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U16  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_RD1/N5 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ), .B1(
        \dp/id_stage/p_addr_wRS1 [2]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n20 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U15  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n20 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [2]) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U14  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n1 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [4]) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U13  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n4 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n19 ) );
  OAI21_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U12  ( .B1(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n18 ), .B2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ), .A(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n19 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [3]) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U11  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n2 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [5]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U10  ( .A1(
        \dp/id_stage/p_addr_wRS1 [1]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ), .B1(
        \dp/id_stage/p_addr_wRS1 [1]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n21 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U9  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n21 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [1]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U8  ( .A1(
        \dp/id_stage/p_addr_wRS1 [0]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ), .B1(
        \dp/id_stage/p_addr_wRS1 [0]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n22 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U7  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n22 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [0]) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U6  ( .A(
        \dp/id_stage/p_addr_wRS1 [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/N5 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U5  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_RD1/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n8 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U4  ( .A1(
        \dp/id_stage/p_addr_wRS1 [4]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n3 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n2 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Conv_RD1/U3  ( .A(
        \dp/id_stage/p_addr_wRS1 [4]), .B(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n3 ), .Z(
        \dp/id_stage/regfile/DataPath/Conv_RD1/n1 ) );
  AOI21_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U20  ( .B1(
        \dp/id_stage/p_addr_wRS2 [3]), .B2(\dp/id_stage/p_addr_wRS2 [2]), .A(
        \dp/id_stage/p_addr_wRS2 [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/N1 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U19  ( .A1(
        \dp/id_stage/p_addr_wRS2 [1]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ), .B1(
        \dp/id_stage/p_addr_wRS2 [1]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n10 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U18  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n10 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [1]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U17  ( .A1(
        \dp/id_stage/p_addr_wRS2 [0]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ), .B1(
        \dp/id_stage/p_addr_wRS2 [0]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n9 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U16  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n9 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [0]) );
  XNOR2_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U15  ( .A(
        \dp/id_stage/p_addr_wRS2 [3]), .B(
        \dp/id_stage/regfile/DataPath/CWP[0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n13 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U14  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n1 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n12 ) );
  OAI21_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U13  ( .B1(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n13 ), .B2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ), .A(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n12 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [3]) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U12  ( .A1(
        \dp/id_stage/p_addr_wRS2 [3]), .A2(\dp/id_stage/p_addr_wRS2 [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n4 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U11  ( .A1(
        \dp/id_stage/p_addr_wRS2 [4]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n3 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U10  ( .A(
        \dp/id_stage/p_addr_wRS2 [4]), .B(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n4 ), .Z(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n2 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U9  ( .A(
        \dp/id_stage/p_addr_wRS2 [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/N5 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U8  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_RD2/N5 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ), .B1(
        \dp/id_stage/p_addr_wRS2 [2]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n11 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U7  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n11 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [2]) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U6  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_RD2/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U5  ( .A(
        \dp/id_stage/p_addr_wRS2 [3]), .B(\dp/id_stage/p_addr_wRS2 [2]), .Z(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n1 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U4  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n3 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [5]) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_RD2/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n2 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_RD2/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [4]) );
  AOI21_X1 \dp/id_stage/regfile/DataPath/Conv_W/U20  ( .B1(
        \dp/id_stage/p_addr_wRD [3]), .B2(\dp/id_stage/p_addr_wRD [2]), .A(
        \dp/id_stage/p_addr_wRD [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/N1 ) );
  XNOR2_X1 \dp/id_stage/regfile/DataPath/Conv_W/U19  ( .A(
        \dp/id_stage/p_addr_wRD [3]), .B(\dp/id_stage/regfile/DataPath/CWP[0] ), .ZN(\dp/id_stage/regfile/DataPath/Conv_W/n13 ) );
  OAI21_X1 \dp/id_stage/regfile/DataPath/Conv_W/U18  ( .B1(
        \dp/id_stage/regfile/DataPath/Conv_W/n13 ), .B2(
        \dp/id_stage/regfile/DataPath/Conv_W/n8 ), .A(
        \dp/id_stage/regfile/DataPath/Conv_W/n12 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_w_p [3]) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Conv_W/U17  ( .A(
        \dp/id_stage/p_addr_wRD [3]), .B(\dp/id_stage/p_addr_wRD [2]), .Z(
        \dp/id_stage/regfile/DataPath/Conv_W/n4 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_W/U16  ( .A1(
        \dp/id_stage/p_addr_wRD [3]), .A2(\dp/id_stage/p_addr_wRD [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/n3 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_W/U15  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_W/n1 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_W/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_w_p [4]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_W/U14  ( .A1(
        \dp/id_stage/p_addr_wRD [1]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_W/n8 ), .B1(
        \dp/id_stage/p_addr_wRD [1]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_W/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/n10 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_W/U13  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_W/n10 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_w_p [1]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_W/U12  ( .A1(
        \dp/id_stage/p_addr_wRD [0]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_W/n8 ), .B1(
        \dp/id_stage/p_addr_wRD [0]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_W/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/n9 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_W/U11  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_W/n9 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_w_p [0]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Conv_W/U10  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_W/N5 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_W/n8 ), .B1(
        \dp/id_stage/p_addr_wRD [2]), .B2(
        \dp/id_stage/regfile/DataPath/Conv_W/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/n11 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_W/U9  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_W/n11 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_w_p [2]) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_W/U8  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_W/n2 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_W/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/addr_w_p [5]) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_W/U7  ( .A(
        \dp/id_stage/p_addr_wRD [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/N5 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Conv_W/U6  ( .A(
        \dp/id_stage/regfile/DataPath/Conv_W/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/n8 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Conv_W/U5  ( .A1(
        \dp/id_stage/p_addr_wRD [4]), .A2(
        \dp/id_stage/regfile/DataPath/Conv_W/n3 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/n2 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Conv_W/U4  ( .A(
        \dp/id_stage/p_addr_wRD [4]), .B(
        \dp/id_stage/regfile/DataPath/Conv_W/n3 ), .Z(
        \dp/id_stage/regfile/DataPath/Conv_W/n1 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Conv_W/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/Conv_W/n4 ), .A2(
        \dp/id_stage/regfile/DataPath/Conv_W/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/Conv_W/n12 ) );
  AOI21_X1 \dp/id_stage/regfile/DataPath/SF_converter/U20  ( .B1(1'b0), .B2(
        \dp/id_stage/regfile/DataPath/addr_sf_in[2] ), .A(1'b0), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/N1 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/SF_converter/U19  ( .A1(1'b0), .A2(
        \dp/id_stage/regfile/DataPath/SF_converter/n2 ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/n4 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/SF_converter/U18  ( .A(1'b0), .B(
        \dp/id_stage/regfile/DataPath/SF_converter/n2 ), .Z(
        \dp/id_stage/regfile/DataPath/SF_converter/n3 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/SF_converter/U17  ( .A1(1'b0), .A2(
        \dp/id_stage/regfile/DataPath/addr_sf_in[2] ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/n2 ) );
  XNOR2_X1 \dp/id_stage/regfile/DataPath/SF_converter/U16  ( .A(1'b0), .B(
        \dp/id_stage/regfile/DataPath/sf_wp[0] ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/n9 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/SF_converter/U15  ( .A1(
        \dp/id_stage/regfile/DataPath/SF_converter/n1 ), .A2(
        \dp/id_stage/regfile/DataPath/SF_converter/n10 ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/n8 ) );
  OAI21_X1 \dp/id_stage/regfile/DataPath/SF_converter/U14  ( .B1(
        \dp/id_stage/regfile/DataPath/SF_converter/n9 ), .B2(
        \dp/id_stage/regfile/DataPath/SF_converter/n10 ), .A(
        \dp/id_stage/regfile/DataPath/SF_converter/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[3] ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/SF_converter/U13  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_sf_in[1] ), .A2(
        \dp/id_stage/regfile/DataPath/SF_converter/n10 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_sf_in[1] ), .B2(
        \dp/id_stage/regfile/DataPath/SF_converter/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/n6 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/SF_converter/U12  ( .A(
        \dp/id_stage/regfile/DataPath/SF_converter/n6 ), .ZN(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[1] ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/SF_converter/U11  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_sf_in[0] ), .A2(
        \dp/id_stage/regfile/DataPath/SF_converter/n10 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_sf_in[0] ), .B2(
        \dp/id_stage/regfile/DataPath/SF_converter/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/n5 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/SF_converter/U10  ( .A(
        \dp/id_stage/regfile/DataPath/SF_converter/n5 ), .ZN(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[0] ) );
  INV_X1 \dp/id_stage/regfile/DataPath/SF_converter/U9  ( .A(
        \dp/id_stage/regfile/DataPath/addr_sf_in[2] ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/N5 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/SF_converter/U8  ( .A1(
        \dp/id_stage/regfile/DataPath/SF_converter/N5 ), .A2(
        \dp/id_stage/regfile/DataPath/SF_converter/n10 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_sf_in[2] ), .B2(
        \dp/id_stage/regfile/DataPath/SF_converter/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/n7 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/SF_converter/U7  ( .A(
        \dp/id_stage/regfile/DataPath/SF_converter/n7 ), .ZN(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[2] ) );
  INV_X1 \dp/id_stage/regfile/DataPath/SF_converter/U6  ( .A(
        \dp/id_stage/regfile/DataPath/SF_converter/N1 ), .ZN(
        \dp/id_stage/regfile/DataPath/SF_converter/n10 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/SF_converter/U5  ( .A(1'b0), .B(
        \dp/id_stage/regfile/DataPath/addr_sf_in[2] ), .Z(
        \dp/id_stage/regfile/DataPath/SF_converter/n1 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/SF_converter/U4  ( .A1(
        \dp/id_stage/regfile/DataPath/SF_converter/n3 ), .A2(
        \dp/id_stage/regfile/DataPath/SF_converter/n10 ), .ZN(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[4] ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/SF_converter/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/SF_converter/n4 ), .A2(
        \dp/id_stage/regfile/DataPath/SF_converter/n10 ), .ZN(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[5] ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Cwp_counter/U6  ( .A(1'b0), .ZN(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n2 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Cwp_counter/U5  ( .A(
        \dp/id_stage/regfile/rst_swp ), .ZN(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n4 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Cwp_counter/U4  ( .A1(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n3 ), .A2(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n2 ), .B1(1'b0), .B2(1'b0), 
        .ZN(\dp/id_stage/regfile/DataPath/Cwp_counter/n1 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Cwp_counter/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n1 ), .A2(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n5 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Cwp_counter/U7  ( .A(
        \dp/id_stage/regfile/cnt_cwp ), .B(
        \dp/id_stage/regfile/DataPath/CWP[0] ), .Z(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n3 ) );
  DFF_X1 \dp/id_stage/regfile/DataPath/Cwp_counter/Q_reg[0]  ( .D(
        \dp/id_stage/regfile/DataPath/Cwp_counter/n5 ), .CK(CLK), .Q(
        \dp/id_stage/regfile/DataPath/CWP[0] ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Swp_counter/U6  ( .A(1'b0), .ZN(
        \dp/id_stage/regfile/DataPath/Swp_counter/n2 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Swp_counter/U5  ( .A(
        \dp/id_stage/regfile/rst_swp ), .ZN(
        \dp/id_stage/regfile/DataPath/Swp_counter/n4 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Swp_counter/U4  ( .A1(
        \dp/id_stage/regfile/DataPath/Swp_counter/n7 ), .A2(
        \dp/id_stage/regfile/DataPath/Swp_counter/n2 ), .B1(1'b0), .B2(1'b0), 
        .ZN(\dp/id_stage/regfile/DataPath/Swp_counter/n8 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Swp_counter/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/Swp_counter/n8 ), .A2(
        \dp/id_stage/regfile/DataPath/Swp_counter/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/Swp_counter/n6 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Swp_counter/U7  ( .A(
        \dp/id_stage/regfile/cnt_swp ), .B(
        \dp/id_stage/regfile/DataPath/Swp_counter/Q[0] ), .Z(
        \dp/id_stage/regfile/DataPath/Swp_counter/n7 ) );
  DFF_X1 \dp/id_stage/regfile/DataPath/Swp_counter/Q_reg[0]  ( .D(
        \dp/id_stage/regfile/DataPath/Swp_counter/n6 ), .CK(CLK), .Q(
        \dp/id_stage/regfile/DataPath/Swp_counter/Q[0] ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U18  ( .A(1'b0), 
        .ZN(\dp/id_stage/regfile/DataPath/Spill_fill_counter/n4 ) );
  XNOR2_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U17  ( .A(1'b1), 
        .B(\dp/id_stage/regfile/DataPath/Spill_fill_counter/n11 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n10 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U16  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_sf_in[1] ), .A2(
        \dp/id_stage/regfile/DataPath/addr_sf_in[0] ), .B1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n11 ), .B2(1'b1), 
        .ZN(\dp/id_stage/regfile/DataPath/Spill_fill_counter/n9 ) );
  XNOR2_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U15  ( .A(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n9 ), .B(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n10 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n7 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U14  ( .A1(1'b0), 
        .A2(1'b0), .B1(\dp/id_stage/regfile/DataPath/Spill_fill_counter/n1 ), 
        .B2(\dp/id_stage/regfile/DataPath/Spill_fill_counter/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n18 ) );
  OR2_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U13  ( .A1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n14 ), .A2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n18 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n17 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U12  ( .A1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n1 ), .A2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n12 ), .B1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n16 ), .B2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n17 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n21 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U11  ( .A1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n10 ), .A2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n4 ), .B1(1'b0), .B2(
        1'b0), .ZN(\dp/id_stage/regfile/DataPath/Spill_fill_counter/n15 ) );
  OR2_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U10  ( .A1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n14 ), .A2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n15 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n13 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U9  ( .A1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n3 ), .A2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n12 ), .B1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n16 ), .B2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n13 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n20 ) );
  OAI21_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U8  ( .B1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n7 ), .B2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n2 ), .A(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n6 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U7  ( .A1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n6 ), .A2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n4 ), .B1(1'b0), .B2(
        1'b0), .ZN(\dp/id_stage/regfile/DataPath/Spill_fill_counter/n5 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U6  ( .A1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n2 ), .A2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n12 ), .B1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n5 ), .B2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n16 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n19 ) );
  NOR3_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U5  ( .A1(
        \dp/id_stage/regfile/rf_enable ), .A2(1'b0), .A3(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n16 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n14 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U4  ( .A(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n14 ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n12 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U3  ( .A(
        \dp/id_stage/regfile/rst_spill_fill ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n16 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U23  ( .A(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n3 ), .B(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n1 ), .Z(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n11 ) );
  NAND3_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/U22  ( .A1(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n7 ), .A2(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n2 ), .A3(
        \dp/id_stage/regfile/rf_enable ), .ZN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n8 ) );
  DFF_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/Q_reg[2]  ( .D(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n19 ), .CK(CLK), .Q(
        \dp/id_stage/regfile/DataPath/addr_sf_in[2] ), .QN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n2 ) );
  DFF_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/Q_reg[1]  ( .D(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n20 ), .CK(CLK), .Q(
        \dp/id_stage/regfile/DataPath/addr_sf_in[1] ), .QN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n3 ) );
  DFF_X1 \dp/id_stage/regfile/DataPath/Spill_fill_counter/Q_reg[0]  ( .D(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n21 ), .CK(CLK), .Q(
        \dp/id_stage/regfile/DataPath/addr_sf_in[0] ), .QN(
        \dp/id_stage/regfile/DataPath/Spill_fill_counter/n1 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/CANSAVE_counter/U6  ( .A(
        \dp/id_stage/regfile/rst_rf ), .ZN(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n4 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/CANSAVE_counter/U5  ( .A1(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n7 ), .A2(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n4 ), .B1(
        \dp/id_stage/regfile/rst_rf ), .B2(1'b0), .ZN(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n8 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/CANSAVE_counter/U4  ( .A(1'b1), .ZN(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n2 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/CANSAVE_counter/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n8 ), .A2(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n2 ), .ZN(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n6 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/CANSAVE_counter/U7  ( .A(
        \dp/id_stage/regfile/cnt_save ), .B(\dp/id_stage/regfile/cansave ), 
        .Z(\dp/id_stage/regfile/DataPath/CANSAVE_counter/n7 ) );
  DFF_X1 \dp/id_stage/regfile/DataPath/CANSAVE_counter/Q_reg[0]  ( .D(
        \dp/id_stage/regfile/DataPath/CANSAVE_counter/n6 ), .CK(CLK), .Q(
        \dp/id_stage/regfile/cansave ) );
  INV_X1 \dp/id_stage/regfile/DataPath/CANRESTORE_counter/U6  ( .A(1'b0), .ZN(
        \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n2 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/CANRESTORE_counter/U5  ( .A(
        \dp/id_stage/regfile/rst_swp ), .ZN(
        \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n4 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/CANRESTORE_counter/U4  ( .A1(
        \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n7 ), .A2(
        \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n2 ), .B1(1'b0), .B2(
        1'b0), .ZN(\dp/id_stage/regfile/DataPath/CANRESTORE_counter/n8 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/CANRESTORE_counter/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n8 ), .A2(
        \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n6 ) );
  XOR2_X1 \dp/id_stage/regfile/DataPath/CANRESTORE_counter/U7  ( .A(
        \dp/id_stage/regfile/cnt_save ), .B(\dp/id_stage/regfile/canrestore ), 
        .Z(\dp/id_stage/regfile/DataPath/CANRESTORE_counter/n7 ) );
  DFF_X1 \dp/id_stage/regfile/DataPath/CANRESTORE_counter/Q_reg[0]  ( .D(
        \dp/id_stage/regfile/DataPath/CANRESTORE_counter/n6 ), .CK(CLK), .Q(
        \dp/id_stage/regfile/canrestore ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U13  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[2] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_rd/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [2]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd/n11 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U12  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_rd/n11 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_rd_out [2]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U11  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[4] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_rd/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [4]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd/n9 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U10  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_rd/n9 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_rd_out [4]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U9  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[3] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_rd/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [3]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd/n10 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U8  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_rd/n10 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_rd_out [3]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U7  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[5] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_rd/n1 ), .B1(
        \dp/id_stage/regfile/cpu_work ), .B2(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd/n8 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U6  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_rd/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_rd_out [5]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U5  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[1] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_rd/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [1]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd/n12 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U4  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_rd/n12 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_rd_out [1]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[0] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_rd/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_rd1_p [0]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd/n13 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U2  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_rd/n13 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_rd_out [0]) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd/U1  ( .A(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd/n1 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U13  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[3] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_wr/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_w_p [3]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr/n5 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U12  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_wr/n5 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_wr_out [3]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U11  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[4] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_wr/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_w_p [4]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr/n6 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U10  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_wr/n6 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_wr_out [4]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U9  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[1] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_wr/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_w_p [1]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr/n3 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U8  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_wr/n3 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_wr_out [1]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U7  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[0] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_wr/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_w_p [0]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr/n2 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U6  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_wr/n2 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_wr_out [0]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U5  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[2] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_wr/n1 ), .B1(
        \dp/id_stage/regfile/DataPath/addr_w_p [2]), .B2(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr/n4 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U4  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_wr/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/spill_fill_addr[5] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_wr/n1 ), .B1(
        \dp/id_stage/regfile/cpu_work ), .B2(
        \dp/id_stage/regfile/DataPath/addr_w_p [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr/n7 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U2  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_wr/n7 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_wr_out [5]) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr/U1  ( .A(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr/n1 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_sf/U3  ( .A(
        \dp/id_stage/regfile/sel_wp ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_sf/n1 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_sf/U2  ( .A1(
        \dp/id_stage/regfile/DataPath/CWP[0] ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_sf/n1 ), .B1(
        \dp/id_stage/regfile/sel_wp ), .B2(
        \dp/id_stage/regfile/DataPath/cwp_1[0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_sf/n3 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_sf/U1  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_sf/n3 ), .ZN(
        \dp/id_stage/regfile/DataPath/sf_wp[0] ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd1_control/U3  ( .A(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd1_control/n2 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_rd1_control/U2  ( .A1(
        \dp/id_stage/regfile/rd_cu ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_rd1_control/n2 ), .B1(
        \dp/id_stage/regfile/cpu_work ), .B2(rf_rs1_en_i), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd1_control/n3 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd1_control/U1  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_rd1_control/n3 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_rd1_control_out ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd2_control/U3  ( .A(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd2_control/n2 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_rd2_control/U2  ( .A1(1'b0), .A2(
        \dp/id_stage/regfile/DataPath/Mux_rd2_control/n2 ), .B1(
        \dp/id_stage/regfile/cpu_work ), .B2(rf_rs2_en_i), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_rd2_control/n4 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_rd2_control/U1  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_rd2_control/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_rd2_control_out ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_wr_control/U3  ( .A1(
        \dp/id_stage/regfile/wr_cu ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_wr_control/n2 ), .B1(
        \dp/id_stage/regfile/cpu_work ), .B2(rf_we_i), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr_control/n4 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr_control/U2  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_wr_control/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_wr_control_out ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_wr_control/U1  ( .A(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_wr_control/n2 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_en_control/U3  ( .A(
        \dp/id_stage/regfile/cpu_work ), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_en_control/n2 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Mux_en_control/U2  ( .A1(
        \dp/id_stage/regfile/rf_enable ), .A2(
        \dp/id_stage/regfile/DataPath/Mux_en_control/n2 ), .B1(
        \dp/id_stage/regfile/cpu_work ), .B2(1'b1), .ZN(
        \dp/id_stage/regfile/DataPath/Mux_en_control/n4 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Mux_en_control/U1  ( .A(
        \dp/id_stage/regfile/DataPath/Mux_en_control/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/mux_en_control_out ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3831  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/N428 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4239 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3830  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/N428 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3829  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/N428 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3828  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/N428 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3827  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/N429 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4235 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3826  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/N429 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3825  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/N429 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3824  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/N429 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3823  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1346 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3822  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1346 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3821  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1346 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3820  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1346 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3819  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1346 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3818  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1346 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3817  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1348 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3816  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1348 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3815  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1348 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3814  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1348 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3813  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1348 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3812  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1348 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3811  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1516 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1226 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3810  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1516 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3809  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1516 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3808  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1516 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3807  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1518 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3806  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1518 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3805  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1518 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1220 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3804  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1585 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3803  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1585 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3802  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1585 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3801  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1585 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3800  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1586 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3799  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1586 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3798  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1687 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1213 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3797  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1687 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3796  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1688 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3795  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1688 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3794  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1688 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3793  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1688 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3792  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1688 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1207 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3791  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1755 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3790  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1755 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3789  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1756 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3788  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1756 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3787  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1756 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3786  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1756 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3785  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1857 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1189 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3784  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1857 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3783  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1857 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3782  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1857 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3781  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1857 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3780  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1857 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3779  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1858 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3778  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1858 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3777  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1858 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3776  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1858 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3775  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1858 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3774  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1858 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ) );
  CLKBUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3773  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1925 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1177 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3772  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_rd2_control_out ), .A2(
        \dp/id_stage/regfile/DataPath/mux_en_control_out ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N429 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3771  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_rd1_control_out ), .A2(
        \dp/id_stage/regfile/DataPath/mux_en_control_out ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N428 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3770  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n450 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n418 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2553 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2541 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3769  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2523 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2524 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2525 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2526 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2522 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3768  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2541 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2542 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2543 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2544 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2521 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3767  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2521 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2522 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N396 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3766  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n450 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n418 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3180 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3168 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3765  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3150 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3151 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3152 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3153 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3149 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3764  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3168 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3169 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3170 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3171 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3148 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3763  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3148 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3149 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N328 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3762  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n451 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n419 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2520 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2513 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3761  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2505 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2506 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2507 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2508 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2504 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3760  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2513 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2514 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2515 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2516 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2503 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3759  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2503 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2504 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N397 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3758  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n451 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n419 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3147 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3140 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3757  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3132 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3133 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3134 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3135 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3131 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3756  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3140 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3141 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3142 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3143 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3130 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3755  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3130 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3131 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N329 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3754  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n452 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n420 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2502 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2495 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3753  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2487 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2488 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2489 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2490 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2486 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3752  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2495 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2496 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2497 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2498 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2485 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3751  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2485 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2486 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N398 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3750  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n452 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n420 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3129 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3122 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3749  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3114 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3115 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3116 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3117 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3113 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3748  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3122 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3123 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3124 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3125 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3112 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3747  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3112 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3113 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N330 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3746  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n453 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n421 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2484 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2477 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3745  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2469 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2470 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2471 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2472 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2468 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3744  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2477 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2478 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2479 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2480 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2467 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3743  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2467 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2468 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N399 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3742  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n453 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n421 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3111 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3104 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3741  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3096 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3097 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3098 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3099 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3095 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3740  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3104 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3105 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3106 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3107 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3094 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3739  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3094 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3095 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N331 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3738  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n454 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n422 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2466 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2459 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3737  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2451 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2452 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2453 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2454 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2450 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3736  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2459 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2460 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2461 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2462 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2449 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3735  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2449 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2450 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N400 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3734  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n454 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n422 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3093 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3086 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3733  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3078 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3079 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3080 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3081 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3077 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3732  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3086 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3087 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3088 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3089 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3076 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3731  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3076 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3077 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N332 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3730  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n455 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n423 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2448 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2441 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3729  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2433 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2434 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2435 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2436 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2432 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3728  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2441 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2442 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2443 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2444 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2431 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3727  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2431 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2432 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N401 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3726  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n455 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n423 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3075 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3068 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3725  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3060 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3061 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3062 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3063 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3059 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3724  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3068 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3069 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3070 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3071 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3058 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3723  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3058 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3059 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N333 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3722  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n456 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n424 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2430 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2423 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3721  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2415 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2416 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2417 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2418 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2414 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3720  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2423 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2424 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2425 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2426 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2413 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3719  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2413 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2414 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N402 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3718  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n456 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n424 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3057 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3050 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3717  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3042 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3043 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3044 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3045 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3041 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3716  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3050 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3051 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3052 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3053 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3040 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3715  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3040 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3041 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N334 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3714  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n457 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n425 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2412 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2405 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3713  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2397 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2398 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2399 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2400 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2396 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3712  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2405 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2406 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2407 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2408 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2395 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3711  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2395 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2396 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N403 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3710  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n457 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n425 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3039 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3032 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3709  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3024 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3025 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3026 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3027 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3023 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3708  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3032 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3033 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3034 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3035 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3022 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3707  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3022 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3023 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N335 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3706  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n458 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n426 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2394 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2387 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3705  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2379 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2380 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2381 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2382 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2378 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3704  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2387 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2388 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2389 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2390 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2377 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3703  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2377 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2378 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N404 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3702  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n458 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n426 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3021 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3014 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3701  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3006 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3007 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3008 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3009 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3005 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3700  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3014 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3015 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3016 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3017 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3004 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3699  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3004 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3005 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N336 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3698  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n459 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n427 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2376 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2369 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3697  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2361 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2362 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2363 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2364 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2360 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3696  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2369 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2370 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2371 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2372 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2359 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3695  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2359 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2360 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N405 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3694  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n459 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n427 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3003 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2996 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3693  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2988 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2989 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2990 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2991 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2987 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3692  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2996 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2997 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2998 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2999 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2986 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3691  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2986 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2987 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N337 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3690  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n460 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n428 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2358 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2351 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3689  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2343 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2344 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2345 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2346 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2342 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3688  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2351 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2352 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2353 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2354 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2341 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3687  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2341 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2342 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N406 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3686  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n460 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n428 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2985 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2978 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3685  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2970 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2971 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2972 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2973 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2969 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3684  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2978 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2979 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2980 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2981 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2968 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3683  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2968 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2969 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N338 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3682  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n461 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n429 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2340 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2333 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3681  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2325 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2326 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2327 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2328 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2324 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3680  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2333 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2334 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2335 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2336 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2323 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3679  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2323 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2324 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N407 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3678  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n461 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n429 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2967 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2960 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3677  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2952 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2953 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2954 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2955 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2951 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3676  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2960 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2961 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2962 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2963 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2950 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3675  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2950 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2951 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N339 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3674  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n462 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n430 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2322 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2315 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3673  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2307 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2308 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2309 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2310 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2306 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3672  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2315 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2316 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2317 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2318 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2305 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3671  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2305 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2306 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N408 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3670  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n462 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n430 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2949 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2942 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3669  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2934 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2935 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2936 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2937 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2933 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3668  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2942 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2943 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2944 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2945 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2932 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3667  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2932 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2933 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N340 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3666  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n463 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n431 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2304 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2297 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3665  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2289 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2290 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2291 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2292 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2288 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3664  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2297 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2298 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2299 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2300 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2287 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3663  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2287 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2288 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N409 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3662  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n463 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n431 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2931 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2924 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3661  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2916 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2917 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2918 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2919 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2915 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3660  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2924 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2925 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2926 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2927 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2914 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3659  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2914 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2915 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N341 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3658  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n464 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n432 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2286 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2279 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3657  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2272 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2273 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2274 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2270 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3656  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2279 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2280 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2281 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2282 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2269 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3655  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2270 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N410 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3654  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n464 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n432 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2913 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2906 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3653  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2898 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2899 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2900 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2901 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2897 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3652  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2906 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2907 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2908 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2909 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2896 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3651  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2896 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2897 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N342 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3650  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n465 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n433 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2268 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2261 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3649  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2254 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2255 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2256 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2252 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3648  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2262 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2263 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2264 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2251 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3647  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2252 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N411 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3646  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n465 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n433 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2895 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2888 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3645  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2880 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2881 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2882 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2883 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2879 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3644  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2889 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2890 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2891 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2878 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3643  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2878 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2879 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N343 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3642  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n466 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n434 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2250 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2243 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3641  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2235 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2236 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2237 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2238 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2234 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3640  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2243 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2244 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2245 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2246 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2233 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3639  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2233 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2234 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N412 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3638  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n466 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n434 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2877 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2870 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3637  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2863 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2864 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2865 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2861 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3636  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2870 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2871 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2872 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2873 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2860 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3635  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2861 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N344 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3634  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n467 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n435 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2232 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2225 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3633  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2217 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2218 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2219 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2220 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2216 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3632  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2225 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2226 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2227 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2228 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2215 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3631  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2215 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2216 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N413 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3630  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n467 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n435 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2859 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2852 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3629  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2844 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2845 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2846 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2847 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2843 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3628  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2852 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2853 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2854 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2855 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2842 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3627  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2842 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2843 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N345 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3626  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n468 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n436 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2214 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2207 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3625  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2199 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2200 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2201 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2202 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2198 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3624  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2207 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2208 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2209 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2210 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2197 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3623  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2197 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2198 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N414 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3622  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n468 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n436 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2841 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2834 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3621  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2826 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2827 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2828 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2829 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2825 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3620  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2835 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2836 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2837 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2824 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3619  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2824 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2825 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N346 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3618  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n469 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n437 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2196 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2189 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3617  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2181 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2182 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2183 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2184 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2180 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3616  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2189 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2190 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2191 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2192 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2179 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3615  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2179 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2180 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N415 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3614  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n469 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n437 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2823 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2816 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3613  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2809 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2810 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2811 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2807 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3612  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2816 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2817 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2818 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2819 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2806 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3611  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2807 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N347 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3610  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n470 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n438 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2178 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2171 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3609  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2163 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2164 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2165 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2166 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2162 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3608  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2171 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2172 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2173 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2174 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2161 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3607  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2161 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2162 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N416 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3606  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n470 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n438 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2805 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2798 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3605  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2790 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2791 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2792 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2793 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2789 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3604  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2798 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2799 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2800 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2801 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2788 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3603  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2788 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2789 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N348 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3602  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n471 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n439 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2153 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3601  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2145 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2146 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2147 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2148 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2144 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3600  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2153 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2154 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2155 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2143 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3599  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2143 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2144 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N417 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3598  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n471 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n439 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2787 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2780 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3597  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2772 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2773 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2774 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2775 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2771 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3596  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2781 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2782 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2783 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2770 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3595  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2770 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2771 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N349 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3594  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n472 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n440 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2142 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2135 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3593  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2127 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2128 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2129 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2130 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2126 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3592  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2135 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2136 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2137 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2138 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2125 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3591  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2125 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2126 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N418 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3590  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n472 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n440 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2769 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2762 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3589  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2755 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2756 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2757 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2753 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3588  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2762 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2763 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2764 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2765 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2752 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3587  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2753 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N350 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3586  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n473 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n441 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2124 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2117 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3585  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2109 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2110 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2111 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2112 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2108 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3584  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2117 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2118 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2119 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2120 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2107 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3583  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2107 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2108 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N419 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3582  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n473 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n441 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2751 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2744 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3581  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2736 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2737 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2738 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2739 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2735 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3580  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2744 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2745 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2746 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2747 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2734 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3579  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2734 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2735 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N351 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3578  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n474 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n442 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2106 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2099 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3577  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2091 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2092 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2093 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2094 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2090 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3576  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2099 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2100 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2101 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2102 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2089 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3575  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2089 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2090 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N420 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3574  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n474 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n442 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2733 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2726 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3573  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2718 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2719 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2720 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2721 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2717 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3572  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2727 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2728 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2729 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2716 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3571  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2716 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2717 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N352 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3570  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n475 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n443 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2088 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2081 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3569  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2073 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2074 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2075 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2076 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2072 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3568  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2081 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2082 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2083 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2084 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2071 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3567  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2071 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2072 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N421 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3566  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n475 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n443 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2715 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2708 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3565  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2701 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2702 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2703 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2699 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3564  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2708 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2709 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2710 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2711 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2698 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3563  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2699 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N353 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3562  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n476 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n444 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2070 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2063 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3561  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2055 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2056 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2057 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2058 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2054 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3560  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2063 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2064 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2065 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2066 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2053 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3559  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2053 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2054 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N422 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3558  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n476 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n444 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2697 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2690 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3557  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2682 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2683 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2684 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2685 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2681 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3556  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2690 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2691 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2692 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2693 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2680 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3555  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2680 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2681 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N354 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3554  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n477 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n445 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2052 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2045 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3553  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2037 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2038 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2039 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2040 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2036 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3552  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2045 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2046 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2047 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2048 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2035 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3551  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2035 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2036 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N423 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3550  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n477 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n445 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2679 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2672 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3549  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2664 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2665 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2666 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2667 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2663 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3548  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2672 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2673 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2674 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2675 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2662 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3547  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2662 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2663 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N355 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3546  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n478 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n446 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2034 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2027 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3545  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2019 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2020 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2021 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2022 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2018 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3544  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2027 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2028 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2029 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2030 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2017 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3543  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2017 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2018 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N424 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3542  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n478 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n446 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2661 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2654 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3541  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2646 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2647 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2648 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2649 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2645 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3540  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2654 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2655 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2656 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2657 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2644 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3539  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2644 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2645 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N356 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3538  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n479 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n447 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2016 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2009 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3537  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2001 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2002 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2003 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2004 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2000 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3536  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2009 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2010 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2011 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2012 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1999 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3535  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1999 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2000 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N425 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3534  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n479 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n447 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2643 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2636 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3533  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2628 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2629 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2630 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2631 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2627 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3532  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2636 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2637 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2638 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2639 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2626 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3531  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2626 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2627 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N357 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3530  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n480 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n448 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1998 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1991 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3529  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1983 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1984 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1985 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1986 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1982 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3528  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1991 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1992 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1993 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1994 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1981 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3527  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1981 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1982 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N426 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3526  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n480 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n448 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2625 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2618 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3525  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2610 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2611 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2612 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2613 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2609 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3524  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2618 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2619 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2620 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2621 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2608 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3523  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2608 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2609 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N358 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3522  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n481 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n449 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1977 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1955 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3521  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1929 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1930 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1931 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1932 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1928 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3520  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1955 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1956 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1957 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1958 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1927 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3519  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1927 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1928 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N427 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3518  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n481 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n449 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2604 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2582 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3517  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2556 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2557 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2558 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2559 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2555 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3516  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2582 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2583 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2584 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2585 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2554 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3515  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2554 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2555 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/N359 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3514  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][20] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2332 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3513  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1037 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1005 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2332 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2325 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3512  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][20] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2959 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3511  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1037 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1005 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2959 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2952 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3510  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][19] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2314 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3509  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1038 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1006 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2314 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2307 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3508  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][19] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2941 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3507  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1038 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1006 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2941 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2934 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3506  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][18] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2296 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3505  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1039 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1007 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2296 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2289 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3504  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][18] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2923 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3503  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1039 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1007 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2923 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2916 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3502  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][17] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2278 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3501  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1040 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1008 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2278 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2271 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3500  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][17] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2905 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3499  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1040 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1008 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2905 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2898 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3498  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][16] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2260 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3497  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1041 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1009 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2260 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2253 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3496  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][16] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2887 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3495  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1041 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1009 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2887 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2880 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3494  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][15] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2242 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3493  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1042 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1010 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2242 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2235 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3492  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][15] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2869 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3491  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1042 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1010 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2869 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2862 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3490  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][14] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2224 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3489  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1043 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1011 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2224 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2217 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3488  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][14] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2851 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3487  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1043 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1011 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2851 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2844 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3486  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][13] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2206 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3485  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1044 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1012 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2206 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2199 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3484  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][13] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2833 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3483  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1044 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1012 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2833 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2826 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3482  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][12] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2188 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3481  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1045 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1013 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2188 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2181 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3480  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][12] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2815 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3479  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1045 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1013 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2815 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2808 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3478  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][11] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2170 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3477  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1046 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1014 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2170 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2163 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3476  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][11] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2797 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3475  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1046 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1014 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2797 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2790 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3474  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][10] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2152 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3473  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1047 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1015 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2152 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2145 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3472  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][10] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2779 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3471  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1047 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1015 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2779 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2772 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3470  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2339 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3469  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n333 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n301 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2339 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2334 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3468  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2331 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3467  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n973 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n941 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2331 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2326 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3466  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2966 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3465  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n333 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n301 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2966 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2961 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3464  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2958 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3463  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n973 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n941 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2958 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2953 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3462  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2321 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3461  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n334 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n302 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2321 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2316 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3460  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2313 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3459  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n974 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n942 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2313 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2308 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3458  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2948 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3457  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n334 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n302 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2948 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2943 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3456  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2940 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3455  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n974 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n942 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2940 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2935 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3454  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2303 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3453  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n335 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n303 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2303 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2298 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3452  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2295 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3451  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n975 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n943 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2295 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2290 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3450  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2930 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3449  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n335 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n303 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2930 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2925 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3448  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2922 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3447  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n975 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n943 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2922 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2917 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3446  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2285 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3445  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n336 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n304 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2285 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2280 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3444  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2277 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3443  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n976 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n944 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2277 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2272 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3442  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2912 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3441  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n336 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n304 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2912 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2907 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3440  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2904 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3439  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n976 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n944 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2904 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2899 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3438  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2267 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3437  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n337 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n305 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2267 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2262 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3436  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2259 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3435  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n977 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n945 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2259 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2254 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3434  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2894 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3433  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n337 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n305 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2894 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2889 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3432  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2886 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3431  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n977 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n945 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2886 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2881 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3430  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2249 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3429  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n338 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n306 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2249 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2244 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3428  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2241 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3427  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n978 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n946 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2241 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2236 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3426  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2876 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3425  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n338 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n306 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2876 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2871 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3424  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2868 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3423  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n978 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n946 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2868 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2863 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3422  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2231 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3421  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n339 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n307 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2231 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2226 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3420  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2223 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3419  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n979 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n947 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2223 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2218 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3418  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2858 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3417  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n339 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n307 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2858 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2853 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3416  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2850 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3415  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n979 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n947 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2850 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2845 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3414  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2213 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3413  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n340 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n308 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2213 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2208 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3412  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2205 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3411  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n980 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n948 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2205 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2200 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3410  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2840 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3409  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n340 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n308 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2840 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2835 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3408  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2832 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3407  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n980 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n948 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2832 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2827 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3406  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2195 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3405  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n341 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n309 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2195 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2190 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3404  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2187 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3403  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n981 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n949 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2187 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2182 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3402  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2822 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3401  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n341 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n309 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2822 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2817 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3400  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2814 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3399  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n981 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n949 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2814 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2809 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3398  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2177 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3397  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n342 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n310 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2177 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2172 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3396  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2169 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3395  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n982 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n950 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2169 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2164 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3394  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2804 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3393  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n342 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n310 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2804 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2799 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3392  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2796 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3391  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n982 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n950 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2796 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2791 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3390  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2159 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3389  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n343 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n311 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2154 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3388  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2151 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3387  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n983 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n951 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2151 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2146 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3386  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2786 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3385  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n343 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n311 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2786 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2781 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3384  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2778 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3383  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n983 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n951 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2778 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2773 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3382  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][9] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2134 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3381  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1048 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1016 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2134 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2127 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3380  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][9] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2761 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3379  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1048 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1016 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2761 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2754 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3378  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][8] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2116 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3377  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1049 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1017 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2116 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2109 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3376  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][8] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2743 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3375  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1049 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1017 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2743 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2736 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3374  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][7] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2098 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3373  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1050 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1018 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2098 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2091 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3372  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][7] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2725 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3371  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1050 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1018 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2725 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2718 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3370  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][6] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2080 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3369  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1051 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1019 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2080 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2073 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3368  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][6] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2707 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3367  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1051 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1019 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2707 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2700 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3366  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][5] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2062 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3365  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1052 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1020 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2062 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2055 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3364  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][5] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2689 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3363  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1052 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1020 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2689 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2682 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3362  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][4] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2044 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3361  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1053 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1021 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2044 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2037 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3360  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][4] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2671 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3359  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1053 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1021 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2671 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2664 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3358  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][3] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2026 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3357  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1054 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1022 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2026 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2019 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3356  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][3] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2653 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3355  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1054 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1022 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2653 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2646 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3354  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][2] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2008 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3353  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1055 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1023 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2008 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2001 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3352  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][2] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2635 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3351  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1055 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1023 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2635 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2628 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3350  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][1] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1990 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3349  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1056 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1024 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1990 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1983 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3348  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][1] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2617 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3347  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1056 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1024 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2617 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2610 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3346  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][0] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1951 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3345  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1057 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1025 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1951 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1929 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3344  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][0] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2578 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3343  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1057 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1025 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2578 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2556 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3342  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][31] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2540 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3341  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1026 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n994 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2540 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2523 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3340  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][31] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3167 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3339  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1026 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n994 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3167 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3150 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3338  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][30] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2512 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3337  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1027 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n995 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2512 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2505 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3336  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][30] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3139 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3335  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1027 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n995 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3139 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3132 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3334  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][29] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2494 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3333  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1028 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n996 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2494 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2487 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3332  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][29] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3121 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3331  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1028 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n996 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3121 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3114 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3330  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][28] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2476 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3329  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1029 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n997 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2476 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2469 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3328  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][28] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3103 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3327  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1029 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n997 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3103 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3096 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3326  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][27] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2458 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3325  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1030 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n998 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2458 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2451 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3324  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][27] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3085 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3323  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1030 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n998 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3085 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3078 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3322  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][26] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2440 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3321  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1031 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n999 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2440 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2433 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3320  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][26] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3067 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3319  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1031 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n999 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3067 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3060 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3318  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][25] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2422 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3317  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1032 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1000 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2422 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2415 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3316  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][25] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3049 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3315  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1032 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1000 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3049 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3042 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3314  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][24] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2404 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3313  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1033 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1001 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2404 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2397 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3312  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][24] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3031 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3311  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1033 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1001 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3031 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3024 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3310  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][23] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2386 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3309  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1034 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1002 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2386 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2379 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3308  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][23] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3013 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3307  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1034 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1002 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3013 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3006 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3306  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][22] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2368 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3305  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1035 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1003 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2368 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2361 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3304  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][22] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2995 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3303  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1035 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1003 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2995 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2988 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3302  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][21] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2350 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3301  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1036 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1004 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2350 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2343 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3300  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][21] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2977 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3299  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1036 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1004 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2977 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2970 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3298  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2141 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3297  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n344 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n312 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2141 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2136 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3296  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2133 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3295  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n984 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n952 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2133 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2128 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3294  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2768 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3293  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n344 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n312 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2768 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2763 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3292  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2760 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3291  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n984 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n952 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2760 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2755 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3290  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2123 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3289  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n345 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n313 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2123 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2118 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3288  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2115 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3287  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n985 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n953 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2115 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2110 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3286  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2750 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3285  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n345 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n313 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2750 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2745 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3284  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2742 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3283  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n985 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n953 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2742 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2737 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3282  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2105 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3281  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n346 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n314 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2105 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2100 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3280  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2097 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3279  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n986 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n954 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2097 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2092 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3278  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2732 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3277  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n346 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n314 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2732 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2727 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3276  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2724 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3275  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n986 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n954 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2724 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2719 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3274  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2087 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3273  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n347 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n315 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2087 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2082 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3272  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2079 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3271  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n987 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n955 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2079 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2074 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3270  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2714 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3269  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n347 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n315 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2714 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2709 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3268  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2706 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3267  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n987 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n955 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2706 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2701 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3266  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2069 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3265  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n348 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n316 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2069 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2064 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3264  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2061 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3263  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n988 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n956 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2061 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2056 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3262  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2696 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3261  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n348 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n316 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2696 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2691 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3260  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2688 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3259  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n988 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n956 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2688 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2683 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3258  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2051 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3257  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n349 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n317 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2051 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2046 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3256  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2043 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3255  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n989 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n957 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2043 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2038 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3254  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2678 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3253  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n349 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n317 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2678 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2673 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3252  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2670 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3251  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n989 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n957 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2670 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2665 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3250  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2033 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3249  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n350 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n318 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2033 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2028 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3248  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2025 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3247  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n990 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n958 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2025 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2020 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3246  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2660 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3245  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n350 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n318 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2660 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2655 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3244  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2652 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3243  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n990 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n958 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2652 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2647 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3242  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2015 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3241  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n351 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n319 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2015 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2010 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3240  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2007 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3239  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n991 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n959 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2007 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2002 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3238  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2642 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3237  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n351 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n319 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2642 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2637 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3236  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2634 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3235  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n991 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n959 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2634 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2629 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3234  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1997 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3233  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n352 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n320 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1997 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1992 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3232  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1989 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3231  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n992 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n960 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1989 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1984 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3230  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2624 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3229  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n352 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n320 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2624 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2619 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3228  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2616 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3227  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n992 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n960 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2616 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2611 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3226  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1972 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3225  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n353 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n321 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1972 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1956 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3224  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1946 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3223  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n993 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n961 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1946 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1930 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3222  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2599 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3221  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n353 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n321 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2599 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2583 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3220  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2573 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3219  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n993 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n961 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2573 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2557 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3218  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2550 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3217  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n322 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n290 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2550 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2542 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3216  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2537 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3215  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n962 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n930 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2537 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2524 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3214  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3177 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3213  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n322 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n290 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3177 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3169 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3212  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3164 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3211  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n962 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n930 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3164 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3151 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3210  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2519 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3209  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n323 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n291 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2519 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2514 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3208  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2511 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3207  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n963 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n931 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2511 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2506 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3206  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3146 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3205  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n323 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n291 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3146 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3141 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3204  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3138 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3203  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n963 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n931 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3138 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3133 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3202  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2501 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3201  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n324 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n292 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2501 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2496 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3200  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2493 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3199  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n964 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n932 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2493 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2488 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3198  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3128 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3197  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n324 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n292 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3128 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3123 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3196  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3120 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3195  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n964 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n932 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3120 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3115 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3194  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2483 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3193  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n325 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n293 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2483 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2478 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3192  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2475 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3191  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n965 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n933 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2475 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2470 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3190  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3110 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3189  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n325 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n293 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3110 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3105 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3188  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3102 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3187  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n965 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n933 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3102 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3097 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3186  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2465 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3185  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n326 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n294 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2465 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2460 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3184  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2457 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3183  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n966 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n934 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2457 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2452 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3182  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3092 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3181  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n326 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n294 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3092 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3087 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3180  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3084 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3179  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n966 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n934 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3084 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3079 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3178  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2447 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3177  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n327 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n295 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2447 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2442 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3176  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2439 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3175  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n967 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n935 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2439 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2434 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3174  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3074 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3173  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n327 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n295 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3074 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3069 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3172  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3066 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3171  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n967 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n935 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3066 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3061 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3170  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2429 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3169  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n328 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n296 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2429 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2424 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3168  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2421 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3167  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n968 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n936 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2421 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2416 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3166  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3056 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3165  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n328 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n296 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3056 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3051 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3164  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3048 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3163  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n968 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n936 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3048 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3043 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3162  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2411 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3161  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n329 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n297 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2411 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2406 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3160  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2403 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3159  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n969 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n937 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2403 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2398 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3158  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3038 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3157  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n329 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n297 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3038 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3033 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3156  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3030 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3155  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n969 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n937 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3030 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3025 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3154  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2393 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3153  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n330 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n298 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2393 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2388 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3152  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2385 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3151  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n970 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n938 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2385 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2380 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3150  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3020 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3149  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n330 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n298 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3020 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3015 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3148  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3012 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3147  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n970 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n938 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3012 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3007 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3146  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2375 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3145  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n331 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n299 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2375 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2370 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3144  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2367 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3143  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n971 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n939 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2367 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2362 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3142  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3002 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3141  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n331 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n299 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3002 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2997 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3140  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2994 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3139  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n971 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n939 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2994 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2989 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3138  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2357 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3137  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n332 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n300 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2357 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2352 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3136  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2349 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3135  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n972 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n940 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2349 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2344 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3134  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2984 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3133  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n332 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n300 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2984 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2979 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3132  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2976 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3131  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n972 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n940 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2976 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2971 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3130  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][20] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2338 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3129  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n173 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n141 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2338 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2335 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3128  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][20] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2330 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3127  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n717 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2330 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2327 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3126  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][20] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2965 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3125  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n173 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n141 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2965 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2962 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3124  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][20] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2957 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3123  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n749 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n717 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2957 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2954 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3122  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][19] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2320 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3121  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n174 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n142 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2320 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2317 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3120  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][19] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2312 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3119  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n718 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2312 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2309 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3118  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][19] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2947 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3117  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n174 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n142 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2947 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2944 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3116  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][19] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2939 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3115  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n750 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n718 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2939 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2936 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3114  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][18] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2302 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3113  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n175 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n143 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2302 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2299 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3112  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][18] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2294 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3111  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2294 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2291 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3110  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][18] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2929 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3109  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n175 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n143 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2929 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2926 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3108  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][18] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2921 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3107  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n751 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2921 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2918 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3106  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][17] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2284 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3105  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n176 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n144 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2284 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2281 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3104  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][17] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2276 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3103  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n752 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2276 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2273 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3102  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][17] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2911 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3101  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n176 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n144 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2911 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2908 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3100  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][17] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2903 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3099  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n752 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2903 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2900 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3098  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][16] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2266 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3097  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n177 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n145 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2266 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2263 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3096  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][16] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2258 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3095  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n753 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2258 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2255 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3094  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][16] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2893 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3093  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n177 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n145 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2893 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2890 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3092  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][16] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2885 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3091  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n753 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2885 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2882 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3090  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][15] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2248 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3089  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n178 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n146 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2248 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2245 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3088  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][15] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2240 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3087  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n754 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n722 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2240 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2237 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3086  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][15] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2875 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3085  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n178 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n146 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2875 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2872 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3084  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][15] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2867 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3083  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n754 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n722 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2867 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2864 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3082  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][14] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2230 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3081  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n179 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n147 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2230 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2227 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3080  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][14] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2222 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3079  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n755 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n723 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2222 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2219 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3078  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][14] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2857 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3077  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n179 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n147 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2857 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2854 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3076  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][14] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2849 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3075  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n755 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n723 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2849 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2846 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3074  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][13] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2212 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3073  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n180 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n148 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2212 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2209 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3072  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][13] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2204 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3071  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n756 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n724 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2204 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2201 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3070  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][13] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2839 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3069  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n180 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n148 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2839 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2836 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3068  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][13] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2831 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3067  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n756 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n724 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2831 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2828 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3066  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][12] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2194 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3065  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n181 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n149 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2194 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2191 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3064  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][12] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2186 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3063  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n757 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n725 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2186 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2183 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3062  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][12] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2821 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3061  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n181 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n149 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2821 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2818 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3060  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][12] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2813 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3059  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n757 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n725 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2813 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2810 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3058  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][11] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2176 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3057  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n182 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n150 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2176 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2173 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3056  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][11] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2168 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3055  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n758 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n726 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2168 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2165 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3054  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][11] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2803 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3053  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n182 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n150 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2803 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2800 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3052  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][11] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2795 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3051  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n758 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n726 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2795 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2792 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3050  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][10] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2158 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3049  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n183 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n151 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2158 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2155 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3048  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][10] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2150 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3047  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n759 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n727 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2150 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2147 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3046  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][10] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2785 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3045  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n183 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n151 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2785 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2782 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3044  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][10] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2777 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3043  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n759 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n727 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2777 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2774 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3042  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][9] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2140 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3041  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n184 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n152 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2140 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2137 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3040  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][9] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2132 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3039  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n760 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n728 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2132 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2129 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3038  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][9] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2767 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3037  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n184 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n152 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2767 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2764 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3036  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][9] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2759 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3035  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n760 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n728 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2759 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2756 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3034  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][8] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2122 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3033  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n185 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n153 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2122 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2119 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3032  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][8] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2114 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3031  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n729 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2114 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2111 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3030  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][8] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2749 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3029  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n185 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n153 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2749 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2746 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3028  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][8] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2741 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3027  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n761 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n729 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2741 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2738 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3026  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][7] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2104 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3025  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n186 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n154 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2104 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2101 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3024  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][7] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2096 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3023  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n730 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2096 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2093 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3022  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][7] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2731 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3021  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n186 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n154 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2731 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2728 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3020  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][7] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2723 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3019  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n762 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n730 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2723 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2720 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3018  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][6] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2086 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3017  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n187 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n155 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2086 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2083 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3016  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][6] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2078 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3015  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n731 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2078 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2075 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3014  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][6] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2713 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3013  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n187 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n155 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2713 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2710 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3012  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][6] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2705 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3011  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n763 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n731 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2705 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2702 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3010  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][5] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2068 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3009  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n188 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n156 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2068 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2065 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3008  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][5] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2060 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3007  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n764 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n732 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2060 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2057 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3006  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][5] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2695 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3005  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n188 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n156 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2695 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2692 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3004  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][5] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2687 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3003  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n764 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n732 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2687 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2684 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3002  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][4] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2050 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3001  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n189 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n157 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2050 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2047 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3000  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][4] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2042 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2999  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n765 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n733 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2042 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2039 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2998  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][4] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2677 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2997  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n189 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n157 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2677 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2674 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2996  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][4] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2669 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2995  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n765 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n733 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2669 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2666 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2994  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][3] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2032 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2993  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n190 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n158 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2032 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2029 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2992  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][3] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2024 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2991  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n766 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n734 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2024 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2021 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2990  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][3] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2659 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2989  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n190 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n158 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2659 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2656 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2988  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][3] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2651 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2987  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n766 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n734 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2651 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2648 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2986  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][2] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2014 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2985  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n191 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n159 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2014 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2011 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2984  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][2] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2006 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2983  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n767 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n735 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2006 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2003 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2982  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][2] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2641 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2981  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n191 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n159 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2641 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2638 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2980  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][2] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2633 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2979  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n767 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n735 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2633 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2630 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2978  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][1] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1996 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2977  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n192 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n160 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1996 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1993 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2976  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][1] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1988 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2975  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n768 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n736 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1988 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1985 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2974  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][1] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2623 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2973  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n192 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n160 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2623 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2620 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2972  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][1] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2615 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2971  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n768 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n736 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2615 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2612 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2970  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][0] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1966 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2969  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n193 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n161 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1966 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1957 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2968  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][0] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1940 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2967  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n769 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n737 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1940 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1931 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2966  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][0] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2593 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2965  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n193 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n161 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2593 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2584 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2964  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][0] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2567 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2963  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n769 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n737 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2567 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2558 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2962  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][31] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2547 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2961  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n162 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n130 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2547 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2543 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2960  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][31] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2534 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2959  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n738 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n706 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2534 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2525 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2958  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][31] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3174 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2957  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n162 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n130 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3174 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3170 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2956  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][31] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3161 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2955  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n738 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n706 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3161 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3152 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2954  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][30] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2518 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2953  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n163 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n131 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2518 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2515 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2952  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][30] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2510 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2951  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n739 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n707 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2510 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2507 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2950  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][30] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3145 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2949  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n163 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n131 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3145 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3142 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2948  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][30] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3137 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2947  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n739 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n707 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3137 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3134 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2946  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][29] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2500 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2945  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n164 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n132 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2500 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2497 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2944  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][29] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2492 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2943  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n740 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n708 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2492 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2489 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2942  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][29] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3127 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2941  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n164 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n132 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3127 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3124 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2940  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][29] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3119 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2939  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n740 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n708 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3119 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3116 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2938  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][28] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2482 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2937  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n165 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n133 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2482 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2479 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2936  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][28] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2474 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2935  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n741 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n709 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2474 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2471 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2934  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][28] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3109 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2933  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n165 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n133 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3109 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3106 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2932  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][28] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3101 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2931  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n741 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n709 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3101 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3098 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2930  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][27] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2464 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2929  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n166 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n134 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2464 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2461 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2928  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][27] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2456 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2927  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n742 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n710 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2456 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2453 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2926  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][27] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3091 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2925  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n166 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n134 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3091 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3088 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2924  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][27] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3083 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2923  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n742 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n710 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3083 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3080 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2922  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][26] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2446 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2921  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n167 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n135 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2446 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2443 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2920  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][26] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2438 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2919  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n743 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n711 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2438 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2435 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2918  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][26] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3073 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2917  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n167 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n135 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3073 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3070 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2916  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][26] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3065 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2915  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n743 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n711 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3065 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3062 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2914  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][25] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2428 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2913  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n168 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n136 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2428 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2425 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2912  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][25] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2420 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2911  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n744 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n712 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2420 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2417 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2910  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][25] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3055 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2909  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n168 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n136 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3055 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3052 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2908  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][25] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3047 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2907  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n744 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n712 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3047 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3044 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2906  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][24] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2410 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2905  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n169 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n137 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2410 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2407 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2904  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][24] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2402 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2903  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n745 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n713 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2402 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2399 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2902  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][24] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3037 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2901  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n169 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n137 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3037 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3034 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2900  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][24] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3029 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2899  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n745 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n713 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3029 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3026 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2898  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][23] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2392 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2897  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n170 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n138 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2392 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2389 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2896  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][23] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2384 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2895  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n746 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n714 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2384 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2381 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2894  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][23] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3019 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2893  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n170 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n138 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3019 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3016 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2892  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][23] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3011 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2891  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n746 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n714 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3011 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3008 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2890  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][22] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2374 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2889  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n171 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n139 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2374 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2371 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2888  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][22] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2366 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2887  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n747 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n715 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2366 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2363 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2886  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][22] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3001 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2885  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n171 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n139 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3001 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2998 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2884  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][22] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2993 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2883  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n747 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n715 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2993 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2990 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2882  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][21] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2356 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2881  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n172 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n140 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2356 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2353 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2880  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][21] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2348 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2879  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n748 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n716 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2348 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2345 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2878  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][21] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2983 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2877  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n172 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n140 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2983 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2980 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2876  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][21] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2975 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2875  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n748 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n716 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2975 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2972 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2874  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2337 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2873  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n45 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n13 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2337 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2336 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2872  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2329 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2871  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n621 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n589 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2329 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2328 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2870  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2964 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2869  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n45 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n13 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2964 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2963 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2868  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2956 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2867  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n621 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n589 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2956 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2955 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2866  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2319 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2865  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n46 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n14 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2319 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2318 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2864  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2311 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2863  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n622 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n590 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2311 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2310 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2862  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2946 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2861  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n46 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n14 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2946 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2945 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2860  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2938 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2859  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n622 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n590 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2938 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2937 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2858  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2301 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2857  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n47 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n15 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2301 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2300 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2856  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2293 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2855  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n623 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n591 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2293 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2292 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2854  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2928 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2853  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n47 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n15 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2928 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2927 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2852  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2920 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2851  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n623 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n591 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2920 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2919 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2850  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2283 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2849  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n48 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n16 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2283 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2282 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2848  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2275 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2847  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n624 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n592 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2275 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2274 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2846  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2910 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2845  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n48 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n16 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2910 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2909 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2844  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2902 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2843  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n624 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n592 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2902 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2901 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2842  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2265 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2841  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n49 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n17 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2265 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2264 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2840  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2257 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2839  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n625 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n593 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2257 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2256 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2838  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2892 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2837  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n49 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n17 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2892 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2891 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2836  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2884 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2835  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n625 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n593 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2884 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2883 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2834  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2247 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2833  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n50 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n18 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2247 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2246 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2832  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2239 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2831  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n626 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n594 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2239 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2238 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2830  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2874 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2829  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n50 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n18 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2874 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2873 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2828  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2866 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2827  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n626 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n594 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2866 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2865 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2826  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2229 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2825  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n51 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n19 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2229 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2228 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2824  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2221 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2823  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n627 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n595 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2221 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2220 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2822  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2856 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2821  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n51 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n19 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2856 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2855 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2820  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2848 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2819  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n627 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n595 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2848 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2847 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2818  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2211 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2817  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n52 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n20 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2211 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2210 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2816  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2203 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2815  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n628 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n596 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2203 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2202 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2814  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2838 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2813  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n52 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n20 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2838 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2837 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2812  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2830 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2811  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n628 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n596 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2830 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2829 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2810  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2193 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2809  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n53 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n21 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2193 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2192 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2808  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2185 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2807  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n629 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n597 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2185 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2184 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2806  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2820 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2805  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n53 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n21 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2820 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2819 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2804  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2812 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2803  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n629 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n597 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2812 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2811 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2802  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2175 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2801  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n54 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n22 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2175 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2174 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2800  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2167 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2799  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n630 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n598 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2167 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2166 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2798  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2802 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2797  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n54 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n22 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2802 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2801 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2796  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2794 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2795  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n630 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n598 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2794 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2793 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2794  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2157 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2793  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n55 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n23 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2156 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2792  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2149 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2791  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n631 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n599 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2149 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2148 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2790  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2784 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2789  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n55 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n23 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2784 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2783 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2788  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2776 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2787  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n631 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n599 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2776 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2775 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2786  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2139 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2785  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n56 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n24 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2139 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2138 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2784  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2131 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2783  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n632 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n600 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2131 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2130 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2782  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2766 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2781  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n56 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n24 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2766 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2765 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2780  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2758 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2779  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n632 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n600 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2758 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2757 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2778  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2121 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2777  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n57 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n25 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2121 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2120 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2776  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2113 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2775  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n633 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n601 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2113 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2112 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2774  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2748 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2773  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n57 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n25 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2748 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2747 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2772  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2740 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2771  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n633 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n601 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2740 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2739 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2770  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2103 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2769  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n58 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n26 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2103 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2102 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2768  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2095 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2767  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n634 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n602 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2095 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2094 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2766  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2730 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2765  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n58 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n26 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2730 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2729 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2764  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2722 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2763  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n634 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n602 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2722 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2721 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2762  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2085 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2761  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n59 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n27 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2085 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2084 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2760  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2077 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2759  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n635 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n603 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2077 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2076 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2758  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2712 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2757  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n59 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n27 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2712 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2711 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2756  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2704 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2755  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n635 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n603 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2704 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2703 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2754  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2067 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2753  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n60 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n28 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2067 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2066 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2752  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2059 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2751  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n636 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n604 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2059 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2058 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2750  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2694 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2749  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n60 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n28 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2694 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2693 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2748  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2686 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2747  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n636 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n604 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2686 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2685 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2746  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2049 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2745  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n61 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n29 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2049 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2048 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2744  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2041 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2743  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n637 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n605 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2041 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2040 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2742  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2676 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2741  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n61 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n29 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2676 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2675 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2740  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2668 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2739  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n637 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n605 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2668 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2667 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2738  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2031 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2737  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n62 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n30 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2031 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2030 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2736  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2023 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2735  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n638 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n606 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2023 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2022 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2734  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2658 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2733  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n62 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n30 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2658 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2657 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2732  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2650 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2731  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n638 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n606 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2650 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2649 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2730  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2013 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2729  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n63 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n31 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2013 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2012 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2728  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2005 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2727  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n639 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n607 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2005 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2004 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2726  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2640 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2725  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n63 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n31 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2640 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2639 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2724  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2632 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2723  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n639 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n607 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2632 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2631 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2722  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1995 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2721  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n64 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n32 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1995 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1994 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2720  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1987 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2719  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n640 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n608 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1987 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1986 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2718  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2622 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2717  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n64 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n32 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2622 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2621 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2716  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2614 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2715  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n640 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n608 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2614 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2613 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2714  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1961 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2713  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n65 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n33 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1961 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1958 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2712  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1935 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2711  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n641 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n609 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1935 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1932 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2710  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2588 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2709  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n65 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n33 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2588 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2585 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2708  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2562 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2707  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n641 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n609 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2562 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2559 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2706  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2545 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2705  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n34 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2545 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2544 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2704  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2527 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2703  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n610 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n578 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2527 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2526 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2702  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3172 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2701  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n34 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3172 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3171 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2700  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3154 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2699  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n610 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n578 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3154 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3153 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2698  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2517 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2697  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n35 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2517 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2516 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2696  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2509 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2695  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n611 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n579 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2509 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2508 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2694  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3144 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2693  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n35 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3144 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3143 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2692  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3136 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2691  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n611 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n579 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3136 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3135 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2690  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2499 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2689  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n36 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2499 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2498 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2688  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2491 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2687  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n612 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n580 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2491 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2490 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2686  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3126 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2685  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n36 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3126 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3125 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2684  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3118 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2683  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n612 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n580 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3118 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3117 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2682  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2481 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2681  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n37 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n5 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2481 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2480 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2680  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2473 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2679  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n613 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n581 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2473 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2472 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2678  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3108 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2677  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n37 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n5 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3108 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3107 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2676  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3100 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2675  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n613 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n581 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3100 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3099 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2674  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2463 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2673  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n38 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n6 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2463 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2462 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2672  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2455 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2671  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n614 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n582 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2455 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2454 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2670  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3090 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2669  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n38 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n6 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3090 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3089 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2668  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3082 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2667  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n614 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n582 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3082 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3081 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2666  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2445 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2665  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n39 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n7 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2445 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2444 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2664  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2437 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2663  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n615 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n583 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2437 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2436 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2662  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3072 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2661  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n39 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n7 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3072 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3071 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2660  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3064 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2659  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n615 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n583 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3064 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3063 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2658  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2427 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2657  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n40 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n8 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2427 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2426 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2656  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2419 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2655  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n616 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n584 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2419 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2418 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2654  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3054 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2653  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n40 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n8 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3054 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3053 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2652  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3046 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2651  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n616 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n584 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3046 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3045 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2650  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2409 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2649  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n41 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n9 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2409 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2408 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2648  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2401 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2647  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n617 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n585 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2401 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2400 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2646  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3036 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2645  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n41 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n9 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3036 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3035 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2644  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3028 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2643  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n617 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n585 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3028 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3027 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2642  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2391 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2641  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n42 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n10 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2391 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2390 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2640  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2383 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2639  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n618 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n586 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2383 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2382 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2638  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3018 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2637  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n42 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n10 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3018 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3017 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2636  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3010 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2635  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n618 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n586 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3010 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3009 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2634  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2373 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2633  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n43 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n11 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2373 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2372 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2632  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2365 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2631  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n619 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n587 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2365 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2364 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2630  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3000 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2629  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n43 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n11 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3000 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2999 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2628  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2992 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2627  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n619 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n587 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2992 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2991 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2626  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2355 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2625  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n44 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n12 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2355 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2354 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2624  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2347 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2623  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n620 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n588 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2347 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2346 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2622  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2982 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2621  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n44 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n12 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2982 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2981 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2620  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2974 ) );
  OAI221_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2619  ( .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n620 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n588 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ), .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2974 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2973 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2618  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][31] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2553 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2617  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][31] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][31] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3180 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2616  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][30] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2520 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2615  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][30] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][30] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3147 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2614  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][29] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2502 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2613  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][29] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][29] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3129 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2612  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][28] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2484 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2611  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][28] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][28] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3111 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2610  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][27] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2466 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2609  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][27] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][27] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3093 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2608  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][26] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2448 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2607  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][26] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][26] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3075 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2606  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][25] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2430 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2605  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][25] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][25] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3057 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2604  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][24] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2412 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2603  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][24] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][24] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3039 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2602  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][23] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2394 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2601  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][23] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][23] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3021 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2600  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][22] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2376 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2599  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][22] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][22] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3003 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2598  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][21] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2358 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2597  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][21] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][21] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2985 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2596  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][20] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2340 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2595  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][20] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][20] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2967 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2594  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][19] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2322 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2593  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][19] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][19] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2949 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2592  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][18] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2304 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2591  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][18] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][18] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2931 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2590  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][17] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2286 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2589  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][17] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][17] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2913 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2588  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][16] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2268 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2587  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][16] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][16] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2895 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2586  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][15] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2250 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2585  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][15] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][15] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2877 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2584  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][14] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2232 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2583  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][14] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][14] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2859 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2582  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][13] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2214 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2581  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][13] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][13] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2841 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2580  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][12] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2196 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2579  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][12] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][12] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2823 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2578  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][11] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2178 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2577  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][11] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][11] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2805 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2576  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][10] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2160 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2575  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][10] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][10] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2787 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2574  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][9] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2142 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2573  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][9] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][9] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2769 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2572  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][8] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2124 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2571  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][8] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][8] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2751 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2570  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][7] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2106 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2569  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][7] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][7] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2733 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2568  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][6] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2088 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2567  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][6] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][6] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2715 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2566  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][5] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2070 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2565  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][5] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][5] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2697 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2564  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][4] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2052 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2563  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][4] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][4] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2679 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2562  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][3] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2034 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2561  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][3] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][3] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2661 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2560  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][2] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2016 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2559  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][2] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][2] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2643 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2558  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][1] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1998 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2557  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][1] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][1] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2625 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2556  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][0] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1977 ) );
  AOI222_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2555  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][0] ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][0] ), .C1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ), .C2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2604 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2554  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3932 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1916 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2553  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1916 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n74 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2552  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3932 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1915 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2551  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1915 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n75 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2550  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3932 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1914 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2549  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1914 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n76 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2548  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3932 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1913 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2547  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1913 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n77 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2546  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3931 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1912 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2545  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1912 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n78 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2544  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3931 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1911 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2543  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1911 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n79 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2542  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3931 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1910 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2541  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1910 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n80 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2540  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3931 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1909 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2539  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1909 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n81 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2538  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3931 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1908 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2537  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1908 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n82 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2536  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3930 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1907 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2535  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1907 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n83 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2534  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3930 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1906 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2533  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1906 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n84 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2532  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3930 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1905 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2531  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1905 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n85 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2530  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3930 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1904 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2529  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1904 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n86 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2528  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3930 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1903 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2527  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1903 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n87 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2526  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3929 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1902 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2525  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1902 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n88 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2524  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3929 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1901 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2523  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1901 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n89 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2522  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3929 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1900 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2521  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1900 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n90 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2520  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3929 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1899 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2519  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1899 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n91 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2518  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3929 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1898 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2517  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1898 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n92 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2516  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3928 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1897 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2515  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1897 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n93 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2514  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3928 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1896 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2513  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1896 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n94 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2512  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3928 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1895 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2511  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1895 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n95 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2510  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3928 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1894 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2509  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1894 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n96 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2508  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3928 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1892 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2507  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1892 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n97 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2506  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3941 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1883 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2505  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1883 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n106 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2504  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3941 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1882 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2503  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1882 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n107 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2502  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3941 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1881 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2501  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1881 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n108 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2500  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3941 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1880 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2499  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1880 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n109 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2498  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3940 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1879 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2497  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1879 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n110 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2496  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3940 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1878 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2495  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1878 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n111 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2494  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3940 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1877 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2493  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1877 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n112 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2492  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3940 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1876 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2491  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1876 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n113 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2490  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3940 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1875 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2489  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1875 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n114 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2488  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3939 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1874 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2487  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1874 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n115 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2486  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3939 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1873 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2485  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1873 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n116 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2484  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3939 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1872 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2483  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1872 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n117 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2482  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3939 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1871 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2481  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1871 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n118 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2480  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3939 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1870 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2479  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1870 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n119 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2478  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3938 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1869 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2477  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1869 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n120 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2476  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3938 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1868 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2475  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1868 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n121 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2474  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3938 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1867 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2473  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1867 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n122 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2472  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3938 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1866 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2471  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1866 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n123 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2470  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3938 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1865 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2469  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1865 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n124 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2468  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3937 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1864 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2467  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1864 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n125 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2466  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3937 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1863 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2465  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1863 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n126 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2464  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3937 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1862 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2463  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1862 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n127 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2462  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3937 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1861 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2461  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1861 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n128 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2460  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3937 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1859 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2459  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1859 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n129 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2458  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3968 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1848 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2457  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1848 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n202 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2456  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3968 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1847 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2455  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1847 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n203 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2454  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3968 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1846 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2453  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1846 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n204 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2452  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3968 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1845 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2451  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1845 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n205 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2450  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3967 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1844 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2449  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1844 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n206 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2448  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3967 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1843 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2447  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1843 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n207 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2446  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3967 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1842 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2445  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1842 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n208 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2444  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3967 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1841 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2443  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1841 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n209 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2442  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3967 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1840 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2441  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1840 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n210 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2440  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3966 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1839 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2439  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1839 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n211 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2438  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3966 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1838 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2437  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1838 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n212 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2436  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3966 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1837 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2435  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1837 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n213 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2434  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3966 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1836 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2433  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1836 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n214 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2432  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3966 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1835 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2431  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1835 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n215 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2430  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3965 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1834 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2429  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1834 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n216 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2428  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3965 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1833 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2427  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1833 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n217 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2426  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3965 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1832 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2425  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1832 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n218 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2424  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3965 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1831 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2423  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1831 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n219 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2422  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3965 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1830 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2421  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1830 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n220 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2420  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3964 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1829 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2419  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1829 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n221 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2418  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3964 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1828 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2417  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1828 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n222 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2416  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3964 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1827 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2415  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1827 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n223 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2414  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3964 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1826 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2413  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1826 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n224 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2412  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3964 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1824 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2411  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1824 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n225 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2410  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3977 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1814 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2409  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1814 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n234 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2408  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3977 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1813 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2407  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1813 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n235 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2406  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3977 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1812 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2405  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1812 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n236 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2404  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3977 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1811 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2403  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1811 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n237 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2402  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3976 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1810 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2401  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1810 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n238 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2400  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3976 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1809 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2399  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1809 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n239 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2398  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3976 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1808 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2397  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1808 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n240 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2396  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3976 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1807 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2395  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1807 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n241 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2394  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3976 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1806 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2393  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1806 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n242 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2392  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3975 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1805 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2391  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1805 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n243 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2390  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3975 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1804 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2389  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1804 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n244 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2388  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3975 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1803 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2387  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1803 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n245 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2386  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3975 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1802 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2385  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1802 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n246 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2384  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3975 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1801 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2383  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1801 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n247 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2382  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3974 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1800 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2381  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1800 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n248 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2380  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3974 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1799 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2379  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1799 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n249 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2378  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3974 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1798 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2377  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1798 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n250 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2376  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3974 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1797 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2375  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1797 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n251 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2374  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3974 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1796 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2373  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1796 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n252 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2372  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3973 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1795 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2371  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1795 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n253 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2370  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3973 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1794 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2369  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1794 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n254 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2368  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3973 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1793 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2367  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1793 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n255 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2366  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3973 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1792 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2365  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1792 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n256 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2364  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3973 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1790 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2363  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1790 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n257 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2362  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3986 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1781 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2361  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1781 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n266 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2360  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3986 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1780 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2359  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1780 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n267 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2358  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3986 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1779 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2357  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1779 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n268 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2356  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3986 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1778 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2355  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1778 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n269 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2354  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3985 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1777 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2353  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1777 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n270 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2352  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3985 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1776 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2351  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1776 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n271 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2350  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3985 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1775 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2349  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1775 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n272 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2348  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3985 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1774 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2347  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1774 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n273 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2346  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3985 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1773 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2345  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1773 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n274 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2344  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3984 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1772 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2343  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1772 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n275 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2342  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3984 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1771 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2341  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1771 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n276 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2340  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3984 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1770 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2339  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1770 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n277 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2338  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3984 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1769 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2337  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1769 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n278 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2336  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3984 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1768 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2335  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1768 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n279 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2334  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3983 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1767 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2333  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1767 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n280 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2332  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3983 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1766 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2331  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1766 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n281 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2330  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3983 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1765 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2329  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1765 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n282 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2328  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3983 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1764 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2327  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1764 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n283 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2326  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3983 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1763 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2325  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1763 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n284 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2324  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3982 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1762 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2323  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1762 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n285 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2322  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3982 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1761 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2321  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1761 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n286 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2320  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3982 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1760 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2319  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1760 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n287 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2318  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3982 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1759 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2317  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1759 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n288 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2316  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3982 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1757 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2315  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1757 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n289 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2314  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4013 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1746 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2313  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1746 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n362 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2312  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4013 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1745 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2311  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1745 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n363 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2310  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4013 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1744 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2309  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1744 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n364 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2308  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4013 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1743 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2307  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1743 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n365 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2306  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4012 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1742 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2305  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1742 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n366 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2304  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4012 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1741 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2303  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1741 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n367 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2302  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4012 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1740 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2301  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1740 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n368 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2300  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4012 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1739 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2299  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1739 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n369 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2298  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4012 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1738 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2297  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1738 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n370 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2296  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4011 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1737 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2295  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1737 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n371 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2294  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4011 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1736 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2293  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1736 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n372 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2292  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4011 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1735 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2291  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1735 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n373 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2290  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4011 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1734 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2289  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1734 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n374 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2288  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4011 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1733 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2287  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1733 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n375 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2286  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4010 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1732 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2285  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1732 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n376 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2284  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4010 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1731 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2283  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1731 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n377 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2282  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4010 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1730 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2281  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1730 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n378 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2280  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4010 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1729 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2279  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1729 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n379 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2278  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4010 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1728 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2277  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1728 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n380 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2276  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4009 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1727 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2275  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1727 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n381 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2274  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4009 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1726 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2273  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1726 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n382 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2272  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4009 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1725 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2271  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1725 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n383 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2270  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4009 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1724 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2269  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1724 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n384 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2268  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4009 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1722 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2267  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1722 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n385 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2266  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4021 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1708 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2265  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1708 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n399 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2264  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4021 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1707 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2263  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1707 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n400 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2262  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4021 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1706 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2261  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1706 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n401 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2260  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4021 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1705 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2259  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1705 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n402 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2258  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4020 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1704 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2257  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1704 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n403 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2256  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4020 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1703 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2255  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1703 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n404 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2254  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4020 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1702 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2253  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1702 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n405 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2252  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4020 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1701 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2251  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1701 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n406 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2250  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4020 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1700 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2249  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1700 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n407 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2248  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4018 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1689 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2247  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1689 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n417 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2246  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4048 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1672 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2245  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1672 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n495 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2244  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4048 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1671 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2243  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1671 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n496 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2242  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4048 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1670 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2241  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1670 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n497 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2240  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4048 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1669 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2239  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1669 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n498 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2238  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4047 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1668 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2237  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1668 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n499 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2236  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4047 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1667 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2235  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1667 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n500 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2234  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4047 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1666 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2233  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1666 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n501 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2232  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4047 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1665 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2231  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1665 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n502 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2230  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4047 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1664 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2229  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1664 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n503 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2228  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4045 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1653 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2227  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1653 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n513 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2226  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4058 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1644 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2225  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1644 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n522 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2224  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4058 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1643 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2223  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1643 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n523 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2222  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4058 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1642 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2221  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1642 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n524 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2220  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4058 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1641 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2219  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1641 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n525 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2218  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4057 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1640 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2217  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1640 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n526 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2216  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4057 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1639 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2215  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1639 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n527 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2214  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4057 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1638 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2213  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1638 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n528 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2212  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4057 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1637 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2211  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1637 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n529 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2210  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4057 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1636 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2209  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1636 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n530 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2208  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4056 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1635 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2207  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1635 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n531 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2206  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4056 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1634 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2205  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1634 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n532 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2204  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4056 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1633 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2203  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1633 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n533 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2202  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4056 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1632 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2201  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1632 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n534 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2200  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4056 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1631 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2199  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1631 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n535 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2198  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4055 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1630 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2197  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1630 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n536 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2196  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4055 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1629 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2195  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1629 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n537 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2194  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4055 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1628 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2193  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1628 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n538 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2192  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4055 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1627 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2191  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1627 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n539 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2190  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4055 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1626 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2189  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1626 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n540 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2188  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4054 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1625 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2187  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1625 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n541 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2186  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4054 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1624 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2185  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1624 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n542 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2184  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4054 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1623 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2183  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1623 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n543 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2182  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4054 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1622 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2181  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1622 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n544 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2180  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4054 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1620 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2179  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1620 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n545 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2178  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4067 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1611 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2177  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1611 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n554 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2176  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4067 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1610 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2175  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1610 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n555 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2174  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4067 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1609 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2173  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1609 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n556 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2172  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4067 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1608 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2171  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1608 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n557 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2170  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4066 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1607 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2169  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1607 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n558 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2168  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4066 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1606 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2167  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1606 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n559 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2166  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4066 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1605 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2165  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1605 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n560 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2164  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4066 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1604 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2163  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1604 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n561 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2162  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4066 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1603 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2161  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1603 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n562 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2160  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4065 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1602 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2159  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1602 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n563 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2158  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4065 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1601 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2157  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1601 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n564 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2156  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4065 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1600 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2155  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1600 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n565 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2154  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4065 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1599 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2153  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1599 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n566 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2152  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4065 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1598 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2151  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1598 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n567 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2150  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4064 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1597 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2149  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1597 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n568 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2148  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4064 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1596 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2147  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1596 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n569 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2146  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4064 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1595 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2145  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1595 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n570 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2144  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4064 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1594 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2143  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1594 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n571 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2142  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4064 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1593 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2141  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1593 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n572 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2140  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4063 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1592 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2139  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1592 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n573 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2138  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4063 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1591 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2137  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1591 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n574 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2136  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4063 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1590 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2135  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1590 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n575 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2134  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4063 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1589 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2133  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1589 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n576 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2132  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4063 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1587 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2131  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1587 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n577 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2130  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4096 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1584 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2129  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1584 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n642 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2128  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4096 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1583 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2127  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1583 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n643 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2126  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4095 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1582 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2125  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1582 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n644 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2124  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4095 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1581 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2123  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1581 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n645 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2122  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4095 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1580 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2121  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1580 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n646 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2120  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4095 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1579 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2119  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1579 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n647 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2118  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4095 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1578 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2117  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1578 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n648 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2116  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4094 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1577 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2115  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1577 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n649 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2114  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4093 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1571 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2113  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1571 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n655 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2112  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4093 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1570 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2111  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1570 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n656 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2110  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4093 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1569 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2109  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1569 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n657 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2108  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4093 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1568 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2107  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1568 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n658 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2106  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4092 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1567 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2105  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1567 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n659 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2104  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4092 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1566 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2103  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1566 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n660 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2102  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4092 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1565 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2101  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1565 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n661 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2100  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4092 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1564 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2099  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1564 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n662 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2098  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4092 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1563 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2097  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1563 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n663 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2096  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4090 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1552 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2095  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1552 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n673 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2094  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4105 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1551 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2093  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1551 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n674 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2092  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4105 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1550 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2091  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1550 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n675 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2090  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4104 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1549 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2089  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1549 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n676 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2088  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4104 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1548 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2087  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1548 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n677 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2086  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4104 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1547 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2085  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1547 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n678 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2084  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4104 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1546 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2083  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1546 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n679 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2082  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4104 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1545 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2081  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1545 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n680 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2080  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4103 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1544 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2079  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1544 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n681 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2078  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4102 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1538 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2077  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1538 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n687 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2076  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4102 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1537 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2075  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1537 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n688 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2074  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4102 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1536 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2073  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1536 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n689 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2072  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4102 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1535 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2071  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1535 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n690 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2070  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4101 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1534 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2069  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1534 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n691 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2068  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4101 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1533 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2067  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n692 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2066  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4101 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1532 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2065  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n693 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2064  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4101 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1531 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2063  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1531 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n694 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2062  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4101 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1530 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2061  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n695 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2060  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4099 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1519 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2059  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1519 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n705 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2058  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4130 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1507 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2057  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1507 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n778 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2056  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4130 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1506 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2055  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1506 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n779 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2054  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4130 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1505 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2053  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1505 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n780 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2052  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4130 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1504 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2051  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1504 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n781 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2050  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4129 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1503 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2049  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1503 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n782 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2048  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4129 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1502 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2047  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1502 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n783 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2046  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4129 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1501 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2045  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1501 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n784 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2044  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4129 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1500 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2043  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1500 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n785 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2042  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4129 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1499 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2041  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1499 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n786 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2040  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4128 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1498 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2039  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1498 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n787 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2038  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4128 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1497 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2037  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1497 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n788 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2036  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4128 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1496 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2035  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1496 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n789 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2034  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4128 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1495 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2033  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1495 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n790 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2032  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4128 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1494 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2031  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1494 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n791 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2030  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4127 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1493 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2029  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1493 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n792 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2028  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4127 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1492 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2027  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1492 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n793 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2026  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4127 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1491 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2025  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1491 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n794 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2024  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4127 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1490 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2023  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1490 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n795 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2022  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4127 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1489 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2021  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1489 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n796 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2020  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4126 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1488 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2019  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1488 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n797 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2018  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4126 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1487 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2017  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1487 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n798 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2016  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4126 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1486 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2015  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1486 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n799 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2014  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4126 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1485 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2013  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1485 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n800 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2012  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4126 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1483 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2011  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1483 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n801 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2010  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4139 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1474 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2009  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1474 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n810 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2008  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4139 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1473 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2007  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1473 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n811 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2006  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4139 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1472 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2005  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1472 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n812 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2004  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4139 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1471 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2003  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1471 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n813 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2002  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4138 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1470 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2001  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1470 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n814 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2000  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4138 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1469 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1999  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1469 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n815 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1998  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4138 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1468 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1997  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1468 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n816 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1996  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4138 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1467 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1995  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1467 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n817 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1994  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4138 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1466 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1993  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1466 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n818 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1992  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4137 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1465 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1991  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1465 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n819 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1990  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4137 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1464 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1989  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1464 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n820 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1988  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4137 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1463 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1987  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1463 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n821 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1986  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4137 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1462 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1985  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1462 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n822 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1984  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4137 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1461 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1983  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1461 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n823 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1982  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4136 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1460 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1981  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1460 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n824 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1980  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4136 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1459 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1979  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1459 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n825 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1978  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4136 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1458 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1977  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1458 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n826 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1976  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4136 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1457 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1975  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1457 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n827 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1974  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4136 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1456 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1973  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1456 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n828 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1972  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4135 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1455 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1971  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1455 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n829 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1970  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4135 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1454 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1969  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1454 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n830 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1968  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4135 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1453 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1967  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1453 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n831 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1966  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4135 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1452 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1965  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1452 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n832 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1964  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4135 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1450 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1963  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1450 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n833 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1962  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4148 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1441 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1961  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1441 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n842 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1960  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4148 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1440 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1959  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1440 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n843 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1958  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4148 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1439 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1957  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1439 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n844 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1956  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4148 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1438 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1955  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1438 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n845 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1954  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4147 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1437 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1953  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1437 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n846 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1952  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4147 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1436 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1951  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1436 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n847 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1950  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4147 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1435 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1949  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1435 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n848 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1948  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4147 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1434 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1947  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1434 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n849 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1946  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4147 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1433 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1945  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1433 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n850 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1944  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4146 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1432 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1943  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1432 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n851 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1942  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4146 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1431 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1941  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1431 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n852 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1940  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4146 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1430 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1939  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1430 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n853 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1938  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4146 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1429 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1937  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1429 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n854 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1936  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4146 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1428 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1935  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1428 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n855 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1934  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4145 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1427 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1933  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1427 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n856 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1932  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4145 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1426 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1931  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1426 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n857 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1930  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4145 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1425 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1929  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1425 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n858 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1928  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4145 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1424 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1927  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1424 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n859 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1926  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4145 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1423 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1925  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1423 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n860 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1924  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4144 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1422 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1923  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1422 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n861 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1922  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4144 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1421 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1921  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1421 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n862 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1920  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4144 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1420 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1919  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1420 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n863 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1918  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4144 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1419 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1917  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1419 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n864 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1916  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4144 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1417 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1915  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1417 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n865 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1914  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4157 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1408 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1913  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1408 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n874 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1912  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4157 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1407 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1911  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1407 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n875 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1910  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4157 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1406 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1909  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1406 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n876 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1908  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4157 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1405 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1907  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1405 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n877 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1906  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4156 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1404 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1905  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1404 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n878 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1904  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4156 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1403 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1903  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1403 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n879 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1902  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4156 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1402 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1901  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1402 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n880 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1900  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4156 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1401 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1899  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1401 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n881 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1898  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4156 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1400 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1897  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1400 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n882 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1896  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4155 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1399 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1895  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1399 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n883 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1894  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4155 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1398 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1893  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1398 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n884 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1892  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4155 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1397 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1891  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1397 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n885 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1890  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4155 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1396 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1889  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1396 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n886 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1888  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4155 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1395 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1887  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1395 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n887 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1886  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4154 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1394 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1885  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1394 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n888 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1884  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4154 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1393 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1883  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1393 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n889 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1882  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4154 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1392 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1881  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1392 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n890 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1880  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4154 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1391 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1879  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1391 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n891 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1878  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4154 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1390 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1877  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1390 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n892 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1876  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4153 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1389 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1875  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1389 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n893 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1874  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4153 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1388 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1873  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1388 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n894 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1872  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4153 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1387 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1871  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1387 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n895 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1870  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4153 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1386 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1869  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1386 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n896 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1868  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4153 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1384 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1867  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1384 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n897 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1866  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4168 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1382 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1865  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1382 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n898 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1864  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4168 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1381 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1863  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1381 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n899 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1862  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4167 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1380 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1861  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1380 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n900 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1860  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4167 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1379 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1859  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1379 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n901 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1858  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4167 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1378 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1857  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1378 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n902 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1856  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4167 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1377 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1855  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1377 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n903 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1854  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4167 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1376 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1853  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1376 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n904 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1852  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4166 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1375 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1851  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1375 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n905 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1850  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4166 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1374 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1849  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1374 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n906 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1848  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4166 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1373 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1847  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1373 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n907 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1846  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4166 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1372 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1845  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1372 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n908 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1844  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4166 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1371 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1843  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1371 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n909 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1842  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4165 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1370 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1841  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1370 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n910 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1840  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4165 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1369 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1839  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1369 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n911 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1838  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4165 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1368 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1837  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1368 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n912 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1836  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4165 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1367 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1835  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1367 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n913 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1834  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4165 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1366 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1833  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1366 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n914 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1832  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4164 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1365 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1831  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1365 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n915 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1830  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4164 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1364 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1829  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1364 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n916 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1828  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4164 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1363 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1827  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1363 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n917 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1826  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4164 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1362 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1825  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1362 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n918 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1824  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4164 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1361 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1823  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1361 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n919 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1822  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4163 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1360 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1821  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1360 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n920 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1820  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4163 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1359 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1819  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1359 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n921 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1818  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4163 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1358 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1817  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1358 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n922 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1816  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4163 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1357 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1815  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1357 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n923 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1814  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4163 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1356 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1813  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1356 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n924 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1812  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4162 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1355 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1811  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1355 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n925 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1810  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4162 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1354 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1809  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1354 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n926 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1808  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4162 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1353 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1807  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1353 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n927 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1806  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4162 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1352 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1805  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1352 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n928 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1804  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4162 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1350 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1803  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1350 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n929 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1802  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4211 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1330 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1801  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1330 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1066 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1800  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4211 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1329 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1799  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1329 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1067 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1798  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4211 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1328 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1797  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1328 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1068 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1796  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4211 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1327 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1795  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1327 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1069 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1794  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4210 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1326 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1793  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1326 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1070 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1792  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4210 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1325 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1791  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1325 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1071 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1790  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4210 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1324 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1789  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1324 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1072 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1788  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4210 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1323 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1787  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1323 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1073 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1786  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4210 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1322 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1785  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1322 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1074 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1784  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4209 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1321 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1783  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1321 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1075 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1782  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4209 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1320 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1781  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1320 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1076 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1780  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4209 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1319 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1779  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1319 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1077 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1778  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4209 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1318 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1777  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1318 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1078 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1776  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4209 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1317 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1775  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1317 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1079 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1774  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4208 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1316 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1773  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1316 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1080 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1772  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4208 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1315 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1771  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1315 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1081 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1770  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4208 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1314 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1769  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1314 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1082 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1768  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4208 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1313 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1767  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1313 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1083 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1766  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4208 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1312 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1765  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1312 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1084 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1764  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4207 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1311 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1763  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1311 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1085 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1762  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4207 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1310 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1761  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1310 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1086 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1760  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4207 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1309 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1759  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1309 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1087 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1758  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4207 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1308 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1757  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1308 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1088 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1756  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4207 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1306 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1755  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1306 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1089 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1754  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4220 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1296 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1753  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1296 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1098 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1752  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4220 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1295 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1751  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1295 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1099 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1750  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4220 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1294 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1749  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1294 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1100 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1748  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4220 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1293 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1747  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1293 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1101 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1746  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4219 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1292 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1745  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1292 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1102 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1744  ( .A1(\dp/n4 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4219 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1291 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1743  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1291 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1103 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1742  ( .A1(
        \dp/wr_data_id_i [17]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4219 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1290 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1741  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1290 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1104 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1740  ( .A1(
        \dp/wr_data_id_i [16]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4219 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1289 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1739  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1289 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1105 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1738  ( .A1(
        \dp/wr_data_id_i [15]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4219 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1288 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1737  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1288 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1106 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1736  ( .A1(
        \dp/wr_data_id_i [14]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4218 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1287 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1735  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1287 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1107 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1734  ( .A1(
        \dp/wr_data_id_i [13]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4218 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1286 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1733  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1286 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1108 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1732  ( .A1(
        \dp/wr_data_id_i [12]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4218 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1285 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1731  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1285 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1109 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1730  ( .A1(
        \dp/wr_data_id_i [11]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4218 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1284 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1729  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1284 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1110 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1728  ( .A1(
        \dp/wr_data_id_i [10]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4218 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1283 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1727  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1283 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1111 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1726  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4217 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1282 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1725  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1282 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1112 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1724  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4217 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1281 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1723  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1281 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1113 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1722  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4217 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1280 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1721  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1280 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1114 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1720  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4217 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1279 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1719  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1279 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1115 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1718  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4217 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1278 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1717  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1278 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1116 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1716  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4216 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1277 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1715  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1277 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1117 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1714  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4216 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1276 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1713  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1276 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1118 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1712  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4216 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1275 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1711  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1275 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1119 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1710  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4216 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1274 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1709  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1274 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1120 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1708  ( .A1(
        \dp/wr_data_id_i [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4216 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1272 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1707  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1272 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1121 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1706  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_control_out ), .A2(
        \dp/id_stage/regfile/DataPath/mux_en_control_out ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1342 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1705  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3910 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3692 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1704  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3910 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3691 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1703  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3910 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3690 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1702  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3910 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n5 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3689 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1701  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3910 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n6 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3688 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1700  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3911 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n7 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3687 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1699  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3911 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3686 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1698  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3911 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n9 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3685 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1697  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3911 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n10 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3684 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1696  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3911 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n11 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3683 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1695  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3912 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n12 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3682 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1694  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3912 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n13 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3681 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1693  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3912 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n14 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3680 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1692  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3912 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n15 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3679 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1691  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3912 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n16 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3678 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1690  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3913 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n17 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3677 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1689  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3913 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n18 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3676 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1688  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3913 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n19 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3675 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1687  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3913 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n20 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3674 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1686  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3913 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n21 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3673 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1685  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3914 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n22 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3672 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1684  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3914 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n23 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3671 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1683  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3914 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n24 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3670 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1682  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3914 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n25 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3669 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1681  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3914 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n26 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3668 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1680  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3915 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n27 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3667 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1679  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3915 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n28 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3666 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1678  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3915 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n29 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3665 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1677  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3915 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n30 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3664 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1676  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3915 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n31 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3663 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1675  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3916 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n32 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3662 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1674  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3916 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n33 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3661 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1673  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3919 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n34 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3660 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1672  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3919 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n35 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3659 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1671  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3919 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n36 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3658 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1670  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3919 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n37 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3657 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1669  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3919 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n38 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3656 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1668  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3920 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n39 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3655 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1667  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3920 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n40 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3654 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1666  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3920 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n41 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3653 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1665  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3920 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n42 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3652 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1664  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3920 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n43 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3651 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1663  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3921 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n44 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3650 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1662  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3921 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n45 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3649 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1661  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3921 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n46 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3648 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1660  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3921 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n47 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3647 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1659  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3921 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n48 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3646 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1658  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3922 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n49 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3645 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1657  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3922 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n50 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3644 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1656  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3922 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n51 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3643 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1655  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3922 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n52 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3642 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1654  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3922 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n53 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3641 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1653  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3923 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n54 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3640 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1652  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3923 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n55 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3639 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1651  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3923 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n56 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3638 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1650  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3923 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n57 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3637 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1649  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3923 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n58 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3636 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1648  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3924 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n59 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3635 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1647  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3924 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n60 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3634 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1646  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3924 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n61 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3633 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1645  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3924 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n62 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3632 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1644  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3924 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n63 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3631 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1643  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3925 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n64 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3630 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1642  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3925 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n65 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3629 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1641  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3946 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n130 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3628 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1640  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3946 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n131 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3627 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1639  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3946 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n132 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3626 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1638  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3946 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n133 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3625 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1637  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3946 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n134 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3624 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1636  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3947 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n135 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3623 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1635  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3947 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n136 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3622 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1634  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3947 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n137 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3621 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1633  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3947 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n138 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3620 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1632  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3947 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n139 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3619 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1631  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3948 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n140 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3618 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1630  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3948 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n141 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3617 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1629  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3948 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n142 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3616 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1628  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3948 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n143 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3615 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1627  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3948 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n144 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3614 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1626  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3949 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n145 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3613 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1625  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3949 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n146 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3612 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1624  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3949 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n147 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3611 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1623  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3949 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n148 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3610 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1622  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3949 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n149 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3609 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1621  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3950 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n150 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3608 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1620  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3950 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n151 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3607 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1619  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3950 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n152 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3606 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1618  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3950 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n153 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3605 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1617  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3950 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n154 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3604 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1616  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3951 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n155 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3603 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1615  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3951 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3602 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1614  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3951 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3601 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1613  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3951 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n158 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3600 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1612  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3951 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3599 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1611  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3952 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3598 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1610  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3952 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n161 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3597 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1609  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3955 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n162 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3596 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1608  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3955 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n163 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3595 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1607  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3955 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n164 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3594 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1606  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3955 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n165 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3593 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1605  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3955 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n166 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3592 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1604  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3956 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n167 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3591 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1603  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3956 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n168 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3590 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1602  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3956 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n169 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3589 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1601  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3956 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n170 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3588 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1600  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3956 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n171 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3587 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1599  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3957 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n172 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3586 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1598  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3957 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n173 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3585 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1597  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3957 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n174 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3584 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1596  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3957 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n175 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3583 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1595  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3957 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n176 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3582 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1594  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3958 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n177 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3581 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1593  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3958 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n178 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3580 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1592  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3958 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n179 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3579 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1591  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3958 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n180 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3578 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1590  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3958 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n181 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3577 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1589  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3959 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n182 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3576 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1588  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3959 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n183 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3575 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1587  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3959 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n184 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3574 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1586  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3959 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n185 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3573 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1585  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3959 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n186 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3572 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1584  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3960 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n187 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3571 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1583  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3960 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n188 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3570 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1582  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3960 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n189 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3569 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1581  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3960 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n190 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3568 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1580  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3960 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n191 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3567 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1579  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3961 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n192 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3566 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1578  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3961 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n193 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3565 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1577  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3991 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n290 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3564 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1576  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3991 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n291 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3563 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1575  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3991 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n292 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3562 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1574  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3991 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n293 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3561 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1573  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3991 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n294 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3560 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1572  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3992 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n295 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3559 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1571  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3992 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n296 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3558 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1570  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3992 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n297 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3557 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1569  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3992 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n298 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3556 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1568  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3992 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n299 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3555 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1567  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3993 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n300 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3554 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1566  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3993 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n301 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3553 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1565  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3993 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n302 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3552 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1564  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3993 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n303 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3551 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1563  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3993 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n304 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3550 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1562  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3994 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n305 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3549 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1561  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3994 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n306 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3548 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1560  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3994 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n307 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3547 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1559  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3994 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n308 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3546 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1558  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3994 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n309 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3545 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1557  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3995 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n310 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3544 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1556  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3995 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n311 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3543 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1555  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3995 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n312 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3542 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1554  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3995 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n313 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3541 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1553  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3995 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n314 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3540 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1552  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3996 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n315 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3539 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1551  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3996 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n316 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3538 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1550  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3996 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n317 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3537 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1549  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3996 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n318 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3536 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1548  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3996 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n319 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3535 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1547  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3997 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n320 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3534 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1546  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3997 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n321 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3533 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1545  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4000 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n322 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3532 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1544  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4000 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n323 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3531 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1543  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4000 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n324 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3530 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1542  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4000 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n325 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3529 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1541  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4000 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n326 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3528 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1540  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4001 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n327 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3527 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1539  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4001 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n328 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3526 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1538  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4001 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n329 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3525 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1537  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4001 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n330 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3524 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1536  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4001 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n331 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3523 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1535  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4002 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n332 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3522 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1534  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4002 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n333 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3521 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1533  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4002 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n334 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3520 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1532  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4002 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n335 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3519 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1531  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4002 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n336 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3518 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1530  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4003 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n337 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3517 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1529  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4003 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n338 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3516 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1528  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4003 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n339 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3515 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1527  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4003 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n340 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3514 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1526  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4003 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n341 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3513 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1525  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4004 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n342 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3512 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1524  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4004 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n343 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3511 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1523  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4004 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n344 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3510 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1522  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4004 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n345 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3509 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1521  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4004 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n346 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3508 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1520  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4005 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n347 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3507 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1519  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4005 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n348 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3506 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1518  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4005 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n349 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3505 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1517  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4005 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n350 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3504 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1516  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4005 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n351 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3503 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1515  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4006 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n352 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3502 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1514  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4006 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n353 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3501 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1513  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4027 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n418 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3500 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1512  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4027 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n419 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3499 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1511  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4027 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n420 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3498 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1510  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4027 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n421 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3497 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1509  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4027 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n422 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3496 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1508  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4028 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n423 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3495 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1507  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4028 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n424 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3494 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1506  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4028 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n425 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3493 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1505  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4028 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n426 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3492 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1504  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4028 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n427 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3491 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1503  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4029 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n428 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3490 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1502  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4029 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n429 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3489 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1501  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4029 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n430 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3488 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1500  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4029 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n431 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3487 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1499  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4029 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n432 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3486 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1498  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4030 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n433 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3485 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1497  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4030 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n434 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3484 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1496  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4030 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n435 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3483 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1495  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4030 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n436 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3482 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1494  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4030 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n437 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3481 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1493  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4031 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n438 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3480 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1492  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4031 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n439 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3479 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1491  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4031 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n440 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3478 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1490  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4031 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n441 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3477 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1489  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4031 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n442 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3476 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1488  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4032 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n443 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3475 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1487  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4032 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n444 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3474 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1486  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4032 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n445 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3473 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1485  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4032 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n446 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3472 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1484  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4032 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n447 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3471 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1483  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4033 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n448 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3470 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1482  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4033 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n449 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3469 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1481  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4036 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n450 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3468 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1480  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4036 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n451 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3467 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1479  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4036 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n452 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3466 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1478  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4036 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n453 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3465 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1477  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4036 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n454 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3464 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1476  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4037 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n455 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3463 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1475  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4037 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n456 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3462 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1474  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4037 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n457 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3461 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1473  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4037 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n458 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3460 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1472  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4037 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n459 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3459 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1471  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4038 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n460 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3458 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1470  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4038 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n461 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3457 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1469  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4038 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n462 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3456 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1468  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4038 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n463 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3455 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1467  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4038 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n464 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3454 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1466  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4039 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n465 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3453 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1465  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4039 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n466 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3452 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1464  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4039 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n467 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3451 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1463  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4039 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n468 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3450 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1462  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4039 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n469 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3449 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1461  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4040 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n470 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3448 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1460  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4040 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n471 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3447 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1459  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4040 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n472 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3446 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1458  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4040 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n473 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3445 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1457  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4040 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n474 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3444 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1456  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4041 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n475 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3443 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1455  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4041 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n476 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3442 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1454  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4041 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n477 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3441 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1453  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4041 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n478 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3440 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1452  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4041 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n479 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3439 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1451  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4042 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n480 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3438 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1450  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4042 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n481 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3437 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1449  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4072 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n578 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3436 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1448  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4072 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n579 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3435 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1447  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4072 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n580 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3434 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1446  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4072 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n581 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3433 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1445  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4072 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n582 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3432 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1444  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4073 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n583 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3431 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1443  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4073 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n584 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3430 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1442  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4073 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n585 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3429 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1441  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4073 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n586 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3428 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1440  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4073 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n587 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3427 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1439  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4074 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n588 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3426 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1438  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4074 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n589 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3425 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1437  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4074 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n590 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3424 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1436  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4074 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n591 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3423 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1435  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4074 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n592 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3422 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1434  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4075 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n593 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3421 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1433  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4075 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n594 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3420 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1432  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4075 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n595 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3419 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1431  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4075 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n596 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3418 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1430  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4075 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n597 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3417 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1429  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4076 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n598 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3416 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1428  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4076 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n599 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3415 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1427  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4076 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n600 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3414 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1426  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4076 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n601 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3413 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1425  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4076 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n602 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3412 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1424  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4077 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n603 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3411 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1423  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4077 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n604 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3410 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1422  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4077 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n605 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3409 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1421  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4077 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n606 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3408 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1420  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4077 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n607 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3407 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1419  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4078 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n608 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3406 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1418  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4078 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n609 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3405 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1417  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4081 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n610 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3404 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1416  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4081 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n611 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3403 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1415  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4081 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n612 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3402 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1414  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4081 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n613 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3401 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1413  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4081 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n614 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3400 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1412  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4082 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n615 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3399 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1411  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4082 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n616 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3398 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1410  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4082 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n617 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3397 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1409  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4082 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n618 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3396 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1408  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4082 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n619 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3395 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1407  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4083 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n620 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3394 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1406  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4083 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n621 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3393 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1405  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4083 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n622 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3392 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1404  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4083 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n623 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3391 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1403  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4083 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n624 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3390 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1402  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4084 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n625 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3389 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1401  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4084 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n626 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3388 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1400  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4084 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n627 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3387 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1399  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4084 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n628 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3386 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1398  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4084 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n629 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3385 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1397  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4085 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n630 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3384 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1396  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4085 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n631 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3383 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1395  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4085 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n632 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3382 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1394  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4085 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n633 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3381 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1393  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4085 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n634 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3380 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1392  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4086 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n635 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3379 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1391  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4086 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n636 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3378 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1390  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4086 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n637 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3377 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1389  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4086 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n638 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3376 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1388  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4086 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n639 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3375 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1387  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4087 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n640 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3374 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1386  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4087 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n641 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3373 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1385  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4108 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n706 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3372 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1384  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4108 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n707 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3371 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1383  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4108 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n708 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3370 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1382  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4108 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n709 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3369 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1381  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4108 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n710 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3368 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1380  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4109 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n711 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3367 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1379  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4109 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n712 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3366 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1378  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4109 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n713 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3365 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1377  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4109 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n714 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3364 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1376  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4109 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n715 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3363 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1375  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4110 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n716 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3362 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1374  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4110 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n717 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3361 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1373  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4110 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n718 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3360 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1372  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4110 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n719 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3359 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1371  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4110 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n720 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3358 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1370  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4111 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n721 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3357 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1369  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4111 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n722 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3356 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1368  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4111 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n723 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3355 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1367  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4111 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n724 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3354 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1366  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4111 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n725 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3353 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1365  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4112 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n726 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3352 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1364  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4112 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n727 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3351 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1363  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4112 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n728 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3350 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1362  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4112 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n729 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3349 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1361  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4112 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n730 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3348 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1360  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4113 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n731 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3347 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1359  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4113 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n732 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3346 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1358  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4113 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n733 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3345 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1357  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4113 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n734 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3344 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1356  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4113 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n735 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3343 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1355  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4114 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n736 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3342 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1354  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4114 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n737 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3341 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1353  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4117 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n738 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3340 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1352  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4117 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n739 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3339 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1351  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4117 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n740 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3338 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1350  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4117 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n741 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3337 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1349  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4117 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n742 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3336 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1348  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4118 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n743 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3335 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1347  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4118 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n744 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3334 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1346  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4118 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n745 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3333 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1345  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4118 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n746 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3332 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1344  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4118 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n747 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3331 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1343  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4119 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n748 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3330 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1342  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4119 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n749 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3329 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1341  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4119 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n750 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3328 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1340  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4119 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n751 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3327 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1339  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4119 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n752 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3326 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1338  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4120 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n753 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3325 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1337  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4120 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n754 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3324 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1336  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4120 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n755 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3323 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1335  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4120 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n756 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3322 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1334  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4120 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n757 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3321 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1333  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4121 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n758 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3320 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1332  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4121 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n759 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3319 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1331  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4121 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n760 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3318 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1330  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4121 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n761 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3317 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1329  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4121 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n762 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3316 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1328  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4122 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n763 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3315 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1327  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4122 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n764 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3314 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1326  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4122 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n765 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3313 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1325  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4122 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n766 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3312 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1324  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4122 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n767 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3311 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1323  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4123 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n768 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3310 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1322  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4123 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n769 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3309 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1321  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4171 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n930 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3308 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1320  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4171 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n931 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3307 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1319  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4171 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n932 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3306 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1318  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4171 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n933 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3305 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1317  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4171 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n934 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3304 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1316  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4172 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n935 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3303 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1315  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4172 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n936 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3302 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1314  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4172 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n937 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3301 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1313  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4172 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n938 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3300 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1312  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4172 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n939 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3299 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1311  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4173 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n940 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3298 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1310  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4173 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n941 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3297 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1309  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4173 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n942 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3296 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1308  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4173 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n943 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3295 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1307  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4173 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n944 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3294 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1306  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4174 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n945 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3293 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1305  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4174 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n946 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3292 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1304  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4174 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n947 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3291 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1303  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4174 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n948 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3290 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1302  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4174 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n949 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3289 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1301  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4175 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n950 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3288 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1300  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4175 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n951 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3287 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1299  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4175 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n952 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3286 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1298  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4175 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n953 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3285 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1297  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4175 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n954 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3284 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1296  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4176 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n955 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3283 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1295  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4176 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n956 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3282 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1294  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4176 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n957 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3281 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1293  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4176 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n958 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3280 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1292  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4176 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n959 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3279 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1291  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4177 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n960 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3278 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1290  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4177 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n961 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3277 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1289  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4180 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n962 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3276 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1288  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4180 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n963 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3275 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1287  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4180 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n964 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3274 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1286  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4180 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n965 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3273 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1285  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4180 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n966 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3272 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1284  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4181 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n967 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3271 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1283  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4181 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n968 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3270 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1282  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4181 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n969 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3269 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1281  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4181 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n970 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3268 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1280  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4181 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n971 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3267 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1279  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4182 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n972 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3266 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1278  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4182 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n973 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3265 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1277  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4182 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n974 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3264 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1276  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4182 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n975 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3263 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1275  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4182 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n976 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3262 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1274  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4183 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n977 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3261 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1273  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4183 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n978 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3260 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1272  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4183 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n979 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3259 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1271  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4183 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n980 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3258 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1270  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4183 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n981 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3257 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1269  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4184 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n982 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3256 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1268  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4184 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n983 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3255 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1267  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4184 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n984 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3254 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1266  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4184 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n985 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3253 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1265  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4184 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n986 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3252 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1264  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4185 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n987 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3251 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1263  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4185 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n988 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3250 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1262  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4185 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n989 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3249 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1261  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4185 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n990 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3248 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1260  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4185 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n991 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3247 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1259  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4186 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n992 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3246 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1258  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4186 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n993 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3245 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1257  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4189 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n994 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3244 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1256  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4189 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n995 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3243 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1255  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4189 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n996 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3242 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1254  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4189 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n997 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3241 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1253  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4189 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n998 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3240 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1252  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4190 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n999 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3239 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1251  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4190 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1000 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3238 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1250  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4190 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1001 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3237 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1249  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4190 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1002 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3236 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1248  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4190 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1003 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3235 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1247  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4191 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1004 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3234 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1246  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4191 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1005 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3233 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1245  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4191 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1006 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3232 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1244  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4191 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1007 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3231 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1243  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4191 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1008 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3230 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1242  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4192 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1009 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3229 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1241  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4192 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1010 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3228 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1240  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4192 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1011 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3227 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1239  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4192 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1012 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3226 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1238  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4192 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1013 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3225 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1237  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4193 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1014 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3224 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1236  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4193 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1015 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3223 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1235  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4193 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1016 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3222 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1234  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4193 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1017 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3221 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1233  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4193 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1018 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3220 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1232  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4194 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1019 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3219 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1231  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4194 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1020 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3218 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1230  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4194 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1021 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3217 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1229  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4194 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1022 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3216 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1228  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4194 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1023 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3215 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1227  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4195 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1024 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3214 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1226  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4195 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1025 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3213 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1225  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4198 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1026 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3212 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1224  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4198 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1027 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3211 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1223  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4198 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1028 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3210 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1222  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4198 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1029 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3209 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1221  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4198 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1030 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3208 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1220  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4199 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1031 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3207 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1219  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4199 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1032 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3206 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1218  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4199 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1033 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3205 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1217  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4199 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1034 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3204 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1216  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4199 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1035 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3203 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1215  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4200 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1036 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3202 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1214  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4200 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1037 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3201 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1213  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4200 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1038 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3200 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1212  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4200 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1039 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3199 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1211  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4200 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1040 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3198 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1210  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4201 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1041 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3197 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1209  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4201 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1042 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3196 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1208  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4201 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1043 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3195 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1207  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4201 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1044 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3194 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1206  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4201 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1045 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3193 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1205  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4202 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1046 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3192 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1204  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4202 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1047 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3191 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1203  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4202 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1048 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3190 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1202  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4202 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1049 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3189 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1201  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4202 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1050 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3188 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1200  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4203 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1051 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3187 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1199  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4203 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1052 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3186 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1198  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4203 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1053 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3185 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1197  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4203 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1054 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3184 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1196  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4203 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1055 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3183 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1195  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4204 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1056 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3182 ) );
  OAI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1194  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4204 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1057 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3181 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1193  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(\dp/n8 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4231 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1269 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1192  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1269 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1122 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1191  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [30]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4231 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1268 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1190  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1268 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1123 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1189  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [29]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4230 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1267 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1188  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1267 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1124 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1187  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [28]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4230 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1266 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1186  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1266 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1125 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1185  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(\dp/n6 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4230 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1265 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1184  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1265 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1126 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1183  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [26]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4230 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1264 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1182  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1264 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1127 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1181  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [25]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4230 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1263 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1180  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1263 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1128 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1179  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [24]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4229 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1262 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1178  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1262 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1129 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1177  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [23]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4229 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1261 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1176  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1261 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1130 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1175  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [22]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4229 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1260 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1174  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1260 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1131 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1173  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [21]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4229 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1259 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1172  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1259 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1132 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1171  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [20]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4229 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1258 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1170  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1258 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1133 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1169  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [19]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4228 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1257 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1168  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1257 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1134 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1167  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(\dp/n4 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4228 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][18] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1256 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1166  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1256 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1135 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1165  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [17]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4228 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][17] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1255 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1164  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1255 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1136 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1163  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [16]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4228 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][16] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1254 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1162  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1254 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1137 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1161  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [15]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4228 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][15] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1253 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1160  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1253 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1138 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1159  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [14]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4227 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][14] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1252 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1158  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1252 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1139 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1157  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [13]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4227 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][13] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1251 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1156  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1251 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1140 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1155  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [12]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4227 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][12] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1250 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1154  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1250 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1141 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1153  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ), .A2(
        \dp/wr_data_id_i [11]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4227 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][11] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1249 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1152  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1249 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1142 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1151  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [10]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4227 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][10] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1248 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1150  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1248 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1143 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1149  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [9]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4226 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1247 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1148  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1247 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1144 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1147  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [8]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4226 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1246 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1146  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1246 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1145 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1145  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [7]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4226 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1245 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1144  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1245 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1146 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1143  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [6]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4226 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1244 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1142  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1244 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1147 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1141  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [5]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4226 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1243 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1140  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1243 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1148 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1139  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [4]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4225 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1242 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1138  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1242 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1149 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1137  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [3]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4225 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1241 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1136  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1241 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1150 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1135  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [2]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4225 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1240 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1134  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1240 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1151 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1133  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [1]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4225 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1239 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1132  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1239 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1152 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1131  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ), .A2(
        \dp/wr_data_id_i [0]), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4225 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][0] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1237 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1130  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1237 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1153 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1129  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3934 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1924 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1128  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1924 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n66 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1127  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3934 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1923 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1126  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1923 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n67 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1125  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3933 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1922 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1124  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1922 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n68 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1123  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3933 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1921 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1122  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1921 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n69 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1121  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3933 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1920 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1120  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1920 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n70 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1119  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3933 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1919 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1118  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1919 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n71 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1117  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3933 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1918 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1116  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1918 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n72 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1115  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3932 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1917 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1114  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1917 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n73 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1113  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3943 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1891 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1112  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1891 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n98 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1111  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3943 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1890 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1110  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1890 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n99 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1109  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3942 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1889 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1108  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1889 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n100 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1107  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3942 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1888 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1106  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1888 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n101 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1105  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3942 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1887 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1104  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1887 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n102 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1103  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3942 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1886 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1102  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1886 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n103 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1101  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3942 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1885 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1100  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1885 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n104 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1099  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3941 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1884 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1098  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1884 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n105 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1097  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3970 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1856 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1096  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1856 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n194 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1095  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3970 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1855 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1094  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1855 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n195 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1093  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3969 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1854 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1092  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1854 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n196 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1091  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3969 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1853 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1090  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1853 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n197 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1089  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3969 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1852 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1088  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1852 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n198 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1087  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3969 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1851 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1086  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1851 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n199 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1085  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3969 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1850 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1084  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1850 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n200 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1083  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3968 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1849 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1082  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1849 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n201 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1081  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3979 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1822 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1080  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1822 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n226 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1079  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3979 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1821 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1078  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1821 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n227 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1077  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3978 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1820 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1076  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1820 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n228 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1075  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3978 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1819 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1074  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1819 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n229 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1073  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3978 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1818 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1072  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1818 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n230 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1071  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3978 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1817 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1070  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1817 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n231 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1069  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3978 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1816 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1068  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1816 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n232 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1067  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3977 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1815 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1066  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1815 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n233 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1065  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3988 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1789 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1064  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1789 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n258 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1063  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3988 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1788 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1062  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1788 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n259 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1061  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3987 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1787 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1060  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1787 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n260 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1059  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3987 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1786 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1058  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1786 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n261 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1057  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3987 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1785 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1056  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1785 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n262 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1055  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3987 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1784 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1054  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1784 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n263 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1053  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3987 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1783 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1052  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1783 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n264 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1051  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3986 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1782 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1050  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1782 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n265 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1049  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4015 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1754 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1048  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1754 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n354 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1047  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4015 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1753 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1046  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1753 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n355 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1045  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4014 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1752 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1044  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1752 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n356 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1043  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4014 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1751 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1042  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1751 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n357 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1041  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4014 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1750 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1040  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1750 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n358 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1039  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4014 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1749 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1038  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1749 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n359 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1037  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4014 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1748 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1036  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1748 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n360 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1035  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4013 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1747 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1034  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1747 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n361 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1033  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4024 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1721 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1032  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1721 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n386 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1031  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4024 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1720 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1030  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1720 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n387 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1029  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4023 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1719 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1028  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1719 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n388 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1027  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4023 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1718 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1026  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1718 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n389 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1025  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4023 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1717 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1024  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1717 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n390 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1023  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4023 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1716 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1022  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1716 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n391 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1021  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4023 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1715 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1020  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1715 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n392 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1019  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4022 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1714 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1018  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1714 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n393 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1017  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4022 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1713 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1016  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1713 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n394 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1015  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4022 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1712 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1014  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1712 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n395 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1013  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4022 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1711 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1012  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1711 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n396 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1011  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4022 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1710 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1010  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1710 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n397 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1009  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4021 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1709 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1008  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1709 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n398 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1007  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4019 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1699 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1006  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1699 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n408 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1005  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4019 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1698 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1004  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1698 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n409 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1003  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4019 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1697 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1002  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1697 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n410 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1001  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4019 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1696 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U1000  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1696 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n411 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U999  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4019 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1695 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U998  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1695 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n412 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U997  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4018 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1694 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U996  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1694 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n413 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U995  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4018 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1693 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U994  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1693 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n414 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U993  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4018 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1692 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U992  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1692 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n415 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U991  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4018 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1691 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U990  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1691 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n416 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U989  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4051 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1685 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U988  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1685 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n482 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U987  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4051 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1684 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U986  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1684 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n483 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U985  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4050 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1683 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U984  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1683 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n484 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U983  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4050 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1682 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U982  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1682 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n485 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U981  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4050 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1681 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U980  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1681 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n486 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U979  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4050 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1680 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U978  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1680 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n487 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U977  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4050 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1679 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U976  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1679 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n488 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U975  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4049 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1678 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U974  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1678 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n489 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U973  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4049 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1677 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U972  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1677 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n490 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U971  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4049 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1676 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U970  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1676 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n491 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U969  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4049 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1675 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U968  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1675 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n492 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U967  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4049 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1674 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U966  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1674 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n493 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U965  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4048 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1673 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U964  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1673 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n494 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U963  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4046 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1663 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U962  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1663 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n504 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U961  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4046 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1662 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U960  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1662 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n505 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U959  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4046 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1661 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U958  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1661 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n506 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U957  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4046 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1660 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U956  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1660 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n507 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U955  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4046 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1659 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U954  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1659 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n508 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U953  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4045 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1658 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U952  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1658 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n509 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U951  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4045 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1657 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U950  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1657 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n510 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U949  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4045 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1656 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U948  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1656 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n511 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U947  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4045 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1655 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U946  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1655 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n512 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U945  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4060 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1652 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U944  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1652 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n514 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U943  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4060 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1651 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U942  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1651 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n515 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U941  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4059 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1650 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U940  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1650 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n516 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U939  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4059 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1649 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U938  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1649 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n517 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U937  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4059 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1648 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U936  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1648 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n518 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U935  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4059 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1647 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U934  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1647 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n519 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U933  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4059 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1646 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U932  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1646 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n520 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U931  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4058 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1645 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U930  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1645 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n521 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U929  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4069 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1619 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U928  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1619 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n546 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U927  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4069 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1618 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U926  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1618 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n547 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U925  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4068 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1617 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U924  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1617 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n548 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U923  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4068 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1616 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U922  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1616 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n549 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U921  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4068 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1615 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U920  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1615 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n550 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U919  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4068 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1614 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U918  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1614 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n551 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U917  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4068 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1613 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U916  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1613 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n552 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U915  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4067 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1612 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U914  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1612 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n553 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U913  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4094 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1576 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U912  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1576 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n650 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U911  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4094 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1575 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U910  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1575 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n651 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U909  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4094 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1574 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U908  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1574 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n652 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U907  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4094 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1573 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U906  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1573 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n653 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U905  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4093 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1572 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U904  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1572 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n654 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U903  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4091 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1562 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U902  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1562 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n664 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U901  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4091 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1561 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U900  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1561 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n665 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U899  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4091 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1560 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U898  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1560 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n666 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U897  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4091 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1559 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U896  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1559 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n667 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U895  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4091 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1558 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U894  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1558 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n668 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U893  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4090 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1557 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U892  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1557 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n669 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U891  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4090 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1556 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U890  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1556 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n670 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U889  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4090 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1555 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U888  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1555 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n671 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U887  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4090 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1554 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U886  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1554 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n672 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U885  ( .A1(
        \dp/wr_data_id_i [23]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4103 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][23] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1543 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U884  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1543 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n682 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U883  ( .A1(
        \dp/wr_data_id_i [22]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4103 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][22] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1542 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U882  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1542 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n683 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U881  ( .A1(
        \dp/wr_data_id_i [21]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4103 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][21] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1541 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U880  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1541 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n684 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U879  ( .A1(
        \dp/wr_data_id_i [20]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4103 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][20] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1540 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U878  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1540 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n685 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U877  ( .A1(
        \dp/wr_data_id_i [19]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4102 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][19] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1539 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U876  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1539 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n686 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U875  ( .A1(
        \dp/wr_data_id_i [9]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4100 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][9] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1529 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U874  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n696 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U873  ( .A1(
        \dp/wr_data_id_i [8]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4100 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][8] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1528 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U872  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1528 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n697 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U871  ( .A1(
        \dp/wr_data_id_i [7]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4100 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][7] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1527 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U870  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1527 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n698 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U869  ( .A1(
        \dp/wr_data_id_i [6]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4100 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][6] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1526 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U868  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1526 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n699 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U867  ( .A1(
        \dp/wr_data_id_i [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4100 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][5] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1525 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U866  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1525 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n700 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U865  ( .A1(
        \dp/wr_data_id_i [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4099 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][4] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1524 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U864  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1524 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n701 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U863  ( .A1(
        \dp/wr_data_id_i [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4099 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][3] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1523 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U862  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1523 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n702 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U861  ( .A1(
        \dp/wr_data_id_i [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4099 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][2] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1522 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U860  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1522 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n703 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U859  ( .A1(
        \dp/wr_data_id_i [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4099 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][1] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1521 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U858  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1521 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n704 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U857  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4132 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1515 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U856  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1515 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n770 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U855  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4132 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1514 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U854  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1514 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n771 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U853  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4131 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1513 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U852  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1513 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n772 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U851  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4131 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1512 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U850  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1512 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n773 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U849  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4131 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1511 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U848  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1511 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n774 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U847  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4131 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1510 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U846  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1510 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n775 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U845  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4131 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1509 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U844  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1509 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n776 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U843  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4130 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1508 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U842  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1508 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n777 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U841  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4141 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1482 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U840  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1482 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n802 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U839  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4141 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1481 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U838  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1481 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n803 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U837  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4140 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1480 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U836  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1480 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n804 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U835  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4140 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1479 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U834  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1479 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n805 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U833  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4140 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1478 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U832  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1478 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n806 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U831  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4140 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1477 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U830  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1477 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n807 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U829  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4140 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1476 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U828  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1476 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n808 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U827  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4139 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1475 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U826  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1475 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n809 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U825  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4150 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1449 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U824  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1449 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n834 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U823  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4150 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1448 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U822  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1448 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n835 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U821  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4149 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1447 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U820  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1447 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n836 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U819  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4149 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1446 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U818  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1446 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n837 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U817  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4149 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1445 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U816  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1445 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n838 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U815  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4149 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1444 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U814  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1444 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n839 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U813  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4149 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1443 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U812  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1443 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n840 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U811  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4148 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1442 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U810  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1442 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n841 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U809  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4159 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1416 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U808  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1416 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n866 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U807  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4159 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1415 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U806  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1415 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n867 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U805  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4158 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1414 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U804  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1414 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n868 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U803  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4158 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1413 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U802  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1413 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n869 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U801  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4158 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1412 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U800  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1412 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n870 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U799  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4158 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1411 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U798  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1411 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n871 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U797  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4158 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1410 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U796  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1410 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n872 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U795  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4157 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1409 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U794  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1409 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n873 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U793  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4213 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1338 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U792  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1338 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1058 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U791  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4213 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1337 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U790  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1337 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1059 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U789  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4212 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1336 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U788  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1336 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1060 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U787  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4212 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1335 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U786  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1335 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1061 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U785  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4212 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1334 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U784  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1334 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1062 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U783  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4212 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1333 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U782  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1333 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1063 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U781  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4212 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1332 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U780  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1332 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1064 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U779  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4211 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1331 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U778  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1331 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1065 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U777  ( .A1(\dp/n8 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4222 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][31] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1304 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U776  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1304 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1090 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U775  ( .A1(
        \dp/wr_data_id_i [30]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4222 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][30] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1303 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U774  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1303 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1091 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U773  ( .A1(
        \dp/wr_data_id_i [29]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4221 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][29] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1302 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U772  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1302 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1092 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U771  ( .A1(
        \dp/wr_data_id_i [28]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4221 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][28] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1301 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U770  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1301 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1093 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U769  ( .A1(\dp/n6 ), 
        .A2(\dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4221 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][27] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1300 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U768  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1300 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1094 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U767  ( .A1(
        \dp/wr_data_id_i [26]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4221 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][26] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1299 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U766  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1299 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1095 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U765  ( .A1(
        \dp/wr_data_id_i [25]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4221 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][25] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1298 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U764  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1298 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1096 ) );
  AOI22_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U763  ( .A1(
        \dp/wr_data_id_i [24]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ), .B1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4220 ), .B2(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][24] ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1297 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U762  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1297 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1097 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U761  ( .A(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [3]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1201 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U760  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4240 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [3]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2536 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U759  ( .A(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [0]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4276 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U758  ( .A(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [1]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4242 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U757  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [0]), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [1]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ) );
  NOR3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U756  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [3]), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [4]), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4241 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2548 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U755  ( .A(
        \dp/id_stage/regfile/DataPath/mux_wr_out [3]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1192 ) );
  AND4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U754  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1342 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1192 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1191 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1271 ) );
  AND4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U753  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [3]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1342 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1191 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1190 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ) );
  AND4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U752  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [4]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1342 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1192 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1190 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ) );
  AND4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U751  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1342 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1192 ), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1191 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1190 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ) );
  AND4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U750  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [4]), .A2(
        \dp/id_stage/regfile/DataPath/mux_wr_out [3]), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1342 ), .A4(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1190 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U749  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2531 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1980 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U748  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2551 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1973 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U747  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2549 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1968 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U746  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2539 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1947 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U745  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2535 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1941 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U744  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2528 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1937 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U743  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1953 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U742  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_rd_out [5]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2580 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U741  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2531 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1979 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U740  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2535 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1943 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U739  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2535 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1942 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U738  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2528 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1936 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U737  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1954 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U736  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1952 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U735  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2581 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U734  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2579 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U733  ( .A(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4240 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U732  ( .A(
        \dp/id_stage/regfile/DataPath/mux_rd_out [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1195 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U731  ( .A(
        \dp/id_stage/regfile/DataPath/mux_rd_out [3]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1196 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U730  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2548 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1969 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U729  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2548 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1967 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U728  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2546 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1963 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U727  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2546 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1962 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U726  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2551 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1975 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U725  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2549 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1970 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U724  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2539 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1944 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U723  ( .A(
        \dp/id_stage/regfile/DataPath/mux_rd_out [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1197 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U722  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1949 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U721  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2576 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U720  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2551 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1976 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U719  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2549 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1971 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U718  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2539 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1945 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U717  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2528 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1939 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U716  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2531 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1934 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U715  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2536 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4241 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2531 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U714  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3179 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3178 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U713  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3163 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3155 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U712  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2536 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2528 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U711  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1195 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [3]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3163 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U710  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1196 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3179 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U709  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1201 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2552 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U708  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4240 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1201 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2538 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U707  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_rd_out [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3165 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3166 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U706  ( .A(
        \dp/id_stage/regfile/DataPath/mux_rd_out [0]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1199 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U705  ( .A(
        \dp/id_stage/regfile/DataPath/mux_rd_out [1]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1198 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U704  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2548 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1964 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U703  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2548 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1965 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U702  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2546 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1959 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U701  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2546 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2529 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1960 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U700  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_rd_out [0]), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [1]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U699  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4242 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4276 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ) );
  NOR3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U698  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_rd_out [3]), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [4]), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1197 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3175 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U697  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1349 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U696  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1344 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U695  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1383 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U694  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1349 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U693  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1349 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U692  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1347 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U691  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1347 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U690  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1344 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U689  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1341 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U688  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1339 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U687  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1339 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U686  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1305 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U685  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1305 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U684  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1270 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U683  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1341 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1271 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U682  ( .A(
        \dp/id_stage/regfile/DataPath/mux_wr_out [0]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1194 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U681  ( .A(
        \dp/id_stage/regfile/DataPath/mux_wr_out [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1191 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U680  ( .A(
        \dp/id_stage/regfile/DataPath/mux_wr_out [1]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1193 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U679  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1347 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U678  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1344 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U677  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1383 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U676  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1344 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U675  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1383 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U674  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1349 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U673  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1383 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U672  ( .A(
        \dp/id_stage/regfile/DataPath/mux_wr_out [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1190 ) );
  AND3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U671  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [0]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1193 ), .A3(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1349 ) );
  AND3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U670  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [1]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1194 ), .A3(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1347 ) );
  AND3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U669  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [1]), .A2(
        \dp/id_stage/regfile/DataPath/mux_wr_out [0]), .A3(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1344 ) );
  AND3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U668  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1194 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1193 ), .A3(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1383 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U667  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1305 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U666  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1823 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1270 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U665  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1341 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U664  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1686 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1270 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U663  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1341 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U662  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1517 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1339 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U661  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1341 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U660  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1339 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U659  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1305 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U658  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1270 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U657  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1339 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1271 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U656  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1305 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1271 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U655  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1270 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1271 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U654  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1347 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1345 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U653  ( .A(\dp/n8 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4275 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U652  ( .A(
        \dp/wr_data_id_i [30]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4274 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U651  ( .A(
        \dp/wr_data_id_i [29]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4273 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U650  ( .A(
        \dp/wr_data_id_i [28]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4272 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U649  ( .A(\dp/n6 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4271 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U648  ( .A(
        \dp/wr_data_id_i [26]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4270 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U647  ( .A(
        \dp/wr_data_id_i [25]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4269 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U646  ( .A(
        \dp/wr_data_id_i [24]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4268 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U645  ( .A(
        \dp/wr_data_id_i [23]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4267 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U644  ( .A(
        \dp/wr_data_id_i [22]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4266 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U643  ( .A(
        \dp/wr_data_id_i [21]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4265 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U642  ( .A(
        \dp/wr_data_id_i [20]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4264 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U641  ( .A(
        \dp/wr_data_id_i [19]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4263 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U640  ( .A(\dp/n4 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4262 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U639  ( .A(
        \dp/wr_data_id_i [17]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4261 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U638  ( .A(
        \dp/wr_data_id_i [16]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4260 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U637  ( .A(
        \dp/wr_data_id_i [15]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4259 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U636  ( .A(
        \dp/wr_data_id_i [14]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4258 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U635  ( .A(
        \dp/wr_data_id_i [13]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4257 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U634  ( .A(
        \dp/wr_data_id_i [12]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4256 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U633  ( .A(
        \dp/wr_data_id_i [11]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4255 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U632  ( .A(
        \dp/wr_data_id_i [10]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4254 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U631  ( .A(
        \dp/wr_data_id_i [9]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4253 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U630  ( .A(
        \dp/wr_data_id_i [8]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4252 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U629  ( .A(
        \dp/wr_data_id_i [7]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4251 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U628  ( .A(
        \dp/wr_data_id_i [6]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4250 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U627  ( .A(
        \dp/wr_data_id_i [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4249 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U626  ( .A(
        \dp/wr_data_id_i [4]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4248 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U625  ( .A(
        \dp/wr_data_id_i [3]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4247 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U624  ( .A(
        \dp/wr_data_id_i [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4246 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U623  ( .A(
        \dp/wr_data_id_i [1]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4245 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U622  ( .A(
        \dp/wr_data_id_i [0]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4244 ) );
  NOR3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U621  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [1]), .A2(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1194 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1339 ) );
  NOR3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U620  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [1]), .A2(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]), .A3(
        \dp/id_stage/regfile/DataPath/mux_wr_out [0]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1341 ) );
  NOR3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U619  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_wr_out [0]), .A2(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1193 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1305 ) );
  NOR3_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U618  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1194 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_wr_out [2]), .A3(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1193 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1270 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U617  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1176 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U616  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1175 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U615  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3158 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2607 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U614  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3178 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2600 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U613  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3176 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2595 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U612  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3166 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2574 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U611  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3162 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2568 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U610  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3155 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2564 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U609  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2551 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1978 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U608  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2549 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1974 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U607  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2535 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1948 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U606  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3178 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2605 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U605  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3158 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2606 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U604  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3162 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2570 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U603  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3162 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2569 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U602  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3155 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2563 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U601  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3175 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2596 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U600  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3175 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2594 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U599  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3173 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2590 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U598  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3173 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2589 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U597  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2538 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4241 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2535 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U596  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3165 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1197 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3162 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U595  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2528 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1938 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U594  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2531 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1933 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U593  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3155 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2565 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U592  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3178 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2602 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U591  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3176 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2597 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U590  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3166 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2571 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U589  ( .A(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4241 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U588  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2539 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2533 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1950 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U587  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3166 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2577 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U586  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3178 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2603 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U585  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3176 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2598 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U584  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3166 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2572 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U583  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3155 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2566 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U582  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3158 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2561 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U581  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2552 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4241 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2549 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U580  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3179 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1197 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3176 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U579  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3163 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1197 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3158 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U578  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2552 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [2]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2551 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U577  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1195 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1196 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3165 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U576  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [2]), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2538 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2539 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U575  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3175 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2591 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U574  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3175 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2592 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U573  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3173 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2586 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U572  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3173 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3156 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2587 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U571  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1975 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3813 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U570  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1970 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3825 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U569  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1964 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3840 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U568  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1959 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3852 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U567  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1949 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3867 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U566  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1944 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3879 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U565  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2576 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3759 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U564  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1976 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3809 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U563  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1971 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3821 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U562  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1965 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3836 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U561  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1960 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3848 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U560  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1945 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3875 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U559  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1939 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3890 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U558  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1934 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3902 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U557  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1976 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3810 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U556  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1971 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3822 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U555  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1965 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3837 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U554  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1960 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3849 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U553  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1945 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3876 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U552  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1939 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3891 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U551  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1934 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3903 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U550  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1980 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3802 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U549  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1969 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3829 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U548  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1954 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3856 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U547  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1943 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3883 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U546  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2581 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3748 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U545  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1937 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3898 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U544  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1963 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3844 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U543  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1979 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3805 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U542  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1968 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3832 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U541  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1953 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3859 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U540  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1942 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3886 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U539  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2580 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3751 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U538  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1975 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3814 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U537  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1970 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3826 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U536  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1964 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3841 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U535  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1959 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3853 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U534  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1949 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3868 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U533  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1944 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3880 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U532  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2576 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3760 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U531  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1973 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3820 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U530  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1947 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3874 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U529  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1936 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3901 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U528  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1962 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3847 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U527  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1967 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3835 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U526  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1952 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3862 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U525  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1941 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3889 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U524  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2579 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3754 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U523  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1976 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3811 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U522  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1971 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3823 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U521  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1965 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3838 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U520  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1960 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3850 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U519  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1945 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3877 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U518  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1939 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3892 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U517  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1934 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3904 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U516  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1980 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3800 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U515  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1969 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3827 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U514  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1954 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3854 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U513  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1943 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3881 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U512  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2581 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3746 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U511  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1980 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3801 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U510  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1969 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3828 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U509  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1954 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3855 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U508  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1943 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3882 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U507  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2581 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3747 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U506  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1963 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3842 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U505  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1937 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3896 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U504  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1963 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3843 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U503  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1937 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3897 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U502  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1979 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3803 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U501  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1968 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3830 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U500  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1953 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3857 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U499  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1942 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3884 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U498  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2580 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3749 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U497  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1979 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3804 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U496  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1968 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3831 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U495  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1953 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3858 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U494  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1942 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3885 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U493  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2580 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3750 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U492  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1975 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3812 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U491  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1970 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3824 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U490  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1964 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3839 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U489  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1959 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3851 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U488  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1949 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3866 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U487  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1944 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3878 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U486  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2576 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3758 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U485  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1973 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3818 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U484  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1962 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3845 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U483  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1947 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3872 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U482  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1936 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3899 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U481  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1973 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3819 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U480  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1962 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3846 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U479  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1947 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3873 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U478  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1936 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3900 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U477  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1967 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3833 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U476  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1952 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3860 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U475  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1941 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3887 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U474  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2579 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3752 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U473  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1967 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3834 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U472  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1952 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3861 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U471  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1941 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3888 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U470  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2579 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3753 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U469  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1198 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1199 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U468  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3970 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U467  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3979 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U466  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4024 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U465  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4051 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U464  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4096 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U463  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4105 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U462  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4168 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U461  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4213 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U460  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4222 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U459  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3934 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U458  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3943 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U457  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3988 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U456  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4015 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U455  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4060 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U454  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4069 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U453  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4132 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U452  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4141 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U451  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4150 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U450  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4159 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U449  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3952 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U448  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3961 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U447  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4033 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U446  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4042 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U445  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4114 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U444  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4123 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U443  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4177 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U442  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4186 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U441  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4195 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U440  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3916 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U439  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3925 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U438  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3997 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U437  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4006 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U436  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4078 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U435  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4087 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U434  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4204 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U433  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3969 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U432  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3968 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U431  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3967 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U430  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3966 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U429  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3965 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U428  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1825 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3964 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U427  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3978 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U426  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3977 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U425  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3976 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U424  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3975 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U423  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3974 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U422  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1791 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3973 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U421  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4023 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U420  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4022 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U419  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4021 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U418  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4020 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U417  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4019 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U416  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1690 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4018 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U415  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4050 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U414  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4049 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U413  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4048 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U412  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4047 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U411  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4046 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U410  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1654 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4045 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U409  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4095 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U408  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4094 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U407  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4093 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U406  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4092 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U405  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4091 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U404  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1553 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4090 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U403  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4104 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U402  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4103 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U401  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4102 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U400  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4101 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U399  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4100 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U398  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1520 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4099 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U397  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4167 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U396  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4166 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U395  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4165 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U394  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4164 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U393  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4163 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U392  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1351 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4162 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U391  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4212 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U390  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4211 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U389  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4210 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U388  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4209 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U387  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4208 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U386  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1307 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4207 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U385  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4221 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U384  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4220 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U383  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4219 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U382  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4218 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U381  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4217 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U380  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1273 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4216 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U379  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4230 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U378  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4229 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U377  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4228 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U376  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4227 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U375  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4226 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U374  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4225 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U373  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3933 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U372  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3932 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U371  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3931 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U370  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3930 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U369  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3929 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U368  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1893 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3928 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U367  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3942 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U366  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3941 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U365  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3940 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U364  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3939 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U363  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3938 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U362  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1860 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3937 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U361  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3987 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U360  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3986 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U359  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3985 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U358  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3984 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U357  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3983 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U356  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1758 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3982 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U355  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4014 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U354  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4013 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U353  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4012 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U352  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4011 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U351  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4010 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U350  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1723 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4009 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U349  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4059 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U348  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4058 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U347  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4057 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U346  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4056 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U345  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4055 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U344  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1621 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4054 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U343  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4068 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U342  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4067 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U341  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4066 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U340  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4065 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U339  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4064 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U338  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1588 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4063 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U337  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4131 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U336  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4130 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U335  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4129 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U334  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4128 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U333  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4127 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U332  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1484 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4126 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U331  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4140 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U330  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4139 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U329  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4138 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U328  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4137 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U327  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4136 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U326  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1451 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4135 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U325  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4149 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U324  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4148 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U323  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4147 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U322  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4146 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U321  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4145 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U320  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1418 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4144 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U319  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4158 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U318  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4157 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U317  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4156 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U316  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4155 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U315  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4154 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U314  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1385 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4153 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U313  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3946 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U312  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3947 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U311  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3948 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U310  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3949 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U309  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3950 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U308  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1166 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3951 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U307  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3955 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U306  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3956 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U305  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3957 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U304  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3958 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U303  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3959 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U302  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1165 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3960 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U301  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4027 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U300  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4028 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U299  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4029 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U298  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4030 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U297  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4031 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U296  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1164 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4032 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U295  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4036 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U294  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4037 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U293  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4038 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U292  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4039 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U291  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4040 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U290  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1163 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4041 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U289  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4108 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U288  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4109 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U287  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4110 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U286  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4111 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U285  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4112 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U284  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1162 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4113 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U283  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4117 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U282  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4118 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U281  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4119 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U280  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4120 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U279  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4121 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U278  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1161 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4122 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U277  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4171 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U276  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4172 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U275  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4173 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U274  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4174 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U273  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4175 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U272  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1168 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4176 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U271  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4180 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U270  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4181 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U269  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4182 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U268  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4183 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U267  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4184 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U266  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4185 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U265  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4189 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U264  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4190 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U263  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4191 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U262  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4192 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U261  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4193 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U260  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1167 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4194 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U259  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3910 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U258  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3911 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U257  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3912 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U256  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3913 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U255  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3914 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U254  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1160 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3915 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U253  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3919 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U252  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3920 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U251  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3921 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U250  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3922 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U249  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3923 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U248  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1159 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3924 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U247  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3991 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U246  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3992 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U245  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3993 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U244  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3994 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U243  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3995 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U242  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1158 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3996 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U241  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4000 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U240  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4001 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U239  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4002 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U238  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4003 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U237  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4004 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U236  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1157 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4005 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U235  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4072 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U234  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4073 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U233  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4074 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U232  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4075 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U231  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4076 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U230  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1156 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4077 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U229  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4081 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U228  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4082 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U227  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4083 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U226  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4084 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U225  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4085 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U224  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1155 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4086 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U223  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4198 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U222  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4199 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U221  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4200 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U220  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4201 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U219  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4202 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U218  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1154 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4203 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U217  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1238 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4231 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U216  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1176 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1169 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U215  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1176 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1170 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U214  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1176 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1171 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U213  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1175 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1172 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U212  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1175 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1173 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U211  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1175 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1174 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U210  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3176 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2601 ) );
  AND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U209  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3162 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2575 ) );
  NAND2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U208  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3158 ), .A2(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3160 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2560 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U207  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1938 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3894 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U206  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1933 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3906 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U205  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2602 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3705 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U204  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2597 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3717 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U203  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2591 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3732 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U202  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2586 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3744 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U201  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2571 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3771 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U200  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2565 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3786 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U199  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1950 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3863 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U198  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2603 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3701 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U197  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2598 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3713 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U196  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2592 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3728 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U195  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2587 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3740 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U194  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2577 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3755 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U193  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2572 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3767 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U192  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2566 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3782 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U191  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2561 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3794 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U190  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1950 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3864 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U189  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2603 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3702 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U188  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2598 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3714 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U187  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2592 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3729 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U186  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2587 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3741 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U185  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2577 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3756 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U184  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2572 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3768 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U183  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2566 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3783 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U182  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2561 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3795 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U181  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2607 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3694 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U180  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2596 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3721 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U179  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2570 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3775 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U178  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1974 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3817 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U177  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1948 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3871 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U176  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2564 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3790 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U175  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2590 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3736 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U174  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2606 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3697 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U173  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2595 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3724 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U172  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2569 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3778 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U171  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1938 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3895 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U170  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1933 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3907 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U169  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2602 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3706 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U168  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2597 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3718 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U167  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2591 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3733 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U166  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2586 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3745 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U165  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2571 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3772 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U164  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2565 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3787 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U163  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2600 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3712 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U162  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2574 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3766 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U161  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2589 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3739 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U160  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2563 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3793 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U159  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1978 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3808 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U158  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2605 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3700 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U157  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2594 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3727 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U156  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2568 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3781 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U155  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1950 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3865 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U154  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2603 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3703 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U153  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2598 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3715 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U152  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2592 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3730 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U151  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2587 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3742 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U150  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2577 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3757 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U149  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2572 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3769 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U148  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2566 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3784 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U147  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2561 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3796 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U146  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2607 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1926 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U145  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2596 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3719 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U144  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2570 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3773 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U143  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2607 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3693 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U142  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2596 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3720 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U141  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2570 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3774 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U140  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1974 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3815 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U139  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1948 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3869 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U138  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2590 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3734 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U137  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2564 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3788 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U136  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1974 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3816 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U135  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1948 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3870 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U134  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2590 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3735 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U133  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2564 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3789 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U132  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2606 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3695 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U131  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2595 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3722 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U130  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2569 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3776 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U129  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2606 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3696 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U128  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2595 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3723 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U127  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2569 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3777 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U126  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1938 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3893 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U125  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1933 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3905 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U124  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2602 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3704 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U123  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2597 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3716 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U122  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2591 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3731 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U121  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2586 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3743 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U120  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2571 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3770 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U119  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2565 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3785 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U118  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2600 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3710 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U117  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2589 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3737 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U116  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2574 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3764 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U115  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2563 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3791 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U114  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2600 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3711 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U113  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2589 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3738 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U112  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2574 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3765 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U111  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2563 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3792 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U110  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1978 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3806 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U109  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2605 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3698 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U108  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2594 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3725 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U107  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2568 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3779 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U106  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1978 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3807 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U105  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2605 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3699 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U104  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2594 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3726 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U103  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2568 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3780 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U102  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4231 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4224 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U101  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4231 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4223 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U100  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3916 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3908 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U99  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3916 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3909 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U98  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3925 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3917 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U97  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3925 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3918 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U96  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3952 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3944 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U95  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3952 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3945 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U94  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3961 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3953 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U93  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3961 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3954 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U92  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3997 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3989 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U91  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3997 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3990 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U90  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4006 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3998 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U89  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4006 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3999 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U88  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4033 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4025 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U87  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4033 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4026 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U86  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4042 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4034 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U85  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4042 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4035 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U84  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4078 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4070 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U83  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4078 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4071 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U82  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4087 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4079 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U81  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4087 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4080 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U80  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4114 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4106 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U79  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4114 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4107 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U78  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4123 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4115 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U77  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4123 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4116 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U76  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4177 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4169 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U75  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4177 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4170 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U74  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4186 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4178 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U73  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4186 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4179 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U72  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4195 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4187 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U71  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4195 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4188 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U70  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4204 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4196 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U69  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4204 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4197 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U68  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3934 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3927 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U67  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3934 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3926 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U66  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3943 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3936 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U65  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3943 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3935 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U64  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3970 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3963 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U63  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3970 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3962 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U62  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3979 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3972 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U61  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3979 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3971 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U60  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3988 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3981 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U59  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3988 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3980 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U58  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4015 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4008 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U57  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4015 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4007 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U56  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4024 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4017 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U55  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4024 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4016 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U54  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4051 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4044 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U53  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4051 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4043 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U52  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4060 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4053 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U51  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4060 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4052 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U50  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4069 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4062 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U49  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4069 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4061 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U48  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4096 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4089 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U47  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4096 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4088 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U46  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4105 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4098 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U45  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4105 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4097 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U44  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4132 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4125 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U43  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4132 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4124 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U42  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4141 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4134 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U41  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4141 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4133 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U40  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4150 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4143 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U39  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4150 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4142 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U38  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4152 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U37  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4159 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4151 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U36  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4168 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4161 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U35  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4168 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4160 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U34  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4213 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4206 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U33  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4213 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4205 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U32  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4222 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4215 ) );
  INV_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U31  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4222 ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4214 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U30  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1169 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1346 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U29  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1169 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1348 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U28  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1170 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1516 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U27  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1170 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1518 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U26  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1171 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1585 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U25  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1171 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1586 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U24  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1171 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1687 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U23  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1172 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1688 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U22  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1172 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1755 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U21  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1172 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1756 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U20  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1173 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1857 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U19  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1174 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1858 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U18  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1174 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1925 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U17  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2560 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3798 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U16  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2601 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3709 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U15  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2575 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3763 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U14  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2560 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3799 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U13  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2601 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3707 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U12  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2575 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3761 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U11  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2601 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3708 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U10  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2575 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3762 ) );
  BUF_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U9  ( .A(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2560 ), .Z(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3797 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U8  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4242 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [0]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2532 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U7  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4276 ), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [1]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2530 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U6  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1198 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [0]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3159 ) );
  NOR2_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U5  ( .A1(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1199 ), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [1]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3157 ) );
  INV_X32 \dp/id_stage/regfile/DataPath/Physical_RF/U4  ( .A(
        \dp/id_stage/regfile/rst_rf ), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U3  ( .A1(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [2]), .A2(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [3]), .A3(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [4]), .A4(
        \dp/id_stage/regfile/DataPath/addr_rd2_p [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2546 ) );
  NOR4_X1 \dp/id_stage/regfile/DataPath/Physical_RF/U2  ( .A1(
        \dp/id_stage/regfile/DataPath/mux_rd_out [2]), .A2(
        \dp/id_stage/regfile/DataPath/mux_rd_out [3]), .A3(
        \dp/id_stage/regfile/DataPath/mux_rd_out [4]), .A4(
        \dp/id_stage/regfile/DataPath/mux_rd_out [5]), .ZN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3173 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n111 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n367 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n879 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1071 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1103 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n128 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n127 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n126 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n125 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n124 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n123 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n122 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n121 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n120 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n110 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n109 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n108 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n107 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n106 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n384 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n383 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n382 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n381 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n380 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n379 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n378 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n377 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n376 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n366 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n365 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n364 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n363 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n362 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n896 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n895 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n894 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n893 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n892 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n891 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n890 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n889 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n888 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n878 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n877 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n876 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n875 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n874 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n129 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n119 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n118 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n117 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n116 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n115 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n114 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n113 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n112 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n385 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n375 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n374 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n373 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n372 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n371 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n370 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n369 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n368 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n897 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n887 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n886 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n885 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n884 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n883 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n882 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n881 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n880 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1088 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1087 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1086 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1085 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1084 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1083 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1082 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1081 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1080 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1070 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1069 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1068 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1067 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1066 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1120 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1119 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1118 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1117 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1116 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1115 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1114 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1113 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1112 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1102 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1101 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1100 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1099 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1098 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1089 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1079 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1078 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1077 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1076 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1075 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1074 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1073 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1072 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1121 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1111 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1110 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1109 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1108 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1107 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1106 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1105 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1104 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1135 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n271 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n527 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n783 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n79 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n559 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n815 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n847 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1153 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1152 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1151 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1150 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1149 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1148 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1147 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1146 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1145 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1144 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1143 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1142 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1141 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1140 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1139 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1138 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1137 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1136 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1134 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1133 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1132 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n288 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n287 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n286 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n285 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n284 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n283 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n282 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n281 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n280 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n270 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n269 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n268 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n267 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n266 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n544 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n543 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n542 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n541 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n540 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n539 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n538 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n537 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n536 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n526 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n525 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n524 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n523 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n522 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n800 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n799 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n798 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n797 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n796 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n795 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n794 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n793 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n792 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n782 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n781 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n780 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n779 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n778 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n289 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n279 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n278 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n277 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n276 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n275 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n274 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n273 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n272 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n545 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n535 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n534 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n533 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n532 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n531 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n530 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n529 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n528 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n801 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n791 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n790 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n789 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n788 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n787 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n786 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n785 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n784 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n96 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n95 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n94 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n93 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n92 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n91 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n90 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n89 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n88 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n78 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n77 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n76 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n75 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n74 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n576 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n575 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n574 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n573 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n572 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n571 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n570 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n569 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n568 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n558 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n557 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n556 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n555 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n554 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n832 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n831 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n830 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n829 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n828 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n827 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n826 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n825 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n824 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n814 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n813 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n812 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n811 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n810 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n864 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n863 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n862 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n861 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n860 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n859 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n858 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n857 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n856 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n846 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n845 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n844 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n843 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n842 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n97 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n87 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n86 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n85 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n84 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n83 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n82 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n81 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n80 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n577 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n567 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n566 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n565 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n564 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n563 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n562 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n561 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n560 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n833 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n823 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n822 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n821 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n820 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n819 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n818 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n817 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n816 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n865 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n855 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n854 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n853 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n852 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n851 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n850 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n849 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n848 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1126 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1122 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1131 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1130 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1129 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1128 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1127 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1125 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1124 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[35][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1123 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[35][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n655 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n687 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n207 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n239 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n672 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n671 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n670 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n669 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n668 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n667 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n666 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n665 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n664 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n654 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n653 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n652 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n651 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n650 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n704 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n703 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n702 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n701 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n700 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n699 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n698 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n697 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n696 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n686 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n685 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n684 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n683 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n682 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n673 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n663 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n662 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n661 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n660 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n659 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n658 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n657 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n656 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n705 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n695 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n694 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n693 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n692 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n691 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n690 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n689 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n688 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n224 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n223 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n222 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n221 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n220 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n219 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n218 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n217 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n216 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n206 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n205 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n204 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n203 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n202 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n256 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n255 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n254 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n253 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n252 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n251 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n250 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n249 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n248 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n238 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n237 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n236 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n235 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n234 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n225 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n215 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n214 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n213 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n212 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n211 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n210 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n209 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n208 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n257 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n247 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n246 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n245 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n244 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n243 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n242 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n241 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n240 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n102 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n98 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n358 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n354 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n870 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n866 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1062 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1058 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1094 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1090 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n105 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n104 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n103 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n101 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n100 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[3][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n99 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[3][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n361 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n360 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n359 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n357 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n356 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[11][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n355 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[11][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n873 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n872 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n871 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n869 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n868 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[27][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n867 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[27][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1065 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1064 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1063 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1061 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1060 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[33][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1059 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[33][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1097 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1096 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1095 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1093 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1092 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[34][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n1091 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[34][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n262 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n258 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n518 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n514 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n774 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n770 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n70 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n66 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n550 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n546 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n806 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n802 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n838 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n834 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n265 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n264 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n263 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n261 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n260 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[8][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n259 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[8][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n521 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n520 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n519 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n517 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n516 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[16][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n515 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[16][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n777 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n776 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n775 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n773 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n772 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[24][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n771 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[24][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n73 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n72 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n71 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n69 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n68 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[2][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n67 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[2][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n553 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n552 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n551 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n549 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n548 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[17][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n547 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[17][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n809 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n808 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n807 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n805 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n804 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[25][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n803 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[25][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n841 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n840 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n839 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n837 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n836 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[26][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n835 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[26][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n646 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n642 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n678 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n674 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n198 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n194 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n230 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n226 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n399 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n649 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n648 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n647 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n645 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n644 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[20][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n643 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[20][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n681 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n680 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n679 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n677 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n676 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[21][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n675 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[21][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n911 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n201 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n200 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n199 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n197 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n196 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[6][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n195 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[6][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n233 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n232 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n231 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n229 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n228 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[7][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n227 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[7][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n416 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n415 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n414 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n413 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n412 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n411 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n410 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n409 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n408 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n398 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n397 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n396 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n395 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n394 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n417 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n407 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n406 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n405 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n404 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n403 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n402 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n401 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n400 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n928 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n927 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n926 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n925 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n924 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n923 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n922 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n921 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n920 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n910 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n909 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n908 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n907 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n906 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n929 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n919 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n918 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n917 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n916 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n915 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n914 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n913 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n912 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n495 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][18] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n512 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][1] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n511 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][2] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n510 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][3] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n509 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][4] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n508 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][5] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n507 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][6] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n506 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][7] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n505 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][8] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n504 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][9] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n494 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][19] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n493 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][20] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n492 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][21] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n491 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][22] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n490 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][23] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n513 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][0] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n503 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][10] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n502 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][11] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n501 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][12] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n500 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][13] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n499 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][14] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n498 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][15] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n497 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][16] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n496 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][17] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n390 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n386 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n902 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n898 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n393 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n392 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n391 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n389 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n388 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[12][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n387 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[12][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n905 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n904 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n903 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n901 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n900 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[28][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n899 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[28][30] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n486 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][27] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n482 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][31] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n489 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][24] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n488 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][25] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n487 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][26] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n485 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][28] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n484 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][29] ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[15][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n483 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4243 ), .Q(
        \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS[15][30] ) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[0]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4239 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N359 ), .Q(
        \dp/id_stage/out1_i [0]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[0]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4235 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N427 ), .Q(
        \dp/id_stage/out2_i [0]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[1]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4239 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N358 ), .Q(
        \dp/id_stage/out1_i [1]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[1]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4235 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N426 ), .Q(
        \dp/id_stage/out2_i [1]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[2]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N357 ), .Q(
        \dp/id_stage/out1_i [2]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[2]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N425 ), .Q(
        \dp/id_stage/out2_i [2]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[3]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N356 ), .Q(
        \dp/id_stage/out1_i [3]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[3]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N424 ), .Q(
        \dp/id_stage/out2_i [3]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[4]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N355 ), .Q(
        \dp/id_stage/out1_i [4]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[4]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N423 ), .Q(
        \dp/id_stage/out2_i [4]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[5]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N354 ), .Q(
        \dp/id_stage/out1_i [5]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[5]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N422 ), .Q(
        \dp/id_stage/out2_i [5]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[6]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N353 ), .Q(
        \dp/id_stage/out1_i [6]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[6]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N421 ), .Q(
        \dp/id_stage/out2_i [6]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[7]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N352 ), .Q(
        \dp/id_stage/out1_i [7]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[7]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N420 ), .Q(
        \dp/id_stage/out2_i [7]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[8]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N351 ), .Q(
        \dp/id_stage/out1_i [8]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[8]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N419 ), .Q(
        \dp/id_stage/out2_i [8]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[9]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N350 ), .Q(
        \dp/id_stage/out1_i [9]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[9]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N418 ), .Q(
        \dp/id_stage/out2_i [9]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[10]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N349 ), .Q(
        \dp/id_stage/out1_i [10]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[10]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N417 ), .Q(
        \dp/id_stage/out2_i [10]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[11]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4238 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N348 ), .Q(
        \dp/id_stage/out1_i [11]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[11]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4234 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N416 ), .Q(
        \dp/id_stage/out2_i [11]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[12]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N347 ), .Q(
        \dp/id_stage/out1_i [12]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[12]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N415 ), .Q(
        \dp/id_stage/out2_i [12]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[13]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N346 ), .Q(
        \dp/id_stage/out1_i [13]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[13]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N414 ), .Q(
        \dp/id_stage/out2_i [13]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[14]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N345 ), .Q(
        \dp/id_stage/out1_i [14]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[14]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N413 ), .Q(
        \dp/id_stage/out2_i [14]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[15]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N344 ), .Q(
        \dp/id_stage/out1_i [15]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[15]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N412 ), .Q(
        \dp/id_stage/out2_i [15]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[16]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N343 ), .Q(
        \dp/id_stage/out1_i [16]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[16]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N411 ), .Q(
        \dp/id_stage/out2_i [16]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[17]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N342 ), .Q(
        \dp/id_stage/out1_i [17]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[17]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N410 ), .Q(
        \dp/id_stage/out2_i [17]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[18]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N341 ), .Q(
        \dp/id_stage/out1_i [18]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[18]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N409 ), .Q(
        \dp/id_stage/out2_i [18]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[19]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N340 ), .Q(
        \dp/id_stage/out1_i [19]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[19]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N408 ), .Q(
        \dp/id_stage/out2_i [19]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[20]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N339 ), .Q(
        \dp/id_stage/out1_i [20]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[20]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N407 ), .Q(
        \dp/id_stage/out2_i [20]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[21]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4237 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N338 ), .Q(
        \dp/id_stage/out1_i [21]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[21]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4233 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N406 ), .Q(
        \dp/id_stage/out2_i [21]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[22]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N337 ), .Q(
        \dp/id_stage/out1_i [22]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[22]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N405 ), .Q(
        \dp/id_stage/out2_i [22]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[23]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N336 ), .Q(
        \dp/id_stage/out1_i [23]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[23]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N404 ), .Q(
        \dp/id_stage/out2_i [23]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[24]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N335 ), .Q(
        \dp/id_stage/out1_i [24]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[24]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N403 ), .Q(
        \dp/id_stage/out2_i [24]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[25]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N334 ), .Q(
        \dp/id_stage/out1_i [25]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[25]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N402 ), .Q(
        \dp/id_stage/out2_i [25]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[26]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N333 ), .Q(
        \dp/id_stage/out1_i [26]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[26]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N401 ), .Q(
        \dp/id_stage/out2_i [26]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[27]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N332 ), .Q(
        \dp/id_stage/out1_i [27]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[27]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N400 ), .Q(
        \dp/id_stage/out2_i [27]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[28]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N331 ), .Q(
        \dp/id_stage/out1_i [28]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[28]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N399 ), .Q(
        \dp/id_stage/out2_i [28]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[29]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N330 ), .Q(
        \dp/id_stage/out1_i [29]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[29]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N398 ), .Q(
        \dp/id_stage/out2_i [29]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[30]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N329 ), .Q(
        \dp/id_stage/out1_i [30]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[30]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N397 ), .Q(
        \dp/id_stage/out2_i [30]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT1_reg[31]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4236 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N328 ), .Q(
        \dp/id_stage/out1_i [31]) );
  DLH_X1 \dp/id_stage/regfile/DataPath/Physical_RF/OUT2_reg[31]  ( .G(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4232 ), .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/N396 ), .Q(
        \dp/id_stage/out2_i [31]) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3181 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1177 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1057 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3182 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1177 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1056 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3183 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1177 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1055 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3184 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1054 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3185 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1053 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3186 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1052 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3187 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1051 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3188 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1050 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3189 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1049 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3190 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1048 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3191 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1047 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3192 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1046 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3193 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1045 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3194 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1178 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1044 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3195 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1043 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3196 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1042 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3197 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1041 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3198 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1040 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3199 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1039 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3200 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1038 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3201 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1037 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3202 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1036 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3203 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1035 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3204 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1034 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3205 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1179 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1033 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3206 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1032 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3207 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1031 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3208 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1030 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3209 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1029 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3210 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1028 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3211 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1027 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[32][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3212 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1026 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3213 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1025 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3214 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1024 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3215 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1023 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3216 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1180 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1022 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3217 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1021 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3218 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1020 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3219 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1019 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3220 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1018 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3221 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1017 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3222 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1016 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3223 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1015 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3224 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1014 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3225 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1013 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3226 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1012 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3227 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1181 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1011 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3228 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1010 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3229 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1009 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3230 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1008 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3231 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1007 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3232 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1006 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3233 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1005 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3234 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1004 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3235 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1003 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3236 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1002 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3237 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1001 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3238 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1182 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1000 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3239 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n999 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3240 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n998 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3241 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n997 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3242 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n996 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3243 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n995 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[31][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3244 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n994 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3245 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n993 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3246 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n992 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3247 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n991 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3248 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n990 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3249 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1183 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n989 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3250 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n988 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3251 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n987 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3252 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n986 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3253 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n985 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3254 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n984 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3255 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n983 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3256 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n982 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3257 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n981 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3258 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n980 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3259 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n979 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3260 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1184 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n978 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3261 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n977 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3262 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n976 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3263 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n975 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3264 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n974 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3265 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n973 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3266 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n972 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3267 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n971 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3268 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n970 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3269 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n969 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3270 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n968 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3271 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1185 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n967 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3272 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n966 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3273 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n965 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3274 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n964 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3275 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n963 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[30][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3276 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n962 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3277 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n961 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3278 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n960 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3279 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n959 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3280 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n958 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3281 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n957 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3282 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1186 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n956 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3283 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n955 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3284 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n954 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3285 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n953 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3286 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n952 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3287 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n951 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3288 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n950 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3289 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n949 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3290 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n948 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3291 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n947 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3292 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n946 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3293 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1187 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n945 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3294 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n944 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3295 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n943 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3296 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n942 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3297 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n941 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3298 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n940 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3299 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n939 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3300 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n938 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3301 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n937 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3302 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n936 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3303 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n935 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3304 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1188 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n934 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3305 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1189 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n933 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3306 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1189 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n932 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3307 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1189 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n931 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[29][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3308 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1189 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n930 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3309 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1172 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n769 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3310 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n768 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3311 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n767 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3312 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n766 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3313 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n765 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3314 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n764 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3315 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n763 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3316 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n762 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3317 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n761 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3318 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n760 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3319 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n759 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3320 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1200 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n758 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3321 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n757 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3322 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n756 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3323 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n755 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3324 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n754 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3325 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n753 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3326 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n752 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3327 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n751 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3328 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n750 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3329 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n749 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3330 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n748 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3331 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1202 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n747 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3332 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n746 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3333 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n745 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3334 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n744 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3335 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n743 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3336 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n742 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3337 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n741 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3338 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n740 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3339 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n739 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[23][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3340 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n738 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3341 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n737 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3342 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1203 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n736 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3343 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n735 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3344 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n734 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3345 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n733 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3346 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n732 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3347 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n731 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3348 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n730 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3349 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n729 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3350 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n728 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3351 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n727 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3352 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n726 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3353 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1204 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n725 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3354 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n724 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3355 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n723 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3356 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n722 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3357 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n721 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3358 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n720 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3359 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n719 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3360 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n718 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3361 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n717 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3362 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n716 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3363 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n715 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3364 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1205 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n714 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3365 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n713 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3366 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n712 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3367 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n711 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3368 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n710 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3369 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n709 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3370 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n708 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3371 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n707 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[22][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3372 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1206 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n706 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3373 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1207 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n641 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3374 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1207 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n640 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3375 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1207 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n639 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3376 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1207 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n638 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3377 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1207 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n637 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3378 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n636 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3379 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n635 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3380 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n634 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3381 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n633 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3382 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n632 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3383 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n631 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3384 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n630 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3385 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n629 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3386 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n628 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3387 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n627 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3388 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1208 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n626 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3389 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n625 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3390 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n624 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3391 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n623 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3392 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n622 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3393 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n621 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3394 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n620 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3395 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n619 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3396 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n618 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3397 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n617 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3398 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n616 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3399 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1209 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n615 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3400 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n614 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3401 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n613 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3402 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n612 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3403 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n611 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[19][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3404 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n610 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3405 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n609 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3406 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n608 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3407 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n607 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3408 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n606 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3409 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n605 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3410 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1210 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n604 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3411 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n603 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3412 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n602 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3413 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n601 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3414 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n600 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3415 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n599 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3416 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n598 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3417 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n597 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3418 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n596 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3419 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n595 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3420 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n594 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3421 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1211 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n593 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3422 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n592 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3423 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n591 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3424 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n590 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3425 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n589 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3426 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n588 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3427 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n587 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3428 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n586 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3429 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n585 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3430 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n584 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3431 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n583 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3432 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1212 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n582 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3433 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1213 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n581 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3434 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1213 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n580 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3435 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1213 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n579 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[18][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3436 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1213 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n578 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3437 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n481 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3438 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n480 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3439 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n479 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3440 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n478 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3441 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n477 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3442 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n476 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3443 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n475 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3444 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n474 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3445 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n473 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3446 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1214 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n472 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3447 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n471 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3448 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n470 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3449 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n469 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3450 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n468 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3451 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n467 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3452 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n466 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3453 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n465 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3454 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n464 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3455 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n463 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3456 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n462 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3457 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1215 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n461 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3458 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n460 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3459 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n459 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3460 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n458 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3461 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n457 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3462 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n456 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3463 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n455 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3464 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n454 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3465 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n453 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3466 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n452 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3467 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n451 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[14][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3468 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1216 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n450 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3469 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n449 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3470 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n448 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3471 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n447 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3472 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n446 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3473 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n445 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3474 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n444 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3475 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n443 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3476 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n442 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3477 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n441 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3478 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n440 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3479 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1217 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n439 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3480 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n438 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3481 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n437 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3482 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n436 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3483 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n435 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3484 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n434 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3485 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n433 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3486 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n432 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3487 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n431 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3488 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n430 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3489 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n429 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3490 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1218 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n428 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3491 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n427 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3492 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n426 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3493 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n425 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3494 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n424 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3495 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n423 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3496 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n422 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3497 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n421 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3498 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n420 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3499 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n419 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[13][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3500 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1219 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n418 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][0]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3501 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1220 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n353 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][1]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3502 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1220 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n352 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][2]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3503 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1220 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n351 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][3]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3504 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n350 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][4]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3505 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n349 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][5]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3506 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n348 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][6]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3507 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n347 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][7]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3508 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n346 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][8]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3509 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n345 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][9]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3510 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n344 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3511 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n343 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3512 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n342 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3513 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n341 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3514 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1221 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n340 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3515 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n339 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3516 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n338 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3517 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n337 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3518 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n336 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3519 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n335 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3520 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n334 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3521 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n333 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3522 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n332 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3523 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n331 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3524 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n330 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3525 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1222 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n329 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3526 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n328 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3527 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n327 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3528 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n326 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3529 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n325 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3530 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n324 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3531 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n323 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[10][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3532 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n322 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3533 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n321 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3534 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n320 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3535 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n319 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3536 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1223 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n318 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3537 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n317 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3538 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n316 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3539 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n315 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3540 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n314 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3541 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n313 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3542 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n312 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3543 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n311 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3544 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n310 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3545 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n309 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3546 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n308 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3547 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1224 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n307 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3548 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n306 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3549 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n305 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3550 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n304 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3551 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n303 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3552 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n302 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3553 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n301 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3554 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n300 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3555 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n299 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3556 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n298 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3557 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n297 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3558 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1225 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n296 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3559 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1226 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n295 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3560 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1226 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n294 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3561 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1226 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n293 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3562 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1226 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n292 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3563 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1226 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n291 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[9][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3564 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1226 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n290 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3565 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n193 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3566 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n192 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3567 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n191 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3568 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n190 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3569 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n189 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3570 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n188 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3571 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n187 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3572 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1227 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n186 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3573 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n185 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3574 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n184 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3575 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n183 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3576 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n182 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3577 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n181 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3578 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n180 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3579 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n179 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3580 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n178 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3581 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n177 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3582 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n176 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3583 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1228 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n175 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3584 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n174 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3585 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n173 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3586 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n172 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3587 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n171 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3588 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n170 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3589 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n169 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3590 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n168 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3591 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n167 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3592 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n166 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3593 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n165 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3594 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1229 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n164 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3595 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n163 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[5][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3596 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n162 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3597 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n161 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3598 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n160 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3599 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n159 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3600 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n158 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3601 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n157 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3602 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n156 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3603 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n155 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3604 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n154 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3605 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1230 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n153 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3606 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n152 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3607 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n151 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3608 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n150 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3609 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n149 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3610 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n148 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3611 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n147 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3612 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n146 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3613 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n145 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3614 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n144 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3615 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n143 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3616 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1231 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n142 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3617 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n141 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3618 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n140 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3619 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n139 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3620 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n138 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3621 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n137 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3622 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n136 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3623 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n135 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3624 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n134 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3625 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n133 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3626 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n132 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3627 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1232 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n131 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[4][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3628 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1169 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n130 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3629 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1169 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n65 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3630 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n64 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3631 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n63 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3632 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n62 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3633 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n61 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3634 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n60 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3635 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n59 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3636 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n58 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3637 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n57 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3638 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n56 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3639 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n55 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3640 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1233 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n54 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3641 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n53 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3642 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n52 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3643 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n51 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3644 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n50 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3645 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n49 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3646 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n48 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3647 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n47 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3648 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n46 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3649 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n45 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3650 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n44 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3651 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1234 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n43 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3652 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n42 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3653 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n41 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3654 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n40 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3655 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n39 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3656 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n38 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3657 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n37 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3658 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n36 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3659 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n35 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[1][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3660 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n34 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][0]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3661 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n33 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][1]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3662 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1235 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n32 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][2]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3663 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n31 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][3]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3664 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n30 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][4]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3665 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n29 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][5]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3666 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n28 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][6]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3667 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n27 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][7]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3668 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n26 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][8]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3669 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n25 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][9]  ( .D(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3670 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n24 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][10]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3671 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n23 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][11]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3672 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n22 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][12]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3673 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1236 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n21 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][13]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3674 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n20 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][14]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3675 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n19 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][15]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3676 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n18 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][16]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3677 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n17 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][17]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3678 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n16 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][18]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3679 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n15 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][19]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3680 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n14 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][20]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3681 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n13 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][21]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3682 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n12 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][22]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3683 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n11 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][23]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3684 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1340 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n10 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][24]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3685 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n9 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][25]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3686 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n8 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][26]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3687 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n7 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][27]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3688 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n6 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][28]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3689 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n5 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][29]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3690 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n4 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][30]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3691 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n3 ) );
  DFFR_X1 \dp/id_stage/regfile/DataPath/Physical_RF/REGISTERS_reg[0][31]  ( 
        .D(\dp/id_stage/regfile/DataPath/Physical_RF/n3692 ), .CK(CLK), .RN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n1343 ), .QN(
        \dp/id_stage/regfile/DataPath/Physical_RF/n2 ) );
  NOR4_X1 \dp/ex_stage/U11  ( .A1(\dp/rf_out1_ex_i [1]), .A2(
        \dp/rf_out1_ex_i [19]), .A3(\dp/rf_out1_ex_i [18]), .A4(
        \dp/rf_out1_ex_i [17]), .ZN(\dp/ex_stage/n5 ) );
  NOR4_X1 \dp/ex_stage/U10  ( .A1(\dp/rf_out1_ex_i [16]), .A2(
        \dp/rf_out1_ex_i [15]), .A3(\dp/rf_out1_ex_i [14]), .A4(
        \dp/rf_out1_ex_i [13]), .ZN(\dp/ex_stage/n4 ) );
  NOR4_X1 \dp/ex_stage/U9  ( .A1(\dp/rf_out1_ex_i [12]), .A2(
        \dp/rf_out1_ex_i [11]), .A3(\dp/rf_out1_ex_i [10]), .A4(
        \dp/rf_out1_ex_i [0]), .ZN(\dp/ex_stage/n3 ) );
  NAND4_X1 \dp/ex_stage/U8  ( .A1(\dp/ex_stage/n3 ), .A2(\dp/ex_stage/n4 ), 
        .A3(\dp/ex_stage/n5 ), .A4(\dp/ex_stage/n6 ), .ZN(\dp/ex_stage/n2 ) );
  NAND4_X1 \dp/ex_stage/U7  ( .A1(\dp/ex_stage/n7 ), .A2(\dp/ex_stage/n8 ), 
        .A3(\dp/ex_stage/n9 ), .A4(\dp/ex_stage/n10 ), .ZN(\dp/ex_stage/n1 )
         );
  OR2_X1 \dp/ex_stage/U6  ( .A1(\dp/ex_stage/n1 ), .A2(\dp/ex_stage/n2 ), .ZN(
        \dp/branch_t_ex_o ) );
  NOR4_X1 \dp/ex_stage/U5  ( .A1(\dp/rf_out1_ex_i [27]), .A2(
        \dp/rf_out1_ex_i [26]), .A3(\dp/rf_out1_ex_i [25]), .A4(
        \dp/rf_out1_ex_i [24]), .ZN(\dp/ex_stage/n7 ) );
  NOR4_X1 \dp/ex_stage/U4  ( .A1(\dp/rf_out1_ex_i [30]), .A2(
        \dp/rf_out1_ex_i [2]), .A3(\dp/rf_out1_ex_i [29]), .A4(
        \dp/rf_out1_ex_i [28]), .ZN(\dp/ex_stage/n8 ) );
  NOR4_X1 \dp/ex_stage/U3  ( .A1(\dp/rf_out1_ex_i [5]), .A2(
        \dp/rf_out1_ex_i [4]), .A3(\dp/rf_out1_ex_i [3]), .A4(
        \dp/rf_out1_ex_i [31]), .ZN(\dp/ex_stage/n9 ) );
  NOR4_X1 \dp/ex_stage/U2  ( .A1(\dp/rf_out1_ex_i [9]), .A2(
        \dp/rf_out1_ex_i [8]), .A3(\dp/rf_out1_ex_i [7]), .A4(
        \dp/rf_out1_ex_i [6]), .ZN(\dp/ex_stage/n10 ) );
  NOR4_X1 \dp/ex_stage/U1  ( .A1(\dp/rf_out1_ex_i [23]), .A2(
        \dp/rf_out1_ex_i [22]), .A3(\dp/rf_out1_ex_i [21]), .A4(
        \dp/rf_out1_ex_i [20]), .ZN(\dp/ex_stage/n6 ) );
  AOI22_X1 \dp/ex_stage/muxA/U78  ( .A1(\dp/rf_out1_ex_i [17]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [17]), .B2(
        \dp/ex_stage/muxA/n11 ), .ZN(\dp/ex_stage/muxA/n87 ) );
  INV_X1 \dp/ex_stage/muxA/U77  ( .A(\dp/ex_stage/muxA/n87 ), .ZN(
        \dp/ex_stage/muxA_out [17]) );
  AOI22_X1 \dp/ex_stage/muxA/U76  ( .A1(\dp/rf_out1_ex_i [21]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [21]), .B2(
        \dp/ex_stage/muxA/n10 ), .ZN(\dp/ex_stage/muxA/n92 ) );
  INV_X1 \dp/ex_stage/muxA/U75  ( .A(\dp/ex_stage/muxA/n92 ), .ZN(
        \dp/ex_stage/muxA_out [21]) );
  AOI22_X1 \dp/ex_stage/muxA/U74  ( .A1(\dp/rf_out1_ex_i [23]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [23]), .B2(
        \dp/ex_stage/muxA/n9 ), .ZN(\dp/ex_stage/muxA/n94 ) );
  INV_X1 \dp/ex_stage/muxA/U73  ( .A(\dp/ex_stage/muxA/n94 ), .ZN(
        \dp/ex_stage/muxA_out [23]) );
  AOI22_X1 \dp/ex_stage/muxA/U72  ( .A1(\dp/rf_out1_ex_i [22]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [22]), .B2(
        \dp/ex_stage/muxA/n9 ), .ZN(\dp/ex_stage/muxA/n93 ) );
  INV_X1 \dp/ex_stage/muxA/U71  ( .A(\dp/ex_stage/muxA/n93 ), .ZN(
        \dp/ex_stage/muxA_out [22]) );
  AOI22_X1 \dp/ex_stage/muxA/U70  ( .A1(\dp/rf_out1_ex_i [29]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [29]), .B2(
        \dp/ex_stage/muxA/n8 ), .ZN(\dp/ex_stage/muxA/n100 ) );
  AOI22_X1 \dp/ex_stage/muxA/U69  ( .A1(\dp/rf_out1_ex_i [31]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [31]), .B2(
        \dp/ex_stage/muxA/n7 ), .ZN(\dp/ex_stage/muxA/n103 ) );
  INV_X1 \dp/ex_stage/muxA/U68  ( .A(\dp/ex_stage/muxA/n103 ), .ZN(
        \dp/ex_stage/alu/shifter/N136 ) );
  AOI22_X1 \dp/ex_stage/muxA/U67  ( .A1(\dp/rf_out1_ex_i [20]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [20]), .B2(
        \dp/ex_stage/muxA/n10 ), .ZN(\dp/ex_stage/muxA/n91 ) );
  INV_X1 \dp/ex_stage/muxA/U66  ( .A(\dp/ex_stage/muxA/n91 ), .ZN(
        \dp/ex_stage/muxA_out [20]) );
  AOI22_X1 \dp/ex_stage/muxA/U65  ( .A1(\dp/rf_out1_ex_i [19]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [19]), .B2(
        \dp/ex_stage/muxA/n11 ), .ZN(\dp/ex_stage/muxA/n89 ) );
  INV_X1 \dp/ex_stage/muxA/U64  ( .A(\dp/ex_stage/muxA/n89 ), .ZN(
        \dp/ex_stage/muxA_out [19]) );
  AOI22_X1 \dp/ex_stage/muxA/U63  ( .A1(\dp/rf_out1_ex_i [30]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [30]), .B2(
        \dp/ex_stage/muxA/n10 ), .ZN(\dp/ex_stage/muxA/n102 ) );
  AOI22_X1 \dp/ex_stage/muxA/U62  ( .A1(\dp/rf_out1_ex_i [18]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [18]), .B2(
        \dp/ex_stage/muxA/n11 ), .ZN(\dp/ex_stage/muxA/n88 ) );
  AOI22_X1 \dp/ex_stage/muxA/U61  ( .A1(\dp/rf_out1_ex_i [26]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [26]), .B2(
        \dp/ex_stage/muxA/n8 ), .ZN(\dp/ex_stage/muxA/n97 ) );
  AOI22_X1 \dp/ex_stage/muxA/U60  ( .A1(\dp/rf_out1_ex_i [25]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [25]), .B2(
        \dp/ex_stage/muxA/n9 ), .ZN(\dp/ex_stage/muxA/n96 ) );
  AOI22_X1 \dp/ex_stage/muxA/U59  ( .A1(\dp/rf_out1_ex_i [24]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [24]), .B2(
        \dp/ex_stage/muxA/n9 ), .ZN(\dp/ex_stage/muxA/n95 ) );
  AOI22_X1 \dp/ex_stage/muxA/U58  ( .A1(\dp/rf_out1_ex_i [28]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [28]), .B2(
        \dp/ex_stage/muxA/n8 ), .ZN(\dp/ex_stage/muxA/n99 ) );
  AOI22_X1 \dp/ex_stage/muxA/U57  ( .A1(\dp/rf_out1_ex_i [27]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [27]), .B2(
        \dp/ex_stage/muxA/n8 ), .ZN(\dp/ex_stage/muxA/n98 ) );
  BUF_X1 \dp/ex_stage/muxA/U56  ( .A(muxA_sel_i), .Z(\dp/ex_stage/muxA/n2 ) );
  BUF_X1 \dp/ex_stage/muxA/U55  ( .A(muxA_sel_i), .Z(\dp/ex_stage/muxA/n3 ) );
  BUF_X1 \dp/ex_stage/muxA/U54  ( .A(muxA_sel_i), .Z(\dp/ex_stage/muxA/n1 ) );
  AOI22_X1 \dp/ex_stage/muxA/U53  ( .A1(\dp/rf_out1_ex_i [1]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [1]), .B2(
        \dp/ex_stage/muxA/n10 ), .ZN(\dp/ex_stage/muxA/n90 ) );
  INV_X1 \dp/ex_stage/muxA/U52  ( .A(\dp/ex_stage/muxA/n90 ), .ZN(
        \dp/ex_stage/muxA_out [1]) );
  AOI22_X1 \dp/ex_stage/muxA/U51  ( .A1(\dp/rf_out1_ex_i [12]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [12]), .B2(
        \dp/ex_stage/muxA/n12 ), .ZN(\dp/ex_stage/muxA/n82 ) );
  INV_X1 \dp/ex_stage/muxA/U50  ( .A(\dp/ex_stage/muxA/n82 ), .ZN(
        \dp/ex_stage/muxA_out [12]) );
  AOI22_X1 \dp/ex_stage/muxA/U49  ( .A1(\dp/rf_out1_ex_i [14]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [14]), .B2(
        \dp/ex_stage/muxA/n12 ), .ZN(\dp/ex_stage/muxA/n84 ) );
  INV_X1 \dp/ex_stage/muxA/U48  ( .A(\dp/ex_stage/muxA/n84 ), .ZN(
        \dp/ex_stage/muxA_out [14]) );
  AOI22_X1 \dp/ex_stage/muxA/U47  ( .A1(\dp/rf_out1_ex_i [15]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [15]), .B2(
        \dp/ex_stage/muxA/n12 ), .ZN(\dp/ex_stage/muxA/n85 ) );
  INV_X1 \dp/ex_stage/muxA/U46  ( .A(\dp/ex_stage/muxA/n85 ), .ZN(
        \dp/ex_stage/muxA_out [15]) );
  AOI22_X1 \dp/ex_stage/muxA/U45  ( .A1(\dp/rf_out1_ex_i [16]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [16]), .B2(
        \dp/ex_stage/muxA/n11 ), .ZN(\dp/ex_stage/muxA/n86 ) );
  INV_X1 \dp/ex_stage/muxA/U44  ( .A(\dp/ex_stage/muxA/n86 ), .ZN(
        \dp/ex_stage/muxA_out [16]) );
  AOI22_X1 \dp/ex_stage/muxA/U43  ( .A1(\dp/rf_out1_ex_i [13]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [13]), .B2(
        \dp/ex_stage/muxA/n12 ), .ZN(\dp/ex_stage/muxA/n83 ) );
  INV_X1 \dp/ex_stage/muxA/U42  ( .A(\dp/ex_stage/muxA/n83 ), .ZN(
        \dp/ex_stage/muxA_out [13]) );
  AOI22_X1 \dp/ex_stage/muxA/U41  ( .A1(\dp/rf_out1_ex_i [5]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [5]), .B2(
        \dp/ex_stage/muxA/n6 ), .ZN(\dp/ex_stage/muxA/n106 ) );
  INV_X1 \dp/ex_stage/muxA/U40  ( .A(\dp/ex_stage/muxA/n106 ), .ZN(
        \dp/ex_stage/muxA_out [5]) );
  AOI22_X1 \dp/ex_stage/muxA/U39  ( .A1(\dp/rf_out1_ex_i [6]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [6]), .B2(
        \dp/ex_stage/muxA/n6 ), .ZN(\dp/ex_stage/muxA/n107 ) );
  AOI22_X1 \dp/ex_stage/muxA/U38  ( .A1(\dp/rf_out1_ex_i [4]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [4]), .B2(
        \dp/ex_stage/muxA/n7 ), .ZN(\dp/ex_stage/muxA/n105 ) );
  AOI22_X1 \dp/ex_stage/muxA/U37  ( .A1(\dp/rf_out1_ex_i [0]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [0]), .B2(
        \dp/ex_stage/muxA/n13 ), .ZN(\dp/ex_stage/muxA/n79 ) );
  AOI22_X1 \dp/ex_stage/muxA/U36  ( .A1(\dp/rf_out1_ex_i [3]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [3]), .B2(
        \dp/ex_stage/muxA/n7 ), .ZN(\dp/ex_stage/muxA/n104 ) );
  AOI22_X1 \dp/ex_stage/muxA/U35  ( .A1(\dp/rf_out1_ex_i [9]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/ex_stage/muxA/n13 ), .B2(
        \dp/npc_ex_i [9]), .ZN(\dp/ex_stage/muxA/n110 ) );
  AOI22_X1 \dp/ex_stage/muxA/U34  ( .A1(\dp/rf_out1_ex_i [2]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [2]), .B2(
        \dp/ex_stage/muxA/n7 ), .ZN(\dp/ex_stage/muxA/n101 ) );
  AOI22_X1 \dp/ex_stage/muxA/U33  ( .A1(\dp/rf_out1_ex_i [7]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [7]), .B2(
        \dp/ex_stage/muxA/n6 ), .ZN(\dp/ex_stage/muxA/n108 ) );
  AOI22_X1 \dp/ex_stage/muxA/U32  ( .A1(\dp/rf_out1_ex_i [8]), .A2(
        \dp/ex_stage/muxA/n5 ), .B1(\dp/npc_ex_i [8]), .B2(
        \dp/ex_stage/muxA/n6 ), .ZN(\dp/ex_stage/muxA/n109 ) );
  AOI22_X1 \dp/ex_stage/muxA/U31  ( .A1(\dp/rf_out1_ex_i [10]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [10]), .B2(
        \dp/ex_stage/muxA/n13 ), .ZN(\dp/ex_stage/muxA/n80 ) );
  AOI22_X1 \dp/ex_stage/muxA/U30  ( .A1(\dp/rf_out1_ex_i [11]), .A2(
        \dp/ex_stage/muxA/n4 ), .B1(\dp/npc_ex_i [11]), .B2(
        \dp/ex_stage/muxA/n13 ), .ZN(\dp/ex_stage/muxA/n81 ) );
  BUF_X1 \dp/ex_stage/muxA/U29  ( .A(\dp/ex_stage/muxA/n2 ), .Z(
        \dp/ex_stage/muxA/n11 ) );
  BUF_X1 \dp/ex_stage/muxA/U28  ( .A(\dp/ex_stage/muxA/n2 ), .Z(
        \dp/ex_stage/muxA/n9 ) );
  BUF_X1 \dp/ex_stage/muxA/U27  ( .A(\dp/ex_stage/muxA/n1 ), .Z(
        \dp/ex_stage/muxA/n8 ) );
  BUF_X1 \dp/ex_stage/muxA/U26  ( .A(\dp/ex_stage/muxA/n3 ), .Z(
        \dp/ex_stage/muxA/n13 ) );
  BUF_X1 \dp/ex_stage/muxA/U25  ( .A(\dp/ex_stage/muxA/n3 ), .Z(
        \dp/ex_stage/muxA/n14 ) );
  BUF_X1 \dp/ex_stage/muxA/U24  ( .A(\dp/ex_stage/muxA/n3 ), .Z(
        \dp/ex_stage/muxA/n12 ) );
  BUF_X1 \dp/ex_stage/muxA/U23  ( .A(\dp/ex_stage/muxA/n2 ), .Z(
        \dp/ex_stage/muxA/n10 ) );
  BUF_X1 \dp/ex_stage/muxA/U22  ( .A(\dp/ex_stage/muxA/n1 ), .Z(
        \dp/ex_stage/muxA/n7 ) );
  BUF_X1 \dp/ex_stage/muxA/U21  ( .A(\dp/ex_stage/muxA/n1 ), .Z(
        \dp/ex_stage/muxA/n6 ) );
  INV_X1 \dp/ex_stage/muxA/U20  ( .A(\dp/ex_stage/muxA/n14 ), .ZN(
        \dp/ex_stage/muxA/n4 ) );
  INV_X1 \dp/ex_stage/muxA/U19  ( .A(\dp/ex_stage/muxA/n14 ), .ZN(
        \dp/ex_stage/muxA/n5 ) );
  INV_X1 \dp/ex_stage/muxA/U18  ( .A(\dp/ex_stage/muxA/n81 ), .ZN(
        \dp/ex_stage/muxA_out [11]) );
  INV_X1 \dp/ex_stage/muxA/U17  ( .A(\dp/ex_stage/muxA/n80 ), .ZN(
        \dp/ex_stage/muxA_out [10]) );
  INV_X1 \dp/ex_stage/muxA/U16  ( .A(\dp/ex_stage/muxA/n88 ), .ZN(
        \dp/ex_stage/muxA_out [18]) );
  INV_X1 \dp/ex_stage/muxA/U15  ( .A(\dp/ex_stage/muxA/n108 ), .ZN(
        \dp/ex_stage/muxA_out [7]) );
  INV_X1 \dp/ex_stage/muxA/U14  ( .A(\dp/ex_stage/muxA/n102 ), .ZN(
        \dp/ex_stage/muxA_out [30]) );
  INV_X1 \dp/ex_stage/muxA/U13  ( .A(\dp/ex_stage/muxA/n100 ), .ZN(
        \dp/ex_stage/muxA_out [29]) );
  INV_X1 \dp/ex_stage/muxA/U12  ( .A(\dp/ex_stage/muxA/n99 ), .ZN(
        \dp/ex_stage/muxA_out [28]) );
  INV_X1 \dp/ex_stage/muxA/U11  ( .A(\dp/ex_stage/muxA/n98 ), .ZN(
        \dp/ex_stage/muxA_out [27]) );
  INV_X1 \dp/ex_stage/muxA/U10  ( .A(\dp/ex_stage/muxA/n97 ), .ZN(
        \dp/ex_stage/muxA_out [26]) );
  INV_X1 \dp/ex_stage/muxA/U9  ( .A(\dp/ex_stage/muxA/n96 ), .ZN(
        \dp/ex_stage/muxA_out [25]) );
  INV_X1 \dp/ex_stage/muxA/U8  ( .A(\dp/ex_stage/muxA/n95 ), .ZN(
        \dp/ex_stage/muxA_out [24]) );
  INV_X1 \dp/ex_stage/muxA/U7  ( .A(\dp/ex_stage/muxA/n110 ), .ZN(
        \dp/ex_stage/muxA_out [9]) );
  INV_X1 \dp/ex_stage/muxA/U6  ( .A(\dp/ex_stage/muxA/n109 ), .ZN(
        \dp/ex_stage/muxA_out [8]) );
  INV_X1 \dp/ex_stage/muxA/U5  ( .A(\dp/ex_stage/muxA/n104 ), .ZN(
        \dp/ex_stage/muxA_out [3]) );
  INV_X1 \dp/ex_stage/muxA/U4  ( .A(\dp/ex_stage/muxA/n101 ), .ZN(
        \dp/ex_stage/muxA_out [2]) );
  INV_X1 \dp/ex_stage/muxA/U3  ( .A(\dp/ex_stage/muxA/n107 ), .ZN(
        \dp/ex_stage/muxA_out [6]) );
  INV_X1 \dp/ex_stage/muxA/U2  ( .A(\dp/ex_stage/muxA/n105 ), .ZN(
        \dp/ex_stage/muxA_out [4]) );
  INV_X1 \dp/ex_stage/muxA/U1  ( .A(\dp/ex_stage/muxA/n79 ), .ZN(
        \dp/ex_stage/alu/shifter/N202 ) );
  AOI22_X1 \dp/ex_stage/muxB/U78  ( .A1(\dp/data_mem_ex_o [23]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [23]), .B2(
        \dp/ex_stage/muxB/n9 ), .ZN(\dp/ex_stage/muxB/n94 ) );
  INV_X1 \dp/ex_stage/muxB/U77  ( .A(\dp/ex_stage/muxB/n94 ), .ZN(
        \dp/ex_stage/muxB_out [23]) );
  AOI22_X1 \dp/ex_stage/muxB/U76  ( .A1(\dp/data_mem_ex_o [19]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [19]), .B2(
        \dp/ex_stage/muxB/n11 ), .ZN(\dp/ex_stage/muxB/n89 ) );
  INV_X1 \dp/ex_stage/muxB/U75  ( .A(\dp/ex_stage/muxB/n89 ), .ZN(
        \dp/ex_stage/muxB_out [19]) );
  AOI22_X1 \dp/ex_stage/muxB/U74  ( .A1(\dp/data_mem_ex_o [27]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [27]), .B2(
        \dp/ex_stage/muxB/n8 ), .ZN(\dp/ex_stage/muxB/n98 ) );
  INV_X1 \dp/ex_stage/muxB/U73  ( .A(\dp/ex_stage/muxB/n98 ), .ZN(
        \dp/ex_stage/muxB_out [27]) );
  AOI22_X1 \dp/ex_stage/muxB/U72  ( .A1(\dp/data_mem_ex_o [15]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [15]), .B2(
        \dp/ex_stage/muxB/n12 ), .ZN(\dp/ex_stage/muxB/n85 ) );
  INV_X1 \dp/ex_stage/muxB/U71  ( .A(\dp/ex_stage/muxB/n85 ), .ZN(
        \dp/ex_stage/muxB_out [15]) );
  AOI22_X1 \dp/ex_stage/muxB/U70  ( .A1(\dp/data_mem_ex_o [25]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [25]), .B2(
        \dp/ex_stage/muxB/n9 ), .ZN(\dp/ex_stage/muxB/n96 ) );
  INV_X1 \dp/ex_stage/muxB/U69  ( .A(\dp/ex_stage/muxB/n96 ), .ZN(
        \dp/ex_stage/muxB_out [25]) );
  AOI22_X1 \dp/ex_stage/muxB/U68  ( .A1(\dp/data_mem_ex_o [21]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [21]), .B2(
        \dp/ex_stage/muxB/n10 ), .ZN(\dp/ex_stage/muxB/n92 ) );
  INV_X1 \dp/ex_stage/muxB/U67  ( .A(\dp/ex_stage/muxB/n92 ), .ZN(
        \dp/ex_stage/muxB_out [21]) );
  AOI22_X1 \dp/ex_stage/muxB/U66  ( .A1(\dp/data_mem_ex_o [17]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [17]), .B2(
        \dp/ex_stage/muxB/n11 ), .ZN(\dp/ex_stage/muxB/n87 ) );
  INV_X1 \dp/ex_stage/muxB/U65  ( .A(\dp/ex_stage/muxB/n87 ), .ZN(
        \dp/ex_stage/muxB_out [17]) );
  AOI22_X1 \dp/ex_stage/muxB/U64  ( .A1(\dp/data_mem_ex_o [13]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [13]), .B2(
        \dp/ex_stage/muxB/n12 ), .ZN(\dp/ex_stage/muxB/n83 ) );
  INV_X1 \dp/ex_stage/muxB/U63  ( .A(\dp/ex_stage/muxB/n83 ), .ZN(
        \dp/ex_stage/muxB_out [13]) );
  AOI22_X1 \dp/ex_stage/muxB/U62  ( .A1(\dp/data_mem_ex_o [24]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [24]), .B2(
        \dp/ex_stage/muxB/n9 ), .ZN(\dp/ex_stage/muxB/n95 ) );
  INV_X1 \dp/ex_stage/muxB/U61  ( .A(\dp/ex_stage/muxB/n95 ), .ZN(
        \dp/ex_stage/muxB_out [24]) );
  AOI22_X1 \dp/ex_stage/muxB/U60  ( .A1(\dp/data_mem_ex_o [20]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [20]), .B2(
        \dp/ex_stage/muxB/n10 ), .ZN(\dp/ex_stage/muxB/n91 ) );
  INV_X1 \dp/ex_stage/muxB/U59  ( .A(\dp/ex_stage/muxB/n91 ), .ZN(
        \dp/ex_stage/muxB_out [20]) );
  AOI22_X1 \dp/ex_stage/muxB/U58  ( .A1(\dp/data_mem_ex_o [16]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [16]), .B2(
        \dp/ex_stage/muxB/n11 ), .ZN(\dp/ex_stage/muxB/n86 ) );
  INV_X1 \dp/ex_stage/muxB/U57  ( .A(\dp/ex_stage/muxB/n86 ), .ZN(
        \dp/ex_stage/muxB_out [16]) );
  AOI22_X1 \dp/ex_stage/muxB/U56  ( .A1(\dp/data_mem_ex_o [31]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [31]), .B2(
        \dp/ex_stage/muxB/n7 ), .ZN(\dp/ex_stage/muxB/n103 ) );
  INV_X1 \dp/ex_stage/muxB/U55  ( .A(\dp/ex_stage/muxB/n103 ), .ZN(
        \dp/ex_stage/muxB_out [31]) );
  AOI22_X1 \dp/ex_stage/muxB/U54  ( .A1(\dp/data_mem_ex_o [26]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [26]), .B2(
        \dp/ex_stage/muxB/n8 ), .ZN(\dp/ex_stage/muxB/n97 ) );
  INV_X1 \dp/ex_stage/muxB/U53  ( .A(\dp/ex_stage/muxB/n97 ), .ZN(
        \dp/ex_stage/muxB_out [26]) );
  AOI22_X1 \dp/ex_stage/muxB/U52  ( .A1(\dp/data_mem_ex_o [22]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [22]), .B2(
        \dp/ex_stage/muxB/n9 ), .ZN(\dp/ex_stage/muxB/n93 ) );
  INV_X1 \dp/ex_stage/muxB/U51  ( .A(\dp/ex_stage/muxB/n93 ), .ZN(
        \dp/ex_stage/muxB_out [22]) );
  AOI22_X1 \dp/ex_stage/muxB/U50  ( .A1(\dp/data_mem_ex_o [18]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [18]), .B2(
        \dp/ex_stage/muxB/n11 ), .ZN(\dp/ex_stage/muxB/n88 ) );
  INV_X1 \dp/ex_stage/muxB/U49  ( .A(\dp/ex_stage/muxB/n88 ), .ZN(
        \dp/ex_stage/muxB_out [18]) );
  AOI22_X1 \dp/ex_stage/muxB/U48  ( .A1(\dp/data_mem_ex_o [14]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [14]), .B2(
        \dp/ex_stage/muxB/n12 ), .ZN(\dp/ex_stage/muxB/n84 ) );
  INV_X1 \dp/ex_stage/muxB/U47  ( .A(\dp/ex_stage/muxB/n84 ), .ZN(
        \dp/ex_stage/muxB_out [14]) );
  AOI22_X1 \dp/ex_stage/muxB/U46  ( .A1(\dp/data_mem_ex_o [30]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [30]), .B2(
        \dp/ex_stage/muxB/n10 ), .ZN(\dp/ex_stage/muxB/n102 ) );
  INV_X1 \dp/ex_stage/muxB/U45  ( .A(\dp/ex_stage/muxB/n102 ), .ZN(
        \dp/ex_stage/muxB_out [30]) );
  AOI22_X1 \dp/ex_stage/muxB/U44  ( .A1(\dp/data_mem_ex_o [28]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [28]), .B2(
        \dp/ex_stage/muxB/n8 ), .ZN(\dp/ex_stage/muxB/n99 ) );
  INV_X1 \dp/ex_stage/muxB/U43  ( .A(\dp/ex_stage/muxB/n99 ), .ZN(
        \dp/ex_stage/muxB_out [28]) );
  AOI22_X1 \dp/ex_stage/muxB/U42  ( .A1(\dp/data_mem_ex_o [29]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [29]), .B2(
        \dp/ex_stage/muxB/n8 ), .ZN(\dp/ex_stage/muxB/n100 ) );
  INV_X1 \dp/ex_stage/muxB/U41  ( .A(\dp/ex_stage/muxB/n100 ), .ZN(
        \dp/ex_stage/muxB_out [29]) );
  BUF_X1 \dp/ex_stage/muxB/U40  ( .A(muxB_sel_i), .Z(\dp/ex_stage/muxB/n1 ) );
  BUF_X1 \dp/ex_stage/muxB/U39  ( .A(muxB_sel_i), .Z(\dp/ex_stage/muxB/n2 ) );
  BUF_X1 \dp/ex_stage/muxB/U38  ( .A(muxB_sel_i), .Z(\dp/ex_stage/muxB/n3 ) );
  AOI22_X1 \dp/ex_stage/muxB/U37  ( .A1(\dp/data_mem_ex_o [1]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [1]), .B2(
        \dp/ex_stage/muxB/n10 ), .ZN(\dp/ex_stage/muxB/n90 ) );
  INV_X1 \dp/ex_stage/muxB/U36  ( .A(\dp/ex_stage/muxB/n90 ), .ZN(
        \dp/ex_stage/muxB_out [1]) );
  AOI22_X1 \dp/ex_stage/muxB/U35  ( .A1(\dp/data_mem_ex_o [4]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [4]), .B2(
        \dp/ex_stage/muxB/n7 ), .ZN(\dp/ex_stage/muxB/n105 ) );
  INV_X1 \dp/ex_stage/muxB/U34  ( .A(\dp/ex_stage/muxB/n105 ), .ZN(
        \dp/ex_stage/muxB_out [4]) );
  AOI22_X1 \dp/ex_stage/muxB/U33  ( .A1(\dp/data_mem_ex_o [2]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [2]), .B2(
        \dp/ex_stage/muxB/n7 ), .ZN(\dp/ex_stage/muxB/n101 ) );
  INV_X1 \dp/ex_stage/muxB/U32  ( .A(\dp/ex_stage/muxB/n101 ), .ZN(
        \dp/ex_stage/muxB_out [2]) );
  AOI22_X1 \dp/ex_stage/muxB/U31  ( .A1(\dp/data_mem_ex_o [11]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [11]), .B2(
        \dp/ex_stage/muxB/n13 ), .ZN(\dp/ex_stage/muxB/n81 ) );
  INV_X1 \dp/ex_stage/muxB/U30  ( .A(\dp/ex_stage/muxB/n81 ), .ZN(
        \dp/ex_stage/muxB_out [11]) );
  AOI22_X1 \dp/ex_stage/muxB/U29  ( .A1(\dp/data_mem_ex_o [12]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [12]), .B2(
        \dp/ex_stage/muxB/n12 ), .ZN(\dp/ex_stage/muxB/n82 ) );
  INV_X1 \dp/ex_stage/muxB/U28  ( .A(\dp/ex_stage/muxB/n82 ), .ZN(
        \dp/ex_stage/muxB_out [12]) );
  AOI22_X1 \dp/ex_stage/muxB/U27  ( .A1(\dp/data_mem_ex_o [5]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [5]), .B2(
        \dp/ex_stage/muxB/n6 ), .ZN(\dp/ex_stage/muxB/n106 ) );
  INV_X1 \dp/ex_stage/muxB/U26  ( .A(\dp/ex_stage/muxB/n106 ), .ZN(
        \dp/ex_stage/muxB_out [5]) );
  AOI22_X1 \dp/ex_stage/muxB/U25  ( .A1(\dp/data_mem_ex_o [9]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/ex_stage/muxB/n13 ), .B2(
        \dp/imm_ex_i [9]), .ZN(\dp/ex_stage/muxB/n110 ) );
  INV_X1 \dp/ex_stage/muxB/U24  ( .A(\dp/ex_stage/muxB/n110 ), .ZN(
        \dp/ex_stage/muxB_out [9]) );
  AOI22_X1 \dp/ex_stage/muxB/U23  ( .A1(\dp/data_mem_ex_o [8]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [8]), .B2(
        \dp/ex_stage/muxB/n6 ), .ZN(\dp/ex_stage/muxB/n109 ) );
  INV_X1 \dp/ex_stage/muxB/U22  ( .A(\dp/ex_stage/muxB/n109 ), .ZN(
        \dp/ex_stage/muxB_out [8]) );
  AOI22_X1 \dp/ex_stage/muxB/U21  ( .A1(\dp/data_mem_ex_o [10]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [10]), .B2(
        \dp/ex_stage/muxB/n13 ), .ZN(\dp/ex_stage/muxB/n80 ) );
  INV_X1 \dp/ex_stage/muxB/U20  ( .A(\dp/ex_stage/muxB/n80 ), .ZN(
        \dp/ex_stage/muxB_out [10]) );
  AOI22_X1 \dp/ex_stage/muxB/U19  ( .A1(\dp/data_mem_ex_o [6]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [6]), .B2(
        \dp/ex_stage/muxB/n6 ), .ZN(\dp/ex_stage/muxB/n107 ) );
  INV_X1 \dp/ex_stage/muxB/U18  ( .A(\dp/ex_stage/muxB/n107 ), .ZN(
        \dp/ex_stage/muxB_out [6]) );
  AOI22_X1 \dp/ex_stage/muxB/U17  ( .A1(\dp/data_mem_ex_o [3]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [3]), .B2(
        \dp/ex_stage/muxB/n7 ), .ZN(\dp/ex_stage/muxB/n104 ) );
  INV_X1 \dp/ex_stage/muxB/U16  ( .A(\dp/ex_stage/muxB/n104 ), .ZN(
        \dp/ex_stage/muxB_out [3]) );
  AOI22_X1 \dp/ex_stage/muxB/U15  ( .A1(\dp/data_mem_ex_o [7]), .A2(
        \dp/ex_stage/muxB/n5 ), .B1(\dp/imm_ex_i [7]), .B2(
        \dp/ex_stage/muxB/n6 ), .ZN(\dp/ex_stage/muxB/n108 ) );
  INV_X1 \dp/ex_stage/muxB/U14  ( .A(\dp/ex_stage/muxB/n108 ), .ZN(
        \dp/ex_stage/muxB_out [7]) );
  AOI22_X1 \dp/ex_stage/muxB/U13  ( .A1(\dp/data_mem_ex_o [0]), .A2(
        \dp/ex_stage/muxB/n4 ), .B1(\dp/imm_ex_i [0]), .B2(
        \dp/ex_stage/muxB/n13 ), .ZN(\dp/ex_stage/muxB/n79 ) );
  INV_X1 \dp/ex_stage/muxB/U12  ( .A(\dp/ex_stage/muxB/n79 ), .ZN(
        \dp/ex_stage/muxB_out [0]) );
  BUF_X1 \dp/ex_stage/muxB/U11  ( .A(\dp/ex_stage/muxB/n1 ), .Z(
        \dp/ex_stage/muxB/n8 ) );
  BUF_X1 \dp/ex_stage/muxB/U10  ( .A(\dp/ex_stage/muxB/n2 ), .Z(
        \dp/ex_stage/muxB/n9 ) );
  BUF_X1 \dp/ex_stage/muxB/U9  ( .A(\dp/ex_stage/muxB/n2 ), .Z(
        \dp/ex_stage/muxB/n11 ) );
  BUF_X1 \dp/ex_stage/muxB/U8  ( .A(\dp/ex_stage/muxB/n3 ), .Z(
        \dp/ex_stage/muxB/n12 ) );
  BUF_X1 \dp/ex_stage/muxB/U7  ( .A(\dp/ex_stage/muxB/n3 ), .Z(
        \dp/ex_stage/muxB/n13 ) );
  BUF_X1 \dp/ex_stage/muxB/U6  ( .A(\dp/ex_stage/muxB/n3 ), .Z(
        \dp/ex_stage/muxB/n14 ) );
  BUF_X1 \dp/ex_stage/muxB/U5  ( .A(\dp/ex_stage/muxB/n1 ), .Z(
        \dp/ex_stage/muxB/n7 ) );
  BUF_X1 \dp/ex_stage/muxB/U4  ( .A(\dp/ex_stage/muxB/n2 ), .Z(
        \dp/ex_stage/muxB/n10 ) );
  BUF_X1 \dp/ex_stage/muxB/U3  ( .A(\dp/ex_stage/muxB/n1 ), .Z(
        \dp/ex_stage/muxB/n6 ) );
  INV_X1 \dp/ex_stage/muxB/U2  ( .A(\dp/ex_stage/muxB/n14 ), .ZN(
        \dp/ex_stage/muxB/n4 ) );
  INV_X1 \dp/ex_stage/muxB/U1  ( .A(\dp/ex_stage/muxB/n14 ), .ZN(
        \dp/ex_stage/muxB/n5 ) );
  INV_X1 \dp/ex_stage/alu/U263  ( .A(\dp/ex_stage/alu/n46 ), .ZN(
        \dp/ex_stage/alu/n45 ) );
  INV_X1 \dp/ex_stage/alu/U262  ( .A(\dp/ex_stage/alu/n38 ), .ZN(
        \dp/ex_stage/alu/n37 ) );
  INV_X1 \dp/ex_stage/alu/U261  ( .A(\dp/ex_stage/alu/n35 ), .ZN(
        \dp/ex_stage/alu/n34 ) );
  INV_X1 \dp/ex_stage/alu/U260  ( .A(\dp/ex_stage/alu/n32 ), .ZN(
        \dp/ex_stage/alu/n31 ) );
  INV_X2 \dp/ex_stage/alu/U259  ( .A(\dp/ex_stage/alu/n30 ), .ZN(
        \dp/ex_stage/alu/n29 ) );
  INV_X1 \dp/ex_stage/alu/U258  ( .A(\dp/ex_stage/alu/n26 ), .ZN(
        \dp/ex_stage/alu/n25 ) );
  CLKBUF_X1 \dp/ex_stage/alu/U257  ( .A(\dp/ex_stage/alu/n221 ), .Z(
        \dp/ex_stage/alu/n18 ) );
  OAI21_X1 \dp/ex_stage/alu/U256  ( .B1(\dp/ex_stage/alu/n93 ), .B2(
        \dp/ex_stage/alu/n223 ), .A(alu_op_i[4]), .ZN(\dp/ex_stage/alu/n207 )
         );
  NOR3_X1 \dp/ex_stage/alu/U255  ( .A1(alu_op_i[1]), .A2(alu_op_i[4]), .A3(
        \dp/ex_stage/alu/n227 ), .ZN(\dp/ex_stage/alu/n205 ) );
  INV_X1 \dp/ex_stage/alu/U254  ( .A(\dp/ex_stage/muxA_out [17]), .ZN(
        \dp/ex_stage/alu/n41 ) );
  INV_X1 \dp/ex_stage/alu/U253  ( .A(\dp/ex_stage/muxA_out [21]), .ZN(
        \dp/ex_stage/alu/n42 ) );
  INV_X1 \dp/ex_stage/alu/U252  ( .A(\dp/ex_stage/muxA_out [23]), .ZN(
        \dp/ex_stage/alu/n46 ) );
  INV_X1 \dp/ex_stage/alu/U251  ( .A(\dp/ex_stage/muxA_out [22]), .ZN(
        \dp/ex_stage/alu/n44 ) );
  NAND2_X1 \dp/ex_stage/alu/U250  ( .A1(alu_op_i[4]), .A2(
        \dp/ex_stage/alu/n88 ), .ZN(\dp/ex_stage/alu/shift_arith_i ) );
  INV_X1 \dp/ex_stage/alu/U249  ( .A(alu_op_i[2]), .ZN(\dp/ex_stage/alu/n224 )
         );
  INV_X1 \dp/ex_stage/alu/U248  ( .A(alu_op_i[4]), .ZN(\dp/ex_stage/alu/n219 )
         );
  INV_X1 \dp/ex_stage/alu/U247  ( .A(alu_op_i[3]), .ZN(\dp/ex_stage/alu/n222 )
         );
  OAI21_X1 \dp/ex_stage/alu/U246  ( .B1(\dp/ex_stage/alu/n90 ), .B2(
        \dp/ex_stage/alu/n222 ), .A(\dp/ex_stage/alu/n91 ), .ZN(
        \dp/ex_stage/alu/N23 ) );
  AOI21_X1 \dp/ex_stage/alu/U245  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n214 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n128 ) );
  OAI221_X1 \dp/ex_stage/alu/U244  ( .B1(\dp/ex_stage/alu/n128 ), .B2(
        \dp/ex_stage/alu/n66 ), .C1(\dp/ex_stage/alu/n129 ), .C2(
        \dp/ex_stage/alu/n214 ), .A(\dp/ex_stage/alu/n130 ), .ZN(
        \dp/alu_out_ex_o [28]) );
  AOI21_X1 \dp/ex_stage/alu/U243  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n215 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n125 ) );
  OAI221_X1 \dp/ex_stage/alu/U242  ( .B1(\dp/ex_stage/alu/n125 ), .B2(
        \dp/ex_stage/alu/n67 ), .C1(\dp/ex_stage/alu/n126 ), .C2(
        \dp/ex_stage/alu/n215 ), .A(\dp/ex_stage/alu/n127 ), .ZN(
        \dp/alu_out_ex_o [29]) );
  AOI21_X1 \dp/ex_stage/alu/U241  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n216 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n119 ) );
  OAI221_X1 \dp/ex_stage/alu/U240  ( .B1(\dp/ex_stage/alu/n119 ), .B2(
        \dp/ex_stage/alu/n68 ), .C1(\dp/ex_stage/alu/n120 ), .C2(
        \dp/ex_stage/alu/n216 ), .A(\dp/ex_stage/alu/n121 ), .ZN(
        \dp/alu_out_ex_o [30]) );
  AOI21_X1 \dp/ex_stage/alu/U239  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n217 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n116 ) );
  OAI221_X1 \dp/ex_stage/alu/U238  ( .B1(\dp/ex_stage/alu/n116 ), .B2(
        \dp/ex_stage/alu/n69 ), .C1(\dp/ex_stage/alu/n117 ), .C2(
        \dp/ex_stage/alu/n217 ), .A(\dp/ex_stage/alu/n118 ), .ZN(
        \dp/alu_out_ex_o [31]) );
  AOI21_X1 \dp/ex_stage/alu/U237  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n70 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n107 ) );
  OAI221_X1 \dp/ex_stage/alu/U236  ( .B1(\dp/ex_stage/alu/n107 ), .B2(
        \dp/ex_stage/alu/n52 ), .C1(\dp/ex_stage/alu/n108 ), .C2(
        \dp/ex_stage/alu/n70 ), .A(\dp/ex_stage/alu/n109 ), .ZN(
        \dp/alu_out_ex_o [5]) );
  AOI21_X1 \dp/ex_stage/alu/U229  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n71 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n104 ) );
  OAI221_X1 \dp/ex_stage/alu/U228  ( .B1(\dp/ex_stage/alu/n104 ), .B2(
        \dp/ex_stage/alu/n53 ), .C1(\dp/ex_stage/alu/n105 ), .C2(
        \dp/ex_stage/alu/n71 ), .A(\dp/ex_stage/alu/n106 ), .ZN(
        \dp/alu_out_ex_o [6]) );
  AOI21_X1 \dp/ex_stage/alu/U227  ( .B1(\dp/ex_stage/alu/n18 ), .B2(
        \dp/ex_stage/alu/n72 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n101 ) );
  OAI221_X1 \dp/ex_stage/alu/U226  ( .B1(\dp/ex_stage/alu/n101 ), .B2(
        \dp/ex_stage/alu/n54 ), .C1(\dp/ex_stage/alu/n102 ), .C2(
        \dp/ex_stage/alu/n72 ), .A(\dp/ex_stage/alu/n103 ), .ZN(
        \dp/alu_out_ex_o [7]) );
  AOI21_X1 \dp/ex_stage/alu/U225  ( .B1(\dp/ex_stage/alu/n18 ), .B2(
        \dp/ex_stage/alu/n73 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n98 ) );
  OAI221_X1 \dp/ex_stage/alu/U224  ( .B1(\dp/ex_stage/alu/n98 ), .B2(
        \dp/ex_stage/alu/n55 ), .C1(\dp/ex_stage/alu/n99 ), .C2(
        \dp/ex_stage/alu/n73 ), .A(\dp/ex_stage/alu/n100 ), .ZN(
        \dp/alu_out_ex_o [8]) );
  AOI21_X1 \dp/ex_stage/alu/U223  ( .B1(\dp/ex_stage/alu/n18 ), .B2(
        \dp/ex_stage/alu/n74 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n94 ) );
  OAI221_X1 \dp/ex_stage/alu/U222  ( .B1(\dp/ex_stage/alu/n94 ), .B2(
        \dp/ex_stage/alu/n56 ), .C1(\dp/ex_stage/alu/n95 ), .C2(
        \dp/ex_stage/alu/n74 ), .A(\dp/ex_stage/alu/n96 ), .ZN(
        \dp/alu_out_ex_o [9]) );
  AOI21_X1 \dp/ex_stage/alu/U221  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n77 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n179 ) );
  OAI221_X1 \dp/ex_stage/alu/U220  ( .B1(\dp/ex_stage/alu/n179 ), .B2(
        \dp/ex_stage/alu/n35 ), .C1(\dp/ex_stage/alu/n180 ), .C2(
        \dp/ex_stage/alu/n77 ), .A(\dp/ex_stage/alu/n181 ), .ZN(
        \dp/alu_out_ex_o [12]) );
  AOI21_X1 \dp/ex_stage/alu/U219  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n82 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n164 ) );
  OAI221_X1 \dp/ex_stage/alu/U218  ( .B1(\dp/ex_stage/alu/n164 ), .B2(
        \dp/ex_stage/alu/n41 ), .C1(\dp/ex_stage/alu/n165 ), .C2(
        \dp/ex_stage/alu/n82 ), .A(\dp/ex_stage/alu/n166 ), .ZN(
        \dp/alu_out_ex_o [17]) );
  AOI21_X1 \dp/ex_stage/alu/U217  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n83 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n161 ) );
  OAI221_X1 \dp/ex_stage/alu/U216  ( .B1(\dp/ex_stage/alu/n161 ), .B2(
        \dp/ex_stage/alu/n59 ), .C1(\dp/ex_stage/alu/n162 ), .C2(
        \dp/ex_stage/alu/n83 ), .A(\dp/ex_stage/alu/n163 ), .ZN(
        \dp/alu_out_ex_o [18]) );
  AOI21_X1 \dp/ex_stage/alu/U215  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n84 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n158 ) );
  OAI221_X1 \dp/ex_stage/alu/U214  ( .B1(\dp/ex_stage/alu/n158 ), .B2(
        \dp/ex_stage/alu/n60 ), .C1(\dp/ex_stage/alu/n159 ), .C2(
        \dp/ex_stage/alu/n84 ), .A(\dp/ex_stage/alu/n160 ), .ZN(
        \dp/alu_out_ex_o [19]) );
  AOI21_X1 \dp/ex_stage/alu/U213  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n85 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n152 ) );
  OAI221_X1 \dp/ex_stage/alu/U212  ( .B1(\dp/ex_stage/alu/n152 ), .B2(
        \dp/ex_stage/alu/n61 ), .C1(\dp/ex_stage/alu/n153 ), .C2(
        \dp/ex_stage/alu/n85 ), .A(\dp/ex_stage/alu/n154 ), .ZN(
        \dp/alu_out_ex_o [20]) );
  AOI21_X1 \dp/ex_stage/alu/U211  ( .B1(\dp/ex_stage/alu/n15 ), .B2(
        \dp/ex_stage/alu/n86 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n149 ) );
  OAI221_X1 \dp/ex_stage/alu/U210  ( .B1(\dp/ex_stage/alu/n149 ), .B2(
        \dp/ex_stage/alu/n42 ), .C1(\dp/ex_stage/alu/n150 ), .C2(
        \dp/ex_stage/alu/n86 ), .A(\dp/ex_stage/alu/n151 ), .ZN(
        \dp/alu_out_ex_o [21]) );
  AOI21_X1 \dp/ex_stage/alu/U209  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n87 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n146 ) );
  OAI221_X1 \dp/ex_stage/alu/U208  ( .B1(\dp/ex_stage/alu/n146 ), .B2(
        \dp/ex_stage/alu/n44 ), .C1(\dp/ex_stage/alu/n147 ), .C2(
        \dp/ex_stage/alu/n87 ), .A(\dp/ex_stage/alu/n148 ), .ZN(
        \dp/alu_out_ex_o [22]) );
  AOI21_X1 \dp/ex_stage/alu/U207  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n209 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n143 ) );
  OAI221_X1 \dp/ex_stage/alu/U206  ( .B1(\dp/ex_stage/alu/n143 ), .B2(
        \dp/ex_stage/alu/n46 ), .C1(\dp/ex_stage/alu/n144 ), .C2(
        \dp/ex_stage/alu/n209 ), .A(\dp/ex_stage/alu/n145 ), .ZN(
        \dp/alu_out_ex_o [23]) );
  AOI21_X1 \dp/ex_stage/alu/U205  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n210 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n140 ) );
  OAI221_X1 \dp/ex_stage/alu/U204  ( .B1(\dp/ex_stage/alu/n140 ), .B2(
        \dp/ex_stage/alu/n62 ), .C1(\dp/ex_stage/alu/n141 ), .C2(
        \dp/ex_stage/alu/n210 ), .A(\dp/ex_stage/alu/n142 ), .ZN(
        \dp/alu_out_ex_o [24]) );
  AOI21_X1 \dp/ex_stage/alu/U203  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n211 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n137 ) );
  OAI221_X1 \dp/ex_stage/alu/U202  ( .B1(\dp/ex_stage/alu/n137 ), .B2(
        \dp/ex_stage/alu/n63 ), .C1(\dp/ex_stage/alu/n138 ), .C2(
        \dp/ex_stage/alu/n211 ), .A(\dp/ex_stage/alu/n139 ), .ZN(
        \dp/alu_out_ex_o [25]) );
  AOI21_X1 \dp/ex_stage/alu/U201  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n212 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n134 ) );
  OAI221_X1 \dp/ex_stage/alu/U200  ( .B1(\dp/ex_stage/alu/n134 ), .B2(
        \dp/ex_stage/alu/n64 ), .C1(\dp/ex_stage/alu/n135 ), .C2(
        \dp/ex_stage/alu/n212 ), .A(\dp/ex_stage/alu/n136 ), .ZN(
        \dp/alu_out_ex_o [26]) );
  AOI21_X1 \dp/ex_stage/alu/U199  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n213 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n131 ) );
  OAI221_X1 \dp/ex_stage/alu/U198  ( .B1(\dp/ex_stage/alu/n131 ), .B2(
        \dp/ex_stage/alu/n65 ), .C1(\dp/ex_stage/alu/n132 ), .C2(
        \dp/ex_stage/alu/n213 ), .A(\dp/ex_stage/alu/n133 ), .ZN(
        \dp/alu_out_ex_o [27]) );
  AOI21_X1 \dp/ex_stage/alu/U197  ( .B1(\dp/ex_stage/alu/n15 ), .B2(
        \dp/ex_stage/alu/n26 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n155 ) );
  OAI221_X1 \dp/ex_stage/alu/U196  ( .B1(\dp/ex_stage/alu/n155 ), .B2(
        \dp/ex_stage/alu/n33 ), .C1(\dp/ex_stage/alu/n156 ), .C2(
        \dp/ex_stage/alu/n26 ), .A(\dp/ex_stage/alu/n157 ), .ZN(
        \dp/alu_out_ex_o [1]) );
  AOI21_X1 \dp/ex_stage/alu/U195  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n28 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n122 ) );
  OAI221_X1 \dp/ex_stage/alu/U194  ( .B1(\dp/ex_stage/alu/n122 ), .B2(
        \dp/ex_stage/alu/n49 ), .C1(\dp/ex_stage/alu/n123 ), .C2(
        \dp/ex_stage/alu/n28 ), .A(\dp/ex_stage/alu/n124 ), .ZN(
        \dp/alu_out_ex_o [2]) );
  AOI21_X1 \dp/ex_stage/alu/U193  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n30 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n113 ) );
  OAI221_X1 \dp/ex_stage/alu/U192  ( .B1(\dp/ex_stage/alu/n113 ), .B2(
        \dp/ex_stage/alu/n50 ), .C1(\dp/ex_stage/alu/n114 ), .C2(
        \dp/ex_stage/alu/n30 ), .A(\dp/ex_stage/alu/n115 ), .ZN(
        \dp/alu_out_ex_o [3]) );
  AOI21_X1 \dp/ex_stage/alu/U191  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n32 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n110 ) );
  OAI221_X1 \dp/ex_stage/alu/U190  ( .B1(\dp/ex_stage/alu/n110 ), .B2(
        \dp/ex_stage/alu/n51 ), .C1(\dp/ex_stage/alu/n111 ), .C2(
        \dp/ex_stage/alu/n32 ), .A(\dp/ex_stage/alu/n112 ), .ZN(
        \dp/alu_out_ex_o [4]) );
  INV_X1 \dp/ex_stage/alu/U189  ( .A(alu_op_i[0]), .ZN(\dp/ex_stage/alu/n227 )
         );
  INV_X1 \dp/ex_stage/alu/U188  ( .A(alu_op_i[1]), .ZN(\dp/ex_stage/alu/n226 )
         );
  NOR2_X1 \dp/ex_stage/alu/U187  ( .A1(alu_op_i[3]), .A2(alu_op_i[2]), .ZN(
        \dp/ex_stage/alu/n92 ) );
  AOI21_X1 \dp/ex_stage/alu/U186  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n78 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n176 ) );
  OAI221_X1 \dp/ex_stage/alu/U185  ( .B1(\dp/ex_stage/alu/n176 ), .B2(
        \dp/ex_stage/alu/n36 ), .C1(\dp/ex_stage/alu/n177 ), .C2(
        \dp/ex_stage/alu/n78 ), .A(\dp/ex_stage/alu/n178 ), .ZN(
        \dp/alu_out_ex_o [13]) );
  AOI21_X1 \dp/ex_stage/alu/U184  ( .B1(\dp/ex_stage/alu/n17 ), .B2(
        \dp/ex_stage/alu/n79 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n173 ) );
  OAI221_X1 \dp/ex_stage/alu/U183  ( .B1(\dp/ex_stage/alu/n173 ), .B2(
        \dp/ex_stage/alu/n38 ), .C1(\dp/ex_stage/alu/n174 ), .C2(
        \dp/ex_stage/alu/n79 ), .A(\dp/ex_stage/alu/n175 ), .ZN(
        \dp/alu_out_ex_o [14]) );
  AOI21_X1 \dp/ex_stage/alu/U182  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n80 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n170 ) );
  OAI221_X1 \dp/ex_stage/alu/U181  ( .B1(\dp/ex_stage/alu/n170 ), .B2(
        \dp/ex_stage/alu/n39 ), .C1(\dp/ex_stage/alu/n171 ), .C2(
        \dp/ex_stage/alu/n80 ), .A(\dp/ex_stage/alu/n172 ), .ZN(
        \dp/alu_out_ex_o [15]) );
  AOI21_X1 \dp/ex_stage/alu/U180  ( .B1(\dp/ex_stage/alu/n16 ), .B2(
        \dp/ex_stage/alu/n81 ), .A(\dp/ex_stage/alu/n6 ), .ZN(
        \dp/ex_stage/alu/n167 ) );
  OAI221_X1 \dp/ex_stage/alu/U179  ( .B1(\dp/ex_stage/alu/n167 ), .B2(
        \dp/ex_stage/alu/n40 ), .C1(\dp/ex_stage/alu/n168 ), .C2(
        \dp/ex_stage/alu/n81 ), .A(\dp/ex_stage/alu/n169 ), .ZN(
        \dp/alu_out_ex_o [16]) );
  AOI21_X1 \dp/ex_stage/alu/U178  ( .B1(\dp/ex_stage/alu/n18 ), .B2(
        \dp/ex_stage/alu/n75 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n185 ) );
  OAI221_X1 \dp/ex_stage/alu/U177  ( .B1(\dp/ex_stage/alu/n185 ), .B2(
        \dp/ex_stage/alu/n57 ), .C1(\dp/ex_stage/alu/n186 ), .C2(
        \dp/ex_stage/alu/n75 ), .A(\dp/ex_stage/alu/n187 ), .ZN(
        \dp/alu_out_ex_o [10]) );
  AOI21_X1 \dp/ex_stage/alu/U176  ( .B1(\dp/ex_stage/alu/n18 ), .B2(
        \dp/ex_stage/alu/n76 ), .A(\dp/ex_stage/alu/n7 ), .ZN(
        \dp/ex_stage/alu/n182 ) );
  OAI221_X1 \dp/ex_stage/alu/U175  ( .B1(\dp/ex_stage/alu/n182 ), .B2(
        \dp/ex_stage/alu/n58 ), .C1(\dp/ex_stage/alu/n183 ), .C2(
        \dp/ex_stage/alu/n76 ), .A(\dp/ex_stage/alu/n184 ), .ZN(
        \dp/alu_out_ex_o [11]) );
  NOR3_X1 \dp/ex_stage/alu/U174  ( .A1(\dp/ex_stage/alu/n223 ), .A2(
        alu_op_i[0]), .A3(\dp/ex_stage/alu/n226 ), .ZN(\dp/ex_stage/alu/n88 )
         );
  NOR4_X1 \dp/ex_stage/alu/U173  ( .A1(\dp/ex_stage/alu/n224 ), .A2(
        \dp/ex_stage/alu/n227 ), .A3(alu_op_i[3]), .A4(alu_op_i[4]), .ZN(
        \dp/ex_stage/alu/n89 ) );
  INV_X1 \dp/ex_stage/alu/U172  ( .A(\dp/ex_stage/muxA_out [1]), .ZN(
        \dp/ex_stage/alu/n33 ) );
  INV_X1 \dp/ex_stage/alu/U171  ( .A(\dp/ex_stage/muxA_out [12]), .ZN(
        \dp/ex_stage/alu/n35 ) );
  INV_X1 \dp/ex_stage/alu/U170  ( .A(\dp/ex_stage/muxA_out [14]), .ZN(
        \dp/ex_stage/alu/n38 ) );
  INV_X1 \dp/ex_stage/alu/U169  ( .A(\dp/ex_stage/muxA_out [15]), .ZN(
        \dp/ex_stage/alu/n39 ) );
  INV_X1 \dp/ex_stage/alu/U168  ( .A(\dp/ex_stage/muxA_out [16]), .ZN(
        \dp/ex_stage/alu/n40 ) );
  INV_X1 \dp/ex_stage/alu/U167  ( .A(\dp/ex_stage/muxB_out [1]), .ZN(
        \dp/ex_stage/alu/n26 ) );
  INV_X1 \dp/ex_stage/alu/U166  ( .A(\dp/ex_stage/muxB_out [4]), .ZN(
        \dp/ex_stage/alu/n32 ) );
  INV_X1 \dp/ex_stage/alu/U165  ( .A(\dp/ex_stage/muxA_out [13]), .ZN(
        \dp/ex_stage/alu/n36 ) );
  INV_X1 \dp/ex_stage/alu/U164  ( .A(\dp/ex_stage/muxB_out [2]), .ZN(
        \dp/ex_stage/alu/n28 ) );
  INV_X1 \dp/ex_stage/alu/U163  ( .A(\dp/ex_stage/alu/n93 ), .ZN(
        \dp/ex_stage/alu/n225 ) );
  NOR3_X1 \dp/ex_stage/alu/U162  ( .A1(\dp/ex_stage/alu/n201 ), .A2(
        alu_op_i[3]), .A3(alu_op_i[0]), .ZN(\dp/ex_stage/alu/n200 ) );
  OAI211_X1 \dp/ex_stage/alu/U161  ( .C1(\dp/ex_stage/alu/n225 ), .C2(
        \dp/ex_stage/alu/n47 ), .A(\dp/ex_stage/alu/n202 ), .B(
        \dp/ex_stage/alu/n203 ), .ZN(\dp/ex_stage/alu/n199 ) );
  AOI21_X1 \dp/ex_stage/alu/U160  ( .B1(alu_op_i[3]), .B2(
        \dp/ex_stage/alu/n199 ), .A(\dp/ex_stage/alu/n200 ), .ZN(
        \dp/ex_stage/alu/n197 ) );
  AOI22_X1 \dp/ex_stage/alu/U159  ( .A1(\dp/ex_stage/alu/N22 ), .A2(
        \dp/ex_stage/alu/n227 ), .B1(\dp/ex_stage/alu/N21 ), .B2(alu_op_i[0]), 
        .ZN(\dp/ex_stage/alu/n196 ) );
  AOI22_X1 \dp/ex_stage/alu/U158  ( .A1(\dp/ex_stage/alu/N17 ), .A2(
        \dp/ex_stage/alu/n226 ), .B1(\dp/ex_stage/alu/N18 ), .B2(alu_op_i[1]), 
        .ZN(\dp/ex_stage/alu/n201 ) );
  AOI222_X1 \dp/ex_stage/alu/U157  ( .A1(\dp/ex_stage/alu/adder_out [0]), .A2(
        \dp/ex_stage/alu/n21 ), .B1(\dp/ex_stage/muxB_out [0]), .B2(
        \dp/ex_stage/alu/n204 ), .C1(\dp/ex_stage/alu/shifter_out [0]), .C2(
        \dp/ex_stage/alu/n24 ), .ZN(\dp/ex_stage/alu/n191 ) );
  NAND2_X1 \dp/ex_stage/alu/U156  ( .A1(\dp/ex_stage/alu/n191 ), .A2(
        \dp/ex_stage/alu/n192 ), .ZN(\dp/alu_out_ex_o [0]) );
  INV_X1 \dp/ex_stage/alu/U155  ( .A(\dp/ex_stage/muxB_out [3]), .ZN(
        \dp/ex_stage/alu/n30 ) );
  OAI21_X1 \dp/ex_stage/alu/U154  ( .B1(\dp/ex_stage/alu/n197 ), .B2(
        \dp/ex_stage/alu/n224 ), .A(\dp/ex_stage/alu/n198 ), .ZN(
        \dp/ex_stage/alu/n194 ) );
  NOR4_X1 \dp/ex_stage/alu/U153  ( .A1(alu_op_i[1]), .A2(
        \dp/ex_stage/alu/n196 ), .A3(\dp/ex_stage/alu/n223 ), .A4(
        \dp/ex_stage/alu/n219 ), .ZN(\dp/ex_stage/alu/n195 ) );
  OAI21_X1 \dp/ex_stage/alu/U152  ( .B1(\dp/ex_stage/muxB_out [0]), .B2(
        \dp/ex_stage/alu/n190 ), .A(\dp/ex_stage/alu/n189 ), .ZN(
        \dp/ex_stage/alu/n193 ) );
  AOI221_X1 \dp/ex_stage/alu/U151  ( .B1(\dp/ex_stage/alu/shifter/N202 ), .B2(
        \dp/ex_stage/alu/n193 ), .C1(\dp/ex_stage/alu/n194 ), .C2(
        \dp/ex_stage/alu/n219 ), .A(\dp/ex_stage/alu/n195 ), .ZN(
        \dp/ex_stage/alu/n192 ) );
  INV_X1 \dp/ex_stage/alu/U150  ( .A(\dp/ex_stage/muxB_out [11]), .ZN(
        \dp/ex_stage/alu/n76 ) );
  INV_X1 \dp/ex_stage/alu/U149  ( .A(\dp/ex_stage/muxB_out [15]), .ZN(
        \dp/ex_stage/alu/n80 ) );
  INV_X1 \dp/ex_stage/alu/U148  ( .A(\dp/ex_stage/muxB_out [19]), .ZN(
        \dp/ex_stage/alu/n84 ) );
  INV_X1 \dp/ex_stage/alu/U147  ( .A(\dp/ex_stage/muxB_out [23]), .ZN(
        \dp/ex_stage/alu/n209 ) );
  INV_X1 \dp/ex_stage/alu/U146  ( .A(\dp/ex_stage/muxB_out [27]), .ZN(
        \dp/ex_stage/alu/n213 ) );
  INV_X1 \dp/ex_stage/alu/U145  ( .A(\dp/ex_stage/muxB_out [13]), .ZN(
        \dp/ex_stage/alu/n78 ) );
  INV_X1 \dp/ex_stage/alu/U144  ( .A(\dp/ex_stage/muxB_out [17]), .ZN(
        \dp/ex_stage/alu/n82 ) );
  INV_X1 \dp/ex_stage/alu/U143  ( .A(\dp/ex_stage/muxB_out [21]), .ZN(
        \dp/ex_stage/alu/n86 ) );
  INV_X1 \dp/ex_stage/alu/U142  ( .A(\dp/ex_stage/muxB_out [25]), .ZN(
        \dp/ex_stage/alu/n211 ) );
  INV_X1 \dp/ex_stage/alu/U141  ( .A(\dp/ex_stage/muxB_out [29]), .ZN(
        \dp/ex_stage/alu/n215 ) );
  INV_X1 \dp/ex_stage/alu/U140  ( .A(\dp/ex_stage/muxB_out [12]), .ZN(
        \dp/ex_stage/alu/n77 ) );
  INV_X1 \dp/ex_stage/alu/U139  ( .A(\dp/ex_stage/muxB_out [16]), .ZN(
        \dp/ex_stage/alu/n81 ) );
  INV_X1 \dp/ex_stage/alu/U138  ( .A(\dp/ex_stage/muxB_out [20]), .ZN(
        \dp/ex_stage/alu/n85 ) );
  INV_X1 \dp/ex_stage/alu/U137  ( .A(\dp/ex_stage/muxB_out [24]), .ZN(
        \dp/ex_stage/alu/n210 ) );
  INV_X1 \dp/ex_stage/alu/U136  ( .A(\dp/ex_stage/muxB_out [28]), .ZN(
        \dp/ex_stage/alu/n214 ) );
  INV_X1 \dp/ex_stage/alu/U135  ( .A(\dp/ex_stage/muxB_out [7]), .ZN(
        \dp/ex_stage/alu/n72 ) );
  INV_X1 \dp/ex_stage/alu/U134  ( .A(\dp/ex_stage/muxB_out [5]), .ZN(
        \dp/ex_stage/alu/n70 ) );
  INV_X1 \dp/ex_stage/alu/U133  ( .A(\dp/ex_stage/muxB_out [9]), .ZN(
        \dp/ex_stage/alu/n74 ) );
  INV_X1 \dp/ex_stage/alu/U132  ( .A(\dp/ex_stage/muxB_out [10]), .ZN(
        \dp/ex_stage/alu/n75 ) );
  INV_X1 \dp/ex_stage/alu/U131  ( .A(\dp/ex_stage/muxB_out [14]), .ZN(
        \dp/ex_stage/alu/n79 ) );
  INV_X1 \dp/ex_stage/alu/U130  ( .A(\dp/ex_stage/muxB_out [18]), .ZN(
        \dp/ex_stage/alu/n83 ) );
  INV_X1 \dp/ex_stage/alu/U129  ( .A(\dp/ex_stage/muxB_out [22]), .ZN(
        \dp/ex_stage/alu/n87 ) );
  INV_X1 \dp/ex_stage/alu/U128  ( .A(\dp/ex_stage/muxB_out [26]), .ZN(
        \dp/ex_stage/alu/n212 ) );
  INV_X1 \dp/ex_stage/alu/U127  ( .A(\dp/ex_stage/muxB_out [8]), .ZN(
        \dp/ex_stage/alu/n73 ) );
  INV_X1 \dp/ex_stage/alu/U126  ( .A(\dp/ex_stage/muxB_out [31]), .ZN(
        \dp/ex_stage/alu/n217 ) );
  INV_X1 \dp/ex_stage/alu/U125  ( .A(\dp/ex_stage/muxB_out [6]), .ZN(
        \dp/ex_stage/alu/n71 ) );
  INV_X1 \dp/ex_stage/alu/U124  ( .A(\dp/ex_stage/muxB_out [30]), .ZN(
        \dp/ex_stage/alu/n216 ) );
  NAND2_X1 \dp/ex_stage/alu/U123  ( .A1(\dp/ex_stage/alu/n205 ), .A2(
        \dp/ex_stage/alu/n92 ), .ZN(\dp/ex_stage/alu/n188 ) );
  INV_X1 \dp/ex_stage/alu/U122  ( .A(\dp/ex_stage/muxA_out [5]), .ZN(
        \dp/ex_stage/alu/n52 ) );
  INV_X1 \dp/ex_stage/alu/U121  ( .A(\dp/ex_stage/alu/shifter/N136 ), .ZN(
        \dp/ex_stage/alu/n69 ) );
  INV_X1 \dp/ex_stage/alu/U120  ( .A(\dp/ex_stage/muxA_out [20]), .ZN(
        \dp/ex_stage/alu/n61 ) );
  INV_X1 \dp/ex_stage/alu/U119  ( .A(\dp/ex_stage/muxA_out [19]), .ZN(
        \dp/ex_stage/alu/n60 ) );
  INV_X1 \dp/ex_stage/alu/U118  ( .A(\dp/ex_stage/muxA_out [30]), .ZN(
        \dp/ex_stage/alu/n68 ) );
  INV_X1 \dp/ex_stage/alu/U117  ( .A(\dp/ex_stage/muxA_out [6]), .ZN(
        \dp/ex_stage/alu/n53 ) );
  INV_X1 \dp/ex_stage/alu/U116  ( .A(\dp/ex_stage/muxA_out [4]), .ZN(
        \dp/ex_stage/alu/n51 ) );
  INV_X1 \dp/ex_stage/alu/U115  ( .A(\dp/ex_stage/muxA_out [29]), .ZN(
        \dp/ex_stage/alu/n67 ) );
  INV_X1 \dp/ex_stage/alu/U114  ( .A(\dp/ex_stage/muxA_out [18]), .ZN(
        \dp/ex_stage/alu/n59 ) );
  NAND2_X1 \dp/ex_stage/alu/U113  ( .A1(\dp/ex_stage/alu/n88 ), .A2(
        \dp/ex_stage/alu/n219 ), .ZN(\dp/ex_stage/alu/n189 ) );
  INV_X1 \dp/ex_stage/alu/U112  ( .A(\dp/ex_stage/muxA_out [24]), .ZN(
        \dp/ex_stage/alu/n62 ) );
  INV_X1 \dp/ex_stage/alu/U111  ( .A(\dp/ex_stage/muxA_out [25]), .ZN(
        \dp/ex_stage/alu/n63 ) );
  INV_X1 \dp/ex_stage/alu/U110  ( .A(\dp/ex_stage/muxA_out [26]), .ZN(
        \dp/ex_stage/alu/n64 ) );
  INV_X1 \dp/ex_stage/alu/U109  ( .A(\dp/ex_stage/muxA_out [27]), .ZN(
        \dp/ex_stage/alu/n65 ) );
  INV_X1 \dp/ex_stage/alu/U108  ( .A(\dp/ex_stage/muxA_out [28]), .ZN(
        \dp/ex_stage/alu/n66 ) );
  INV_X1 \dp/ex_stage/alu/U107  ( .A(\dp/ex_stage/muxA_out [3]), .ZN(
        \dp/ex_stage/alu/n50 ) );
  INV_X1 \dp/ex_stage/alu/U106  ( .A(\dp/ex_stage/muxA_out [9]), .ZN(
        \dp/ex_stage/alu/n56 ) );
  INV_X1 \dp/ex_stage/alu/U105  ( .A(\dp/ex_stage/muxA_out [2]), .ZN(
        \dp/ex_stage/alu/n49 ) );
  INV_X1 \dp/ex_stage/alu/U104  ( .A(\dp/ex_stage/muxA_out [7]), .ZN(
        \dp/ex_stage/alu/n54 ) );
  INV_X1 \dp/ex_stage/alu/U103  ( .A(\dp/ex_stage/muxA_out [8]), .ZN(
        \dp/ex_stage/alu/n55 ) );
  INV_X1 \dp/ex_stage/alu/U102  ( .A(\dp/ex_stage/muxA_out [10]), .ZN(
        \dp/ex_stage/alu/n57 ) );
  INV_X1 \dp/ex_stage/alu/U101  ( .A(\dp/ex_stage/muxA_out [11]), .ZN(
        \dp/ex_stage/alu/n58 ) );
  INV_X1 \dp/ex_stage/alu/U100  ( .A(\dp/ex_stage/alu/n190 ), .ZN(
        \dp/ex_stage/alu/n221 ) );
  BUF_X1 \dp/ex_stage/alu/U99  ( .A(\dp/ex_stage/alu/n97 ), .Z(
        \dp/ex_stage/alu/n21 ) );
  BUF_X1 \dp/ex_stage/alu/U98  ( .A(\dp/ex_stage/alu/n97 ), .Z(
        \dp/ex_stage/alu/n20 ) );
  BUF_X1 \dp/ex_stage/alu/U97  ( .A(\dp/ex_stage/alu/n97 ), .Z(
        \dp/ex_stage/alu/n19 ) );
  BUF_X1 \dp/ex_stage/alu/U96  ( .A(\dp/ex_stage/alu/n89 ), .Z(
        \dp/ex_stage/alu/n23 ) );
  BUF_X1 \dp/ex_stage/alu/U95  ( .A(\dp/ex_stage/alu/n89 ), .Z(
        \dp/ex_stage/alu/n22 ) );
  INV_X1 \dp/ex_stage/alu/U94  ( .A(\dp/ex_stage/alu/shifter/N202 ), .ZN(
        \dp/ex_stage/alu/n48 ) );
  OAI221_X1 \dp/ex_stage/alu/U93  ( .B1(\dp/ex_stage/alu/shifter/N202 ), .B2(
        \dp/ex_stage/alu/n190 ), .C1(\dp/ex_stage/alu/n188 ), .C2(
        \dp/ex_stage/alu/n48 ), .A(\dp/ex_stage/alu/n189 ), .ZN(
        \dp/ex_stage/alu/n204 ) );
  AOI221_X1 \dp/ex_stage/alu/U92  ( .B1(\dp/ex_stage/muxA_out [2]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n49 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n123 ) );
  AOI221_X1 \dp/ex_stage/alu/U91  ( .B1(\dp/ex_stage/muxA_out [3]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n50 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n114 ) );
  AOI221_X1 \dp/ex_stage/alu/U90  ( .B1(\dp/ex_stage/muxA_out [4]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n51 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n111 ) );
  AOI221_X1 \dp/ex_stage/alu/U89  ( .B1(\dp/ex_stage/muxA_out [5]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n52 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n108 ) );
  AOI221_X1 \dp/ex_stage/alu/U88  ( .B1(\dp/ex_stage/muxA_out [6]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n53 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n105 ) );
  AOI221_X1 \dp/ex_stage/alu/U87  ( .B1(\dp/ex_stage/muxA_out [7]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n54 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n102 ) );
  AOI221_X1 \dp/ex_stage/alu/U86  ( .B1(\dp/ex_stage/muxA_out [8]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n55 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n99 ) );
  AOI221_X1 \dp/ex_stage/alu/U85  ( .B1(\dp/ex_stage/muxA_out [28]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n66 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n129 ) );
  AOI221_X1 \dp/ex_stage/alu/U84  ( .B1(\dp/ex_stage/muxA_out [29]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n67 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n126 ) );
  AOI221_X1 \dp/ex_stage/alu/U83  ( .B1(\dp/ex_stage/muxA_out [30]), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n68 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n120 ) );
  AOI221_X1 \dp/ex_stage/alu/U82  ( .B1(\dp/ex_stage/alu/shifter/N136 ), .B2(
        \dp/ex_stage/alu/n8 ), .C1(\dp/ex_stage/alu/n11 ), .C2(
        \dp/ex_stage/alu/n69 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n117 ) );
  AOI221_X1 \dp/ex_stage/alu/U81  ( .B1(\dp/ex_stage/muxA_out [10]), .B2(
        \dp/ex_stage/alu/n10 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n57 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n186 ) );
  AOI221_X1 \dp/ex_stage/alu/U80  ( .B1(\dp/ex_stage/muxA_out [11]), .B2(
        \dp/ex_stage/alu/n10 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n58 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n183 ) );
  AOI221_X1 \dp/ex_stage/alu/U79  ( .B1(\dp/ex_stage/alu/n34 ), .B2(
        \dp/ex_stage/alu/n10 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n35 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n180 ) );
  AOI221_X1 \dp/ex_stage/alu/U78  ( .B1(\dp/ex_stage/muxA_out [13]), .B2(
        \dp/ex_stage/alu/n10 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n36 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n177 ) );
  AOI221_X1 \dp/ex_stage/alu/U77  ( .B1(\dp/ex_stage/alu/n37 ), .B2(
        \dp/ex_stage/alu/n10 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n38 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n174 ) );
  AOI221_X1 \dp/ex_stage/alu/U76  ( .B1(\dp/ex_stage/muxA_out [15]), .B2(
        \dp/ex_stage/alu/n10 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n39 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n171 ) );
  AOI221_X1 \dp/ex_stage/alu/U75  ( .B1(\dp/ex_stage/muxA_out [16]), .B2(
        \dp/ex_stage/alu/n10 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n40 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n168 ) );
  AOI221_X1 \dp/ex_stage/alu/U74  ( .B1(\dp/ex_stage/muxA_out [1]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n33 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n156 ) );
  AOI221_X1 \dp/ex_stage/alu/U73  ( .B1(\dp/ex_stage/alu/n8 ), .B2(
        \dp/ex_stage/muxA_out [9]), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n56 ), .A(\dp/ex_stage/alu/n3 ), .ZN(
        \dp/ex_stage/alu/n95 ) );
  AOI221_X1 \dp/ex_stage/alu/U72  ( .B1(\dp/ex_stage/muxA_out [17]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n41 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n165 ) );
  AOI221_X1 \dp/ex_stage/alu/U71  ( .B1(\dp/ex_stage/muxA_out [18]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n59 ), .A(\dp/ex_stage/alu/n5 ), .ZN(
        \dp/ex_stage/alu/n162 ) );
  AOI221_X1 \dp/ex_stage/alu/U70  ( .B1(\dp/ex_stage/muxA_out [19]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n15 ), .C2(
        \dp/ex_stage/alu/n60 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n159 ) );
  AOI221_X1 \dp/ex_stage/alu/U69  ( .B1(\dp/ex_stage/muxA_out [20]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n61 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n153 ) );
  AOI221_X1 \dp/ex_stage/alu/U68  ( .B1(\dp/ex_stage/muxA_out [21]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n42 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n150 ) );
  AOI221_X1 \dp/ex_stage/alu/U67  ( .B1(\dp/ex_stage/alu/n43 ), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n44 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n147 ) );
  AOI221_X1 \dp/ex_stage/alu/U66  ( .B1(\dp/ex_stage/alu/n45 ), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n46 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n144 ) );
  AOI221_X1 \dp/ex_stage/alu/U65  ( .B1(\dp/ex_stage/muxA_out [24]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n62 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n141 ) );
  AOI221_X1 \dp/ex_stage/alu/U64  ( .B1(\dp/ex_stage/muxA_out [25]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n63 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n138 ) );
  AOI221_X1 \dp/ex_stage/alu/U63  ( .B1(\dp/ex_stage/muxA_out [26]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n64 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n135 ) );
  AOI221_X1 \dp/ex_stage/alu/U62  ( .B1(\dp/ex_stage/muxA_out [27]), .B2(
        \dp/ex_stage/alu/n9 ), .C1(\dp/ex_stage/alu/n14 ), .C2(
        \dp/ex_stage/alu/n65 ), .A(\dp/ex_stage/alu/n4 ), .ZN(
        \dp/ex_stage/alu/n132 ) );
  INV_X1 \dp/ex_stage/alu/U61  ( .A(\dp/ex_stage/alu/n92 ), .ZN(
        \dp/ex_stage/alu/n223 ) );
  AND2_X1 \dp/ex_stage/alu/U60  ( .A1(\dp/ex_stage/alu/n226 ), .A2(
        \dp/ex_stage/alu/n24 ), .ZN(\dp/ex_stage/alu/n208 ) );
  NAND4_X1 \dp/ex_stage/alu/U59  ( .A1(\dp/ex_stage/alu/n227 ), .A2(
        \dp/ex_stage/alu/n226 ), .A3(\dp/ex_stage/alu/n224 ), .A4(
        \dp/ex_stage/alu/n219 ), .ZN(\dp/ex_stage/alu/n90 ) );
  AOI22_X1 \dp/ex_stage/alu/U58  ( .A1(\dp/ex_stage/alu/shifter_out [4]), .A2(
        \dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [4]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n112 ) );
  AOI22_X1 \dp/ex_stage/alu/U57  ( .A1(\dp/ex_stage/alu/shifter_out [8]), .A2(
        \dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [8]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n100 ) );
  AOI22_X1 \dp/ex_stage/alu/U56  ( .A1(\dp/ex_stage/alu/shifter_out [12]), 
        .A2(\dp/ex_stage/alu/n24 ), .B1(\dp/ex_stage/alu/adder_out [12]), .B2(
        \dp/ex_stage/alu/n21 ), .ZN(\dp/ex_stage/alu/n181 ) );
  BUF_X1 \dp/ex_stage/alu/U55  ( .A(\dp/ex_stage/alu/n89 ), .Z(
        \dp/ex_stage/alu/n24 ) );
  NOR2_X1 \dp/ex_stage/alu/U54  ( .A1(\dp/ex_stage/alu/n227 ), .A2(
        \dp/ex_stage/alu/n226 ), .ZN(\dp/ex_stage/alu/n93 ) );
  INV_X1 \dp/ex_stage/alu/U53  ( .A(\dp/ex_stage/alu/n44 ), .ZN(
        \dp/ex_stage/alu/n43 ) );
  NAND2_X1 \dp/ex_stage/alu/U52  ( .A1(\dp/ex_stage/alu/N19 ), .A2(
        \dp/ex_stage/alu/n226 ), .ZN(\dp/ex_stage/alu/n203 ) );
  INV_X1 \dp/ex_stage/alu/U51  ( .A(\dp/ex_stage/alu/n28 ), .ZN(
        \dp/ex_stage/alu/n27 ) );
  INV_X1 \dp/ex_stage/alu/U50  ( .A(\dp/ex_stage/alu/n189 ), .ZN(
        \dp/ex_stage/alu/n218 ) );
  INV_X1 \dp/ex_stage/alu/U49  ( .A(\dp/ex_stage/alu/n188 ), .ZN(
        \dp/ex_stage/alu/n220 ) );
  BUF_X1 \dp/ex_stage/alu/U48  ( .A(\dp/ex_stage/alu/n221 ), .Z(
        \dp/ex_stage/alu/n15 ) );
  BUF_X1 \dp/ex_stage/alu/U47  ( .A(\dp/ex_stage/alu/n221 ), .Z(
        \dp/ex_stage/alu/n14 ) );
  BUF_X1 \dp/ex_stage/alu/U46  ( .A(\dp/ex_stage/alu/n221 ), .Z(
        \dp/ex_stage/alu/n11 ) );
  BUF_X1 \dp/ex_stage/alu/U45  ( .A(\dp/ex_stage/alu/n221 ), .Z(
        \dp/ex_stage/alu/n17 ) );
  BUF_X1 \dp/ex_stage/alu/U44  ( .A(\dp/ex_stage/alu/n221 ), .Z(
        \dp/ex_stage/alu/n16 ) );
  AOI22_X1 \dp/ex_stage/alu/U43  ( .A1(\dp/ex_stage/alu/shifter_out [15]), 
        .A2(\dp/ex_stage/alu/n24 ), .B1(\dp/ex_stage/alu/adder_out [15]), .B2(
        \dp/ex_stage/alu/n21 ), .ZN(\dp/ex_stage/alu/n172 ) );
  AOI22_X1 \dp/ex_stage/alu/U42  ( .A1(\dp/ex_stage/alu/shifter_out [23]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [23]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n145 ) );
  AOI22_X1 \dp/ex_stage/alu/U41  ( .A1(\dp/ex_stage/alu/shifter_out [27]), 
        .A2(\dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [27]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n133 ) );
  AOI22_X1 \dp/ex_stage/alu/U40  ( .A1(\dp/ex_stage/alu/shifter_out [31]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [31]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n118 ) );
  AOI22_X1 \dp/ex_stage/alu/U39  ( .A1(\dp/ex_stage/alu/shifter_out [19]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [19]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n160 ) );
  AOI22_X1 \dp/ex_stage/alu/U38  ( .A1(\dp/ex_stage/alu/shifter_out [1]), .A2(
        \dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [1]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n157 ) );
  AOI22_X1 \dp/ex_stage/alu/U37  ( .A1(\dp/ex_stage/alu/shifter_out [2]), .A2(
        \dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [2]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n124 ) );
  AOI22_X1 \dp/ex_stage/alu/U36  ( .A1(\dp/ex_stage/alu/shifter_out [3]), .A2(
        \dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [3]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n115 ) );
  AOI22_X1 \dp/ex_stage/alu/U35  ( .A1(\dp/ex_stage/alu/shifter_out [5]), .A2(
        \dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [5]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n109 ) );
  AOI22_X1 \dp/ex_stage/alu/U34  ( .A1(\dp/ex_stage/alu/shifter_out [6]), .A2(
        \dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [6]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n106 ) );
  AOI22_X1 \dp/ex_stage/alu/U33  ( .A1(\dp/ex_stage/alu/shifter_out [7]), .A2(
        \dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [7]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n103 ) );
  AOI22_X1 \dp/ex_stage/alu/U32  ( .A1(\dp/ex_stage/alu/shifter_out [9]), .A2(
        \dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [9]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n96 ) );
  AOI22_X1 \dp/ex_stage/alu/U31  ( .A1(\dp/ex_stage/alu/shifter_out [17]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [17]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n166 ) );
  AOI22_X1 \dp/ex_stage/alu/U30  ( .A1(\dp/ex_stage/alu/shifter_out [18]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [18]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n163 ) );
  AOI22_X1 \dp/ex_stage/alu/U29  ( .A1(\dp/ex_stage/alu/shifter_out [20]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [20]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n154 ) );
  AOI22_X1 \dp/ex_stage/alu/U28  ( .A1(\dp/ex_stage/alu/shifter_out [21]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [21]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n151 ) );
  AOI22_X1 \dp/ex_stage/alu/U27  ( .A1(\dp/ex_stage/alu/shifter_out [22]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [22]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n148 ) );
  AOI22_X1 \dp/ex_stage/alu/U26  ( .A1(\dp/ex_stage/alu/shifter_out [24]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [24]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n142 ) );
  AOI22_X1 \dp/ex_stage/alu/U25  ( .A1(\dp/ex_stage/alu/shifter_out [25]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [25]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n139 ) );
  AOI22_X1 \dp/ex_stage/alu/U24  ( .A1(\dp/ex_stage/alu/shifter_out [26]), 
        .A2(\dp/ex_stage/alu/n23 ), .B1(\dp/ex_stage/alu/adder_out [26]), .B2(
        \dp/ex_stage/alu/n20 ), .ZN(\dp/ex_stage/alu/n136 ) );
  AOI22_X1 \dp/ex_stage/alu/U23  ( .A1(\dp/ex_stage/alu/shifter_out [28]), 
        .A2(\dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [28]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n130 ) );
  AOI22_X1 \dp/ex_stage/alu/U22  ( .A1(\dp/ex_stage/alu/shifter_out [29]), 
        .A2(\dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [29]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n127 ) );
  AOI22_X1 \dp/ex_stage/alu/U21  ( .A1(\dp/ex_stage/alu/shifter_out [30]), 
        .A2(\dp/ex_stage/alu/n22 ), .B1(\dp/ex_stage/alu/adder_out [30]), .B2(
        \dp/ex_stage/alu/n19 ), .ZN(\dp/ex_stage/alu/n121 ) );
  AOI22_X1 \dp/ex_stage/alu/U20  ( .A1(\dp/ex_stage/alu/shifter_out [10]), 
        .A2(\dp/ex_stage/alu/n24 ), .B1(\dp/ex_stage/alu/adder_out [10]), .B2(
        \dp/ex_stage/alu/n21 ), .ZN(\dp/ex_stage/alu/n187 ) );
  AOI22_X1 \dp/ex_stage/alu/U19  ( .A1(\dp/ex_stage/alu/shifter_out [11]), 
        .A2(\dp/ex_stage/alu/n24 ), .B1(\dp/ex_stage/alu/adder_out [11]), .B2(
        \dp/ex_stage/alu/n21 ), .ZN(\dp/ex_stage/alu/n184 ) );
  AOI22_X1 \dp/ex_stage/alu/U18  ( .A1(\dp/ex_stage/alu/shifter_out [13]), 
        .A2(\dp/ex_stage/alu/n24 ), .B1(\dp/ex_stage/alu/adder_out [13]), .B2(
        \dp/ex_stage/alu/n21 ), .ZN(\dp/ex_stage/alu/n178 ) );
  AOI22_X1 \dp/ex_stage/alu/U17  ( .A1(\dp/ex_stage/alu/shifter_out [14]), 
        .A2(\dp/ex_stage/alu/n24 ), .B1(\dp/ex_stage/alu/adder_out [14]), .B2(
        \dp/ex_stage/alu/n21 ), .ZN(\dp/ex_stage/alu/n175 ) );
  AOI22_X1 \dp/ex_stage/alu/U16  ( .A1(\dp/ex_stage/alu/shifter_out [16]), 
        .A2(\dp/ex_stage/alu/n24 ), .B1(\dp/ex_stage/alu/adder_out [16]), .B2(
        \dp/ex_stage/alu/n21 ), .ZN(\dp/ex_stage/alu/n169 ) );
  INV_X1 \dp/ex_stage/alu/U15  ( .A(\dp/ex_stage/alu/N21 ), .ZN(
        \dp/ex_stage/alu/n47 ) );
  BUF_X1 \dp/ex_stage/alu/U14  ( .A(\dp/ex_stage/alu/n218 ), .Z(
        \dp/ex_stage/alu/n2 ) );
  BUF_X1 \dp/ex_stage/alu/U13  ( .A(\dp/ex_stage/alu/n218 ), .Z(
        \dp/ex_stage/alu/n1 ) );
  BUF_X1 \dp/ex_stage/alu/U12  ( .A(\dp/ex_stage/alu/n220 ), .Z(
        \dp/ex_stage/alu/n10 ) );
  BUF_X1 \dp/ex_stage/alu/U11  ( .A(\dp/ex_stage/alu/n220 ), .Z(
        \dp/ex_stage/alu/n8 ) );
  BUF_X1 \dp/ex_stage/alu/U10  ( .A(\dp/ex_stage/alu/n220 ), .Z(
        \dp/ex_stage/alu/n9 ) );
  BUF_X1 \dp/ex_stage/alu/U9  ( .A(\dp/ex_stage/alu/n1 ), .Z(
        \dp/ex_stage/alu/n5 ) );
  BUF_X1 \dp/ex_stage/alu/U8  ( .A(\dp/ex_stage/alu/n2 ), .Z(
        \dp/ex_stage/alu/n6 ) );
  BUF_X1 \dp/ex_stage/alu/U7  ( .A(\dp/ex_stage/alu/n2 ), .Z(
        \dp/ex_stage/alu/n7 ) );
  BUF_X1 \dp/ex_stage/alu/U5  ( .A(\dp/ex_stage/alu/n1 ), .Z(
        \dp/ex_stage/alu/n4 ) );
  BUF_X1 \dp/ex_stage/alu/U4  ( .A(\dp/ex_stage/alu/n1 ), .Z(
        \dp/ex_stage/alu/n3 ) );
  NAND3_X1 \dp/ex_stage/alu/U235  ( .A1(alu_op_i[1]), .A2(
        \dp/ex_stage/alu/n224 ), .A3(alu_op_i[3]), .ZN(\dp/ex_stage/alu/n206 )
         );
  NAND3_X1 \dp/ex_stage/alu/U234  ( .A1(\dp/ex_stage/alu/n206 ), .A2(
        \dp/ex_stage/alu/n90 ), .A3(\dp/ex_stage/alu/n207 ), .ZN(
        \dp/ex_stage/alu/n97 ) );
  NAND3_X1 \dp/ex_stage/alu/U233  ( .A1(alu_op_i[3]), .A2(
        \dp/ex_stage/alu/n224 ), .A3(\dp/ex_stage/alu/n205 ), .ZN(
        \dp/ex_stage/alu/n190 ) );
  NAND3_X1 \dp/ex_stage/alu/U232  ( .A1(alu_op_i[1]), .A2(
        \dp/ex_stage/alu/n227 ), .A3(\dp/ex_stage/alu/N20 ), .ZN(
        \dp/ex_stage/alu/n202 ) );
  NAND3_X1 \dp/ex_stage/alu/U231  ( .A1(\dp/ex_stage/alu/n93 ), .A2(
        \dp/ex_stage/alu/n92 ), .A3(\dp/ex_stage/alu/N16 ), .ZN(
        \dp/ex_stage/alu/n198 ) );
  NAND3_X1 \dp/ex_stage/alu/U230  ( .A1(alu_op_i[4]), .A2(
        \dp/ex_stage/alu/n92 ), .A3(\dp/ex_stage/alu/n93 ), .ZN(
        \dp/ex_stage/alu/n91 ) );
  BUF_X1 \dp/ex_stage/alu/adder/U36  ( .A(\dp/ex_stage/alu/N23 ), .Z(
        \dp/ex_stage/alu/adder/n3 ) );
  BUF_X1 \dp/ex_stage/alu/adder/U35  ( .A(\dp/ex_stage/alu/N23 ), .Z(
        \dp/ex_stage/alu/adder/n2 ) );
  BUF_X1 \dp/ex_stage/alu/adder/U34  ( .A(\dp/ex_stage/alu/N23 ), .Z(
        \dp/ex_stage/alu/adder/n1 ) );
  OR2_X1 \dp/ex_stage/alu/adder/U1  ( .A1(\dp/ex_stage/alu/N23 ), .A2(
        \dp/ex_stage/alu/adder/n3 ), .ZN(\dp/ex_stage/alu/adder/carries [0])
         );
  XOR2_X1 \dp/ex_stage/alu/adder/U33  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [0]), .Z(\dp/ex_stage/alu/adder/B_xor[0] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U32  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [10]), .Z(\dp/ex_stage/alu/adder/B_xor[10] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U31  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [11]), .Z(\dp/ex_stage/alu/adder/B_xor[11] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U30  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [12]), .Z(\dp/ex_stage/alu/adder/B_xor[12] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U29  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [13]), .Z(\dp/ex_stage/alu/adder/B_xor[13] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U28  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [14]), .Z(\dp/ex_stage/alu/adder/B_xor[14] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U27  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [15]), .Z(\dp/ex_stage/alu/adder/B_xor[15] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U26  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [16]), .Z(\dp/ex_stage/alu/adder/B_xor[16] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U25  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [17]), .Z(\dp/ex_stage/alu/adder/B_xor[17] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U24  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [18]), .Z(\dp/ex_stage/alu/adder/B_xor[18] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U23  ( .A(\dp/ex_stage/alu/adder/n1 ), .B(
        \dp/ex_stage/muxB_out [19]), .Z(\dp/ex_stage/alu/adder/B_xor[19] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U22  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/alu/n25 ), .Z(\dp/ex_stage/alu/adder/B_xor[1] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U21  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [20]), .Z(\dp/ex_stage/alu/adder/B_xor[20] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U20  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [21]), .Z(\dp/ex_stage/alu/adder/B_xor[21] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U19  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [22]), .Z(\dp/ex_stage/alu/adder/B_xor[22] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U18  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [23]), .Z(\dp/ex_stage/alu/adder/B_xor[23] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U17  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [24]), .Z(\dp/ex_stage/alu/adder/B_xor[24] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U16  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [25]), .Z(\dp/ex_stage/alu/adder/B_xor[25] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U15  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [26]), .Z(\dp/ex_stage/alu/adder/B_xor[26] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U14  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [27]), .Z(\dp/ex_stage/alu/adder/B_xor[27] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U13  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [28]), .Z(\dp/ex_stage/alu/adder/B_xor[28] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U12  ( .A(\dp/ex_stage/alu/adder/n2 ), .B(
        \dp/ex_stage/muxB_out [29]), .Z(\dp/ex_stage/alu/adder/B_xor[29] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U11  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/alu/n27 ), .Z(\dp/ex_stage/alu/adder/B_xor[2] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U10  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/muxB_out [30]), .Z(\dp/ex_stage/alu/adder/B_xor[30] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U9  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/muxB_out [31]), .Z(\dp/ex_stage/alu/adder/B_xor[31] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U8  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/alu/n29 ), .Z(\dp/ex_stage/alu/adder/B_xor[3] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U7  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/alu/n31 ), .Z(\dp/ex_stage/alu/adder/B_xor[4] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U6  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/muxB_out [5]), .Z(\dp/ex_stage/alu/adder/B_xor[5] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U5  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/muxB_out [6]), .Z(\dp/ex_stage/alu/adder/B_xor[6] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U4  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/muxB_out [7]), .Z(\dp/ex_stage/alu/adder/B_xor[7] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U3  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/muxB_out [8]), .Z(\dp/ex_stage/alu/adder/B_xor[8] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/U2  ( .A(\dp/ex_stage/alu/adder/n3 ), .B(
        \dp/ex_stage/muxB_out [9]), .Z(\dp/ex_stage/alu/adder/B_xor[9] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_1/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[0] ), .A2(\dp/ex_stage/alu/shifter/N202 ), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[1][1] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_1/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[0] ), .B(\dp/ex_stage/alu/shifter/N202 ), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[1][1] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_2/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[1] ), .A2(\dp/ex_stage/muxA_out [1]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[2][2] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_2/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[1] ), .B(\dp/ex_stage/muxA_out [1]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[2][2] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_3/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[2] ), .A2(\dp/ex_stage/muxA_out [2]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[3][3] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_3/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[2] ), .B(\dp/ex_stage/muxA_out [2]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[3][3] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_4/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[3] ), .A2(\dp/ex_stage/muxA_out [3]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[4][4] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_4/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[3] ), .B(\dp/ex_stage/muxA_out [3]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[4][4] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_5/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[4] ), .A2(\dp/ex_stage/muxA_out [4]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[5][5] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_5/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[4] ), .B(\dp/ex_stage/muxA_out [4]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[5][5] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_6/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[5] ), .A2(\dp/ex_stage/muxA_out [5]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[6][6] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_6/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[5] ), .B(\dp/ex_stage/muxA_out [5]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[6][6] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_7/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[6] ), .A2(\dp/ex_stage/muxA_out [6]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[7][7] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_7/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[6] ), .B(\dp/ex_stage/muxA_out [6]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[7][7] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_8/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[7] ), .A2(\dp/ex_stage/muxA_out [7]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[8][8] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_8/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[7] ), .B(\dp/ex_stage/muxA_out [7]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[8][8] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_9/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[8] ), .A2(\dp/ex_stage/muxA_out [8]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[9][9] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_9/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[8] ), .B(\dp/ex_stage/muxA_out [8]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[9][9] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_10/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[9] ), .A2(\dp/ex_stage/muxA_out [9]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[10][10] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_10/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[9] ), .B(\dp/ex_stage/muxA_out [9]), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[10][10] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_11/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[10] ), .A2(\dp/ex_stage/muxA_out [10]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[11][11] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_11/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[10] ), .B(\dp/ex_stage/muxA_out [10]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[11][11] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_12/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[11] ), .A2(\dp/ex_stage/muxA_out [11]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[12][12] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_12/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[11] ), .B(\dp/ex_stage/muxA_out [11]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[12][12] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_13/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[12] ), .A2(\dp/ex_stage/alu/n34 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[13][13] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_13/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[12] ), .B(\dp/ex_stage/alu/n34 ), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[13][13] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_14/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[13] ), .A2(\dp/ex_stage/muxA_out [13]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[14][14] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_14/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[13] ), .B(\dp/ex_stage/muxA_out [13]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[14][14] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_15/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[14] ), .A2(\dp/ex_stage/alu/n37 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[15][15] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_15/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[14] ), .B(\dp/ex_stage/alu/n37 ), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[15][15] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_16/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[15] ), .A2(\dp/ex_stage/muxA_out [15]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[16][16] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_16/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[15] ), .B(\dp/ex_stage/muxA_out [15]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[16][16] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_17/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[16] ), .A2(\dp/ex_stage/muxA_out [16]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[17][17] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_17/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[16] ), .B(\dp/ex_stage/muxA_out [16]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[17][17] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_18/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[17] ), .A2(\dp/ex_stage/muxA_out [17]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[18][18] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_18/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[17] ), .B(\dp/ex_stage/muxA_out [17]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[18][18] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_19/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[18] ), .A2(\dp/ex_stage/muxA_out [18]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[19][19] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_19/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[18] ), .B(\dp/ex_stage/muxA_out [18]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[19][19] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_20/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[19] ), .A2(\dp/ex_stage/muxA_out [19]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[20][20] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_20/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[19] ), .B(\dp/ex_stage/muxA_out [19]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[20][20] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_21/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[20] ), .A2(\dp/ex_stage/muxA_out [20]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[21][21] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_21/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[20] ), .B(\dp/ex_stage/muxA_out [20]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[21][21] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_22/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[21] ), .A2(\dp/ex_stage/muxA_out [21]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[22][22] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_22/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[21] ), .B(\dp/ex_stage/muxA_out [21]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[22][22] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_23/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[22] ), .A2(\dp/ex_stage/alu/n43 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[23][23] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_23/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[22] ), .B(\dp/ex_stage/alu/n43 ), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[23][23] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_24/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[23] ), .A2(\dp/ex_stage/alu/n45 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][24] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_24/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[23] ), .B(\dp/ex_stage/alu/n45 ), .Z(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][24] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_25/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[24] ), .A2(\dp/ex_stage/muxA_out [24]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[25][25] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_25/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[24] ), .B(\dp/ex_stage/muxA_out [24]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[25][25] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_26/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[25] ), .A2(\dp/ex_stage/muxA_out [25]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[26][26] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_26/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[25] ), .B(\dp/ex_stage/muxA_out [25]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[26][26] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_27/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[26] ), .A2(\dp/ex_stage/muxA_out [26]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[27][27] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_27/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[26] ), .B(\dp/ex_stage/muxA_out [26]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[27][27] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_28/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[27] ), .A2(\dp/ex_stage/muxA_out [27]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[28][28] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_28/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[27] ), .B(\dp/ex_stage/muxA_out [27]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[28][28] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_29/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[28] ), .A2(\dp/ex_stage/muxA_out [28]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[29][29] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_29/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[28] ), .B(\dp/ex_stage/muxA_out [28]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[29][29] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_30/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[29] ), .A2(\dp/ex_stage/muxA_out [29]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[30][30] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_30/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[29] ), .B(\dp/ex_stage/muxA_out [29]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[30][30] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_31/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[30] ), .A2(\dp/ex_stage/muxA_out [30]), 
        .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[31][31] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_31/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[30] ), .B(\dp/ex_stage/muxA_out [30]), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[31][31] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_32/U1  ( .A1(
        \dp/ex_stage/alu/adder/B_xor[31] ), .A2(\dp/ex_stage/alu/shifter/N136 ), .ZN(\dp/ex_stage/alu/adder/SparseTree/gen[32][32] ) );
  XOR2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_net_i_32/U2  ( .A(
        \dp/ex_stage/alu/adder/B_xor[31] ), .B(\dp/ex_stage/alu/shifter/N136 ), 
        .Z(\dp/ex_stage/alu/adder/SparseTree/prop[32][32] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G10/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[1][1] ), .B2(
        \dp/ex_stage/alu/adder/carries [0]), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[1][1] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G10/n2 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G10/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G10/n2 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[1][0] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G20_1/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[2][2] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/gen[1][0] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[2][2] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G20_1/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G20_1/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G20_1/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[2][0] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_0/U3  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[3][3] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[4][4] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[4][4] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_0/n2 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_0/U2  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_0/n2 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[4][3] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_0/U1  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[3][3] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[4][4] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[4][3] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_1/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[5][5] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[6][6] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[6][5] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_1/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[5][5] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[6][6] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[6][6] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_1/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_1/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_1/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[6][5] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_2/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[7][7] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[8][8] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[8][7] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_2/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[7][7] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[8][8] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[8][8] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_2/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_2/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_2/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[8][7] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_3/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[9][9] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[10][10] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[10][9] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_3/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[9][9] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[10][10] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[10][10] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_3/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_3/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_3/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[10][9] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_4/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[11][11] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[12][12] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[12][11] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_4/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[11][11] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[12][12] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[12][12] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_4/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_4/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_4/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[12][11] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_5/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[13][13] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[14][14] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[14][13] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_5/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[13][13] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[14][14] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[14][14] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_5/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_5/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_5/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[14][13] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_6/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[15][15] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][16] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][15] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_6/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[15][15] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][16] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[16][16] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_6/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_6/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_6/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[16][15] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_7/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[17][17] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[18][18] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[18][17] ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_7/U2  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_7/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[18][17] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_7/U1  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[17][17] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[18][18] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[18][18] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_7/n3 ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_8/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[19][19] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[20][20] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[20][19] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_8/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[19][19] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[20][20] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[20][20] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_8/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_8/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_8/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[20][19] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_9/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[21][21] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[22][22] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[22][21] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_9/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[21][21] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[22][22] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[22][22] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_9/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_9/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_9/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[22][21] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_10/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[23][23] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][24] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][23] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_10/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[23][23] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][24] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][24] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_10/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_10/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_10/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][23] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_11/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[25][25] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[26][26] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[26][25] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_11/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[25][25] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[26][26] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[26][26] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_11/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_11/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_11/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[26][25] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_12/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[27][27] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][28] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][27] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_12/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[27][27] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][28] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[28][28] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_12/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_12/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_12/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[28][27] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_13/U3  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[29][29] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[30][30] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[30][30] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_13/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_13/U2  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_13/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[30][29] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_13/U1  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[29][29] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[30][30] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[30][29] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_14/U3  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[31][31] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][32] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][32] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_14/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_14/U2  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_14/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][31] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_1_14/U1  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[31][31] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][32] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][31] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_2/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[4][3] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/gen[2][0] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[4][3] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_2/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_2/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_2/n3 ), .ZN(
        \dp/ex_stage/alu/adder/carries [1]) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_0/U3  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[6][5] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[8][7] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[8][7] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_0/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_0/U2  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_0/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[8][5] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_0/U1  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[6][5] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[8][7] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[8][5] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_1/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[10][9] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[12][11] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[12][9] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_1/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[10][9] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[12][11] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[12][11] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_1/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_1/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_1/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[12][9] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_2/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[14][13] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][15] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][13] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_2/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[14][13] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][15] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[16][15] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_2/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_2/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_2/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[16][13] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_3/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[18][17] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[20][19] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[20][17] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_3/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[18][17] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[20][19] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[20][19] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_3/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_3/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_3/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[20][17] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_4/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[22][21] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][23] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][21] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_4/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[22][21] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][23] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][23] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_4/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_4/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_4/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][21] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_5/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[26][25] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][27] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][25] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_5/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[26][25] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][27] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[28][27] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_5/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_5/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_5/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[28][25] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_6/U3  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[30][29] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][31] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][29] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_6/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[30][29] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][31] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][31] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_6/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_6/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_2_6/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][29] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_3/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[8][5] ), .B2(
        \dp/ex_stage/alu/adder/carries [1]), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[8][5] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_3/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_3/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_3/n3 ), .ZN(
        \dp/ex_stage/alu/adder/carries [2]) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_0/U3  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_0/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[16][9] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_0/U2  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[12][9] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][13] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][9] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_0/U1  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[12][9] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][13] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[16][13] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_0/n3 ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_1/U3  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[20][17] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][21] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][21] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_1/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_1/U2  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_1/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][17] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_1/U1  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[20][17] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][21] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][17] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_2/U3  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[28][25] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][29] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][29] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_2/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_2/U2  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_2/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][25] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_3_2/U1  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][25] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][29] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][25] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_4/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[16][9] ), .B2(
        \dp/ex_stage/alu/adder/carries [2]), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[16][9] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_4/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_4/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_4/n3 ), .ZN(
        \dp/ex_stage/alu/adder/carries [4]) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G_2n_0_4_1/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[12][9] ), .B2(
        \dp/ex_stage/alu/adder/carries [2]), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[12][9] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G_2n_0_4_1/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G_2n_0_4_1/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G_2n_0_4_1/n3 ), .ZN(
        \dp/ex_stage/alu/adder/carries [3]) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_0_0/U3  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][17] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][25] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][25] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_0_0/n3 ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_0_0/U2  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][17] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][25] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][17] ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_0_0/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_0_0/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][17] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_1_0/U3  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][17] ), .B2(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][25] ), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[28][25] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_1_0/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_1_0/U2  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_1_0/n3 ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/gen[28][17] ) );
  AND2_X1 \dp/ex_stage/alu/adder/SparseTree/PG_ij_4_1_0/U1  ( .A1(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][17] ), .A2(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][25] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][17] ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_5/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[32][17] ), .B2(
        \dp/ex_stage/alu/adder/carries [4]), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[32][17] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_5/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_5/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G_2exp_0_5/n3 ), .ZN(
        \dp/ex_stage/alu/adder/Cout ) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_1/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[28][17] ), .B2(
        \dp/ex_stage/alu/adder/carries [4]), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[28][17] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_1/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_1/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_1/n3 ), .ZN(
        \dp/ex_stage/alu/adder/carries [7]) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_2/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[24][17] ), .B2(
        \dp/ex_stage/alu/adder/carries [4]), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[24][17] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_2/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_2/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_2/n3 ), .ZN(
        \dp/ex_stage/alu/adder/carries [6]) );
  AOI21_X1 \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_3/U2  ( .B1(
        \dp/ex_stage/alu/adder/SparseTree/prop[20][17] ), .B2(
        \dp/ex_stage/alu/adder/carries [4]), .A(
        \dp/ex_stage/alu/adder/SparseTree/gen[20][17] ), .ZN(
        \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_3/n3 ) );
  INV_X1 \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_3/U1  ( .A(
        \dp/ex_stage/alu/adder/SparseTree/G_2n_0_5_3/n3 ), .ZN(
        \dp/ex_stage/alu/adder/carries [5]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [3]), .B(\dp/ex_stage/alu/adder/B_xor[3] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [2]), .B(\dp/ex_stage/alu/adder/B_xor[2] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [1]), .B(\dp/ex_stage/alu/adder/B_xor[1] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/alu/shifter/N202 ), .B(
        \dp/ex_stage/alu/adder/B_xor[0] ), .CI(1'b0), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA0/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 [0]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [3]), .B(\dp/ex_stage/alu/adder/B_xor[3] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [2]), .B(\dp/ex_stage/alu/adder/B_xor[2] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [1]), .B(\dp/ex_stage/alu/adder/B_xor[1] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/alu/shifter/N202 ), .B(
        \dp/ex_stage/alu/adder/B_xor[0] ), .CI(1'b1), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/RCA1/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 [0]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U9  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 [0]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 [0]), .B2(
        \dp/ex_stage/alu/adder/carries [0]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n9 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U8  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n9 ), .ZN(
        \dp/ex_stage/alu/adder_out [0]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U7  ( .A(
        \dp/ex_stage/alu/adder/carries [0]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n5 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U6  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 [1]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 [1]), .B2(
        \dp/ex_stage/alu/adder/carries [0]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n8 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U5  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n8 ), .ZN(
        \dp/ex_stage/alu/adder_out [1]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U4  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 [2]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 [2]), .B2(
        \dp/ex_stage/alu/adder/carries [0]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n7 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U3  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n7 ), .ZN(
        \dp/ex_stage/alu/adder_out [2]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U2  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out0 [3]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/carries [0]), .B2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/rca_out1 [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n6 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/U1  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_0/Mux/n6 ), .ZN(
        \dp/ex_stage/alu/adder_out [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [7]), .B(\dp/ex_stage/alu/adder/B_xor[7] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [6]), .B(\dp/ex_stage/alu/adder/B_xor[6] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [5]), .B(\dp/ex_stage/alu/adder/B_xor[5] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [4]), .B(\dp/ex_stage/alu/adder/B_xor[4] ), 
        .CI(1'b0), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA0/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 [0]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [7]), .B(\dp/ex_stage/alu/adder/B_xor[7] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [6]), .B(\dp/ex_stage/alu/adder/B_xor[6] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [5]), .B(\dp/ex_stage/alu/adder/B_xor[5] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [4]), .B(\dp/ex_stage/alu/adder/B_xor[4] ), 
        .CI(1'b1), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/RCA1/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 [0]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U9  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 [0]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 [0]), .B2(
        \dp/ex_stage/alu/adder/carries [1]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n10 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U8  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n10 ), .ZN(
        \dp/ex_stage/alu/adder_out [4]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U7  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 [1]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 [1]), .B2(
        \dp/ex_stage/alu/adder/carries [1]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n11 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U6  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n11 ), .ZN(
        \dp/ex_stage/alu/adder_out [5]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U5  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 [2]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 [2]), .B2(
        \dp/ex_stage/alu/adder/carries [1]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n12 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U4  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n12 ), .ZN(
        \dp/ex_stage/alu/adder_out [6]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U3  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out0 [3]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/carries [1]), .B2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/rca_out1 [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n13 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U2  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n13 ), .ZN(
        \dp/ex_stage/alu/adder_out [7]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/U1  ( .A(
        \dp/ex_stage/alu/adder/carries [1]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_1/Mux/n5 ) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [11]), .B(\dp/ex_stage/alu/adder/B_xor[11] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [10]), .B(\dp/ex_stage/alu/adder/B_xor[10] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [9]), .B(\dp/ex_stage/alu/adder/B_xor[9] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [8]), .B(\dp/ex_stage/alu/adder/B_xor[8] ), 
        .CI(1'b0), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA0/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 [0]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [11]), .B(\dp/ex_stage/alu/adder/B_xor[11] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [10]), .B(\dp/ex_stage/alu/adder/B_xor[10] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [9]), .B(\dp/ex_stage/alu/adder/B_xor[9] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [8]), .B(\dp/ex_stage/alu/adder/B_xor[8] ), 
        .CI(1'b1), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/RCA1/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 [0]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U9  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 [0]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 [0]), .B2(
        \dp/ex_stage/alu/adder/carries [2]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n10 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U8  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n10 ), .ZN(
        \dp/ex_stage/alu/adder_out [8]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U7  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 [1]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 [1]), .B2(
        \dp/ex_stage/alu/adder/carries [2]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n11 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U6  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n11 ), .ZN(
        \dp/ex_stage/alu/adder_out [9]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U5  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 [2]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 [2]), .B2(
        \dp/ex_stage/alu/adder/carries [2]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n12 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U4  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n12 ), .ZN(
        \dp/ex_stage/alu/adder_out [10]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U3  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out0 [3]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/carries [2]), .B2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/rca_out1 [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n13 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U2  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n13 ), .ZN(
        \dp/ex_stage/alu/adder_out [11]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/U1  ( .A(
        \dp/ex_stage/alu/adder/carries [2]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_2/Mux/n5 ) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [15]), .B(\dp/ex_stage/alu/adder/B_xor[15] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/alu/n37 ), .B(\dp/ex_stage/alu/adder/B_xor[14] ), .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [13]), .B(\dp/ex_stage/alu/adder/B_xor[13] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/alu/n34 ), .B(\dp/ex_stage/alu/adder/B_xor[12] ), .CI(
        1'b0), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA0/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 [0]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [15]), .B(\dp/ex_stage/alu/adder/B_xor[15] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/alu/n37 ), .B(\dp/ex_stage/alu/adder/B_xor[14] ), .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [13]), .B(\dp/ex_stage/alu/adder/B_xor[13] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/alu/n34 ), .B(\dp/ex_stage/alu/adder/B_xor[12] ), .CI(
        1'b1), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/RCA1/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 [0]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U9  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 [0]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 [0]), .B2(
        \dp/ex_stage/alu/adder/carries [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n10 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U8  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n10 ), .ZN(
        \dp/ex_stage/alu/adder_out [12]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U7  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n13 ), .ZN(
        \dp/ex_stage/alu/adder_out [15]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U6  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 [1]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 [1]), .B2(
        \dp/ex_stage/alu/adder/carries [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n11 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U5  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 [3]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/carries [3]), .B2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n13 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U4  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n11 ), .ZN(
        \dp/ex_stage/alu/adder_out [13]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U3  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n12 ), .ZN(
        \dp/ex_stage/alu/adder_out [14]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U2  ( .A(
        \dp/ex_stage/alu/adder/carries [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n5 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/U1  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out0 [2]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/rca_out1 [2]), .B2(
        \dp/ex_stage/alu/adder/carries [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_3/Mux/n12 ) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [19]), .B(\dp/ex_stage/alu/adder/B_xor[19] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [18]), .B(\dp/ex_stage/alu/adder/B_xor[18] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [17]), .B(\dp/ex_stage/alu/adder/B_xor[17] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [16]), .B(\dp/ex_stage/alu/adder/B_xor[16] ), 
        .CI(1'b0), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA0/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 [0]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [19]), .B(\dp/ex_stage/alu/adder/B_xor[19] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [18]), .B(\dp/ex_stage/alu/adder/B_xor[18] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [17]), .B(\dp/ex_stage/alu/adder/B_xor[17] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [16]), .B(\dp/ex_stage/alu/adder/B_xor[16] ), 
        .CI(1'b1), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/RCA1/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 [0]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U9  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 [3]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/carries [4]), .B2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n13 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U8  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 [0]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 [0]), .B2(
        \dp/ex_stage/alu/adder/carries [4]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n10 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U7  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n13 ), .ZN(
        \dp/ex_stage/alu/adder_out [19]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U6  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 [1]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 [1]), .B2(
        \dp/ex_stage/alu/adder/carries [4]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n11 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U5  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out0 [2]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/rca_out1 [2]), .B2(
        \dp/ex_stage/alu/adder/carries [4]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n12 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U4  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n11 ), .ZN(
        \dp/ex_stage/alu/adder_out [17]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U3  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n12 ), .ZN(
        \dp/ex_stage/alu/adder_out [18]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U2  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n10 ), .ZN(
        \dp/ex_stage/alu/adder_out [16]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/U1  ( .A(
        \dp/ex_stage/alu/adder/carries [4]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_4/Mux/n5 ) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/alu/n45 ), .B(\dp/ex_stage/alu/adder/B_xor[23] ), .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/alu/n43 ), .B(\dp/ex_stage/alu/adder/B_xor[22] ), .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [21]), .B(\dp/ex_stage/alu/adder/B_xor[21] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [20]), .B(\dp/ex_stage/alu/adder/B_xor[20] ), 
        .CI(1'b0), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA0/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 [0]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/alu/n45 ), .B(\dp/ex_stage/alu/adder/B_xor[23] ), .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/alu/n43 ), .B(\dp/ex_stage/alu/adder/B_xor[22] ), .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [21]), .B(\dp/ex_stage/alu/adder/B_xor[21] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [20]), .B(\dp/ex_stage/alu/adder/B_xor[20] ), 
        .CI(1'b1), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/RCA1/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 [0]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U9  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 [0]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 [0]), .B2(
        \dp/ex_stage/alu/adder/carries [5]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n10 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U8  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n13 ), .ZN(
        \dp/ex_stage/alu/adder_out [23]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U7  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 [1]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 [1]), .B2(
        \dp/ex_stage/alu/adder/carries [5]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n11 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U6  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 [3]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/carries [5]), .B2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n13 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U5  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n10 ), .ZN(
        \dp/ex_stage/alu/adder_out [20]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U4  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n11 ), .ZN(
        \dp/ex_stage/alu/adder_out [21]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U3  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n12 ), .ZN(
        \dp/ex_stage/alu/adder_out [22]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U2  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out0 [2]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/rca_out1 [2]), .B2(
        \dp/ex_stage/alu/adder/carries [5]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n12 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/U1  ( .A(
        \dp/ex_stage/alu/adder/carries [5]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_5/Mux/n5 ) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [27]), .B(\dp/ex_stage/alu/adder/B_xor[27] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [26]), .B(\dp/ex_stage/alu/adder/B_xor[26] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [25]), .B(\dp/ex_stage/alu/adder/B_xor[25] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [24]), .B(\dp/ex_stage/alu/adder/B_xor[24] ), 
        .CI(1'b0), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA0/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 [0]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/muxA_out [27]), .B(\dp/ex_stage/alu/adder/B_xor[27] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [26]), .B(\dp/ex_stage/alu/adder/B_xor[26] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [25]), .B(\dp/ex_stage/alu/adder/B_xor[25] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [24]), .B(\dp/ex_stage/alu/adder/B_xor[24] ), 
        .CI(1'b1), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/RCA1/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 [0]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U9  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 [0]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 [0]), .B2(
        \dp/ex_stage/alu/adder/carries [6]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n10 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U8  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 [3]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/carries [6]), .B2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n13 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U7  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n13 ), .ZN(
        \dp/ex_stage/alu/adder_out [27]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U6  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 [1]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 [1]), .B2(
        \dp/ex_stage/alu/adder/carries [6]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n11 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U5  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out0 [2]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/rca_out1 [2]), .B2(
        \dp/ex_stage/alu/adder/carries [6]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n12 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U4  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n10 ), .ZN(
        \dp/ex_stage/alu/adder_out [24]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U3  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n11 ), .ZN(
        \dp/ex_stage/alu/adder_out [25]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U2  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n12 ), .ZN(
        \dp/ex_stage/alu/adder_out [26]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/U1  ( .A(
        \dp/ex_stage/alu/adder/carries [6]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_6/Mux/n5 ) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/alu/shifter/N136 ), .B(
        \dp/ex_stage/alu/adder/B_xor[31] ), .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [30]), .B(\dp/ex_stage/alu/adder/B_xor[30] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [29]), .B(\dp/ex_stage/alu/adder/B_xor[29] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [28]), .B(\dp/ex_stage/alu/adder/B_xor[28] ), 
        .CI(1'b0), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA0/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 [0]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/U1_3  ( 
        .A(\dp/ex_stage/alu/shifter/N136 ), .B(
        \dp/ex_stage/alu/adder/B_xor[31] ), .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[3] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/Co ), .S(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 [3]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/U1_2  ( 
        .A(\dp/ex_stage/muxA_out [30]), .B(\dp/ex_stage/alu/adder/B_xor[30] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[2] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[3] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 [2]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/U1_1  ( 
        .A(\dp/ex_stage/muxA_out [29]), .B(\dp/ex_stage/alu/adder/B_xor[29] ), 
        .CI(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[1] ), .CO(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[2] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 [1]) );
  FA_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/U1_0  ( 
        .A(\dp/ex_stage/muxA_out [28]), .B(\dp/ex_stage/alu/adder/B_xor[28] ), 
        .CI(1'b1), .CO(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/RCA1/add_1_root_add_27_2/carry[1] ), .S(\dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 [0]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U9  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 [0]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 [0]), .B2(
        \dp/ex_stage/alu/adder/carries [7]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n10 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U8  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 [3]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/carries [7]), .B2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 [3]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n13 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U7  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n13 ), .ZN(
        \dp/ex_stage/alu/adder_out [31]) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U6  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 [1]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 [1]), .B2(
        \dp/ex_stage/alu/adder/carries [7]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n11 ) );
  AOI22_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U5  ( .A1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out0 [2]), .A2(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n5 ), .B1(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/rca_out1 [2]), .B2(
        \dp/ex_stage/alu/adder/carries [7]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n12 ) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U4  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n10 ), .ZN(
        \dp/ex_stage/alu/adder_out [28]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U3  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n11 ), .ZN(
        \dp/ex_stage/alu/adder_out [29]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U2  ( .A(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n12 ), .ZN(
        \dp/ex_stage/alu/adder_out [30]) );
  INV_X1 \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/U1  ( .A(
        \dp/ex_stage/alu/adder/carries [7]), .ZN(
        \dp/ex_stage/alu/adder/SumGen/CS_Bn_7/Mux/n5 ) );
  CLKBUF_X1 \dp/ex_stage/alu/shifter/U133  ( .A(\dp/ex_stage/alu/n31 ), .Z(
        \dp/ex_stage/alu/shifter/n99 ) );
  CLKBUF_X1 \dp/ex_stage/alu/shifter/U132  ( .A(\dp/ex_stage/alu/n31 ), .Z(
        \dp/ex_stage/alu/shifter/n98 ) );
  CLKBUF_X1 \dp/ex_stage/alu/shifter/U131  ( .A(\dp/ex_stage/alu/n31 ), .Z(
        \dp/ex_stage/alu/shifter/n97 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/U130  ( .A1(\dp/ex_stage/alu/shifter/n101 ), 
        .A2(1'b1), .ZN(\dp/ex_stage/alu/shifter/n26 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/U129  ( .A1(\dp/ex_stage/alu/n208 ), .A2(
        1'b1), .ZN(\dp/ex_stage/alu/shifter/n28 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/U128  ( .A1(\dp/ex_stage/alu/shift_arith_i ), .A2(1'b1), .ZN(\dp/ex_stage/alu/shifter/n91 ) );
  INV_X1 \dp/ex_stage/alu/shifter/U127  ( .A(1'b1), .ZN(
        \dp/ex_stage/alu/shifter/n100 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/U126  ( .A1(\dp/ex_stage/alu/shifter/n100 ), 
        .A2(\dp/ex_stage/alu/shift_arith_i ), .ZN(
        \dp/ex_stage/alu/shifter/n92 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U125  ( .A(\dp/ex_stage/alu/shifter/n28 ), 
        .Z(\dp/ex_stage/alu/shifter/n3 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U124  ( .A(\dp/ex_stage/alu/shifter/n26 ), 
        .Z(\dp/ex_stage/alu/shifter/n9 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U123  ( .A(\dp/ex_stage/alu/shifter/n26 ), 
        .Z(\dp/ex_stage/alu/shifter/n7 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U122  ( .A(\dp/ex_stage/alu/shifter/n26 ), 
        .Z(\dp/ex_stage/alu/shifter/n8 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U121  ( .A(\dp/ex_stage/alu/shifter/n28 ), 
        .Z(\dp/ex_stage/alu/shifter/n1 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U120  ( .A(\dp/ex_stage/alu/shifter/n28 ), 
        .Z(\dp/ex_stage/alu/shifter/n2 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/U119  ( .A1(\dp/ex_stage/alu/n208 ), .A2(
        \dp/ex_stage/alu/shifter/n92 ), .ZN(\dp/ex_stage/alu/shifter/n23 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U118  ( .A1(
        \dp/ex_stage/alu/shifter/N202 ), .A2(\dp/ex_stage/alu/shifter/n94 ), 
        .B1(\dp/ex_stage/alu/shifter/N105 ), .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N137 ), .C2(\dp/ex_stage/alu/shifter/n10 ), 
        .ZN(\dp/ex_stage/alu/shifter/n90 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U117  ( .A1(\dp/ex_stage/alu/shifter/N39 ), .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N234 ), .B2(
        \dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N7 ), .C2(
        \dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n89 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U116  ( .A1(\dp/ex_stage/alu/shifter/n89 ), 
        .A2(\dp/ex_stage/alu/shifter/n90 ), .ZN(
        \dp/ex_stage/alu/shifter_out [0]) );
  AND2_X1 \dp/ex_stage/alu/shifter/U115  ( .A1(\dp/ex_stage/alu/shifter/n91 ), 
        .A2(\dp/ex_stage/alu/shifter/n101 ), .ZN(\dp/ex_stage/alu/shifter/n25 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/U114  ( .A1(\dp/ex_stage/alu/shifter/n92 ), 
        .A2(\dp/ex_stage/alu/shifter/n101 ), .ZN(\dp/ex_stage/alu/shifter/n24 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/U113  ( .A1(\dp/ex_stage/alu/n208 ), .A2(
        \dp/ex_stage/alu/shifter/n91 ), .ZN(\dp/ex_stage/alu/shifter/n27 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U112  ( .A1(\dp/ex_stage/alu/shifter/n37 ), 
        .A2(\dp/ex_stage/alu/shifter/n38 ), .ZN(
        \dp/ex_stage/alu/shifter_out [4]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U111  ( .A1(\dp/ex_stage/alu/shifter/n29 ), 
        .A2(\dp/ex_stage/alu/shifter/n30 ), .ZN(
        \dp/ex_stage/alu/shifter_out [8]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U110  ( .A1(\dp/ex_stage/alu/shifter/n83 ), 
        .A2(\dp/ex_stage/alu/shifter/n84 ), .ZN(
        \dp/ex_stage/alu/shifter_out [12]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U109  ( .A1(
        \dp/ex_stage/alu/shifter/N233 ), .A2(\dp/ex_stage/alu/shifter/n96 ), 
        .B1(\dp/ex_stage/alu/shifter/N136 ), .B2(\dp/ex_stage/alu/shifter/n93 ), .C1(\dp/ex_stage/alu/shifter/N168 ), .C2(\dp/ex_stage/alu/shifter/n12 ), 
        .ZN(\dp/ex_stage/alu/shifter/n42 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U108  ( .A1(\dp/ex_stage/alu/shifter/N54 ), .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N249 ), .B2(
        \dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N22 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n77 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U107  ( .A1(\dp/ex_stage/alu/shifter/n77 ), 
        .A2(\dp/ex_stage/alu/shifter/n78 ), .ZN(
        \dp/ex_stage/alu/shifter_out [15]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U106  ( .A1(\dp/ex_stage/alu/shifter/N62 ), .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N257 ), .B2(
        \dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N30 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n59 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U105  ( .A1(\dp/ex_stage/alu/shifter/n59 ), 
        .A2(\dp/ex_stage/alu/shifter/n60 ), .ZN(
        \dp/ex_stage/alu/shifter_out [23]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U104  ( .A1(\dp/ex_stage/alu/shifter/N66 ), .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N261 ), .B2(
        \dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N34 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n51 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U103  ( .A1(\dp/ex_stage/alu/shifter/n51 ), 
        .A2(\dp/ex_stage/alu/shifter/n52 ), .ZN(
        \dp/ex_stage/alu/shifter_out [27]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U102  ( .A1(\dp/ex_stage/alu/shifter/N70 ), .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N265 ), .B2(
        \dp/ex_stage/alu/shifter/n6 ), .C1(\dp/ex_stage/alu/shifter/N38 ), 
        .C2(\dp/ex_stage/alu/shifter/n3 ), .ZN(\dp/ex_stage/alu/shifter/n41 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U101  ( .A1(\dp/ex_stage/alu/shifter/n41 ), 
        .A2(\dp/ex_stage/alu/shifter/n42 ), .ZN(
        \dp/ex_stage/alu/shifter_out [31]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U100  ( .A1(\dp/ex_stage/alu/shifter/N58 ), .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N253 ), .B2(
        \dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N26 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n69 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U99  ( .A1(\dp/ex_stage/alu/shifter/n69 ), 
        .A2(\dp/ex_stage/alu/shifter/n70 ), .ZN(
        \dp/ex_stage/alu/shifter_out [19]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U98  ( .A1(\dp/ex_stage/alu/shifter/N47 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N242 ), 
        .B2(\dp/ex_stage/alu/shifter/n6 ), .C1(\dp/ex_stage/alu/shifter/N15 ), 
        .C2(\dp/ex_stage/alu/shifter/n3 ), .ZN(\dp/ex_stage/alu/shifter/n29 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U97  ( .A1(\dp/ex_stage/alu/shifter/N48 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N243 ), 
        .B2(\dp/ex_stage/alu/shifter/n6 ), .C1(\dp/ex_stage/alu/shifter/N16 ), 
        .C2(\dp/ex_stage/alu/shifter/n3 ), .ZN(\dp/ex_stage/alu/shifter/n21 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U96  ( .A1(\dp/ex_stage/alu/shifter/N49 ), 
        .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N244 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N17 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n87 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U95  ( .A1(\dp/ex_stage/alu/shifter/N50 ), 
        .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N245 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N18 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n85 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U94  ( .A1(\dp/ex_stage/alu/shifter/N51 ), 
        .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N246 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N19 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n83 )
         );
  INV_X1 \dp/ex_stage/alu/shifter/U93  ( .A(\dp/ex_stage/alu/n208 ), .ZN(
        \dp/ex_stage/alu/shifter/n101 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U92  ( .A1(\dp/ex_stage/alu/shifter/N45 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N240 ), 
        .B2(\dp/ex_stage/alu/shifter/n6 ), .C1(\dp/ex_stage/alu/shifter/N13 ), 
        .C2(\dp/ex_stage/alu/shifter/n3 ), .ZN(\dp/ex_stage/alu/shifter/n33 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U91  ( .A1(\dp/ex_stage/alu/shifter/N46 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N241 ), 
        .B2(\dp/ex_stage/alu/shifter/n6 ), .C1(\dp/ex_stage/alu/shifter/N14 ), 
        .C2(\dp/ex_stage/alu/shifter/n3 ), .ZN(\dp/ex_stage/alu/shifter/n31 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U90  ( .A1(\dp/ex_stage/alu/shifter/N41 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N236 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N9 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n45 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U89  ( .A1(\dp/ex_stage/alu/shifter/N42 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N237 ), 
        .B2(\dp/ex_stage/alu/shifter/n6 ), .C1(\dp/ex_stage/alu/shifter/N10 ), 
        .C2(\dp/ex_stage/alu/shifter/n3 ), .ZN(\dp/ex_stage/alu/shifter/n39 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U88  ( .A1(\dp/ex_stage/alu/shifter/N43 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N238 ), 
        .B2(\dp/ex_stage/alu/shifter/n6 ), .C1(\dp/ex_stage/alu/shifter/N11 ), 
        .C2(\dp/ex_stage/alu/shifter/n3 ), .ZN(\dp/ex_stage/alu/shifter/n37 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U87  ( .A1(\dp/ex_stage/alu/shifter/N44 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N239 ), 
        .B2(\dp/ex_stage/alu/shifter/n6 ), .C1(\dp/ex_stage/alu/shifter/N12 ), 
        .C2(\dp/ex_stage/alu/shifter/n3 ), .ZN(\dp/ex_stage/alu/shifter/n35 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U86  ( .A1(\dp/ex_stage/alu/shifter/n67 ), 
        .A2(\dp/ex_stage/alu/shifter/n68 ), .ZN(
        \dp/ex_stage/alu/shifter_out [1]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U85  ( .A1(\dp/ex_stage/alu/shifter/n45 ), 
        .A2(\dp/ex_stage/alu/shifter/n46 ), .ZN(
        \dp/ex_stage/alu/shifter_out [2]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U84  ( .A1(\dp/ex_stage/alu/shifter/n39 ), 
        .A2(\dp/ex_stage/alu/shifter/n40 ), .ZN(
        \dp/ex_stage/alu/shifter_out [3]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U83  ( .A1(\dp/ex_stage/alu/shifter/n35 ), 
        .A2(\dp/ex_stage/alu/shifter/n36 ), .ZN(
        \dp/ex_stage/alu/shifter_out [5]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U82  ( .A1(\dp/ex_stage/alu/shifter/n33 ), 
        .A2(\dp/ex_stage/alu/shifter/n34 ), .ZN(
        \dp/ex_stage/alu/shifter_out [6]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U81  ( .A1(\dp/ex_stage/alu/shifter/n31 ), 
        .A2(\dp/ex_stage/alu/shifter/n32 ), .ZN(
        \dp/ex_stage/alu/shifter_out [7]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U80  ( .A1(\dp/ex_stage/alu/shifter/n21 ), 
        .A2(\dp/ex_stage/alu/shifter/n22 ), .ZN(
        \dp/ex_stage/alu/shifter_out [9]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U79  ( .A1(\dp/ex_stage/alu/shifter/N56 ), 
        .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N251 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N24 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n73 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U78  ( .A1(\dp/ex_stage/alu/shifter/n73 ), 
        .A2(\dp/ex_stage/alu/shifter/n74 ), .ZN(
        \dp/ex_stage/alu/shifter_out [17]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U77  ( .A1(\dp/ex_stage/alu/shifter/N57 ), 
        .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N252 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N25 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n71 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U76  ( .A1(\dp/ex_stage/alu/shifter/n71 ), 
        .A2(\dp/ex_stage/alu/shifter/n72 ), .ZN(
        \dp/ex_stage/alu/shifter_out [18]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U75  ( .A1(\dp/ex_stage/alu/shifter/N59 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N254 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N27 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n65 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U74  ( .A1(\dp/ex_stage/alu/shifter/n65 ), 
        .A2(\dp/ex_stage/alu/shifter/n66 ), .ZN(
        \dp/ex_stage/alu/shifter_out [20]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U73  ( .A1(\dp/ex_stage/alu/shifter/N60 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N255 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N28 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n63 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U72  ( .A1(\dp/ex_stage/alu/shifter/n63 ), 
        .A2(\dp/ex_stage/alu/shifter/n64 ), .ZN(
        \dp/ex_stage/alu/shifter_out [21]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U71  ( .A1(\dp/ex_stage/alu/shifter/N61 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N256 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N29 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n61 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U70  ( .A1(\dp/ex_stage/alu/shifter/n61 ), 
        .A2(\dp/ex_stage/alu/shifter/n62 ), .ZN(
        \dp/ex_stage/alu/shifter_out [22]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U69  ( .A1(\dp/ex_stage/alu/shifter/N63 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N258 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N31 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n57 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U68  ( .A1(\dp/ex_stage/alu/shifter/n57 ), 
        .A2(\dp/ex_stage/alu/shifter/n58 ), .ZN(
        \dp/ex_stage/alu/shifter_out [24]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U67  ( .A1(\dp/ex_stage/alu/shifter/N64 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N259 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N32 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n55 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U66  ( .A1(\dp/ex_stage/alu/shifter/n55 ), 
        .A2(\dp/ex_stage/alu/shifter/n56 ), .ZN(
        \dp/ex_stage/alu/shifter_out [25]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U65  ( .A1(\dp/ex_stage/alu/shifter/N65 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N260 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N33 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n53 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U64  ( .A1(\dp/ex_stage/alu/shifter/n53 ), 
        .A2(\dp/ex_stage/alu/shifter/n54 ), .ZN(
        \dp/ex_stage/alu/shifter_out [26]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U63  ( .A1(\dp/ex_stage/alu/shifter/N67 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N262 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N35 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n49 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U62  ( .A1(\dp/ex_stage/alu/shifter/n49 ), 
        .A2(\dp/ex_stage/alu/shifter/n50 ), .ZN(
        \dp/ex_stage/alu/shifter_out [28]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U61  ( .A1(\dp/ex_stage/alu/shifter/N68 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N263 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N36 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n47 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U60  ( .A1(\dp/ex_stage/alu/shifter/n47 ), 
        .A2(\dp/ex_stage/alu/shifter/n48 ), .ZN(
        \dp/ex_stage/alu/shifter_out [29]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U59  ( .A1(\dp/ex_stage/alu/shifter/N69 ), 
        .A2(\dp/ex_stage/alu/shifter/n9 ), .B1(\dp/ex_stage/alu/shifter/N264 ), 
        .B2(\dp/ex_stage/alu/shifter/n5 ), .C1(\dp/ex_stage/alu/shifter/N37 ), 
        .C2(\dp/ex_stage/alu/shifter/n2 ), .ZN(\dp/ex_stage/alu/shifter/n43 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U58  ( .A1(\dp/ex_stage/alu/shifter/n43 ), 
        .A2(\dp/ex_stage/alu/shifter/n44 ), .ZN(
        \dp/ex_stage/alu/shifter_out [30]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U57  ( .A1(\dp/ex_stage/alu/shifter/n87 ), 
        .A2(\dp/ex_stage/alu/shifter/n88 ), .ZN(
        \dp/ex_stage/alu/shifter_out [10]) );
  NAND2_X1 \dp/ex_stage/alu/shifter/U56  ( .A1(\dp/ex_stage/alu/shifter/n85 ), 
        .A2(\dp/ex_stage/alu/shifter/n86 ), .ZN(
        \dp/ex_stage/alu/shifter_out [11]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U55  ( .A1(\dp/ex_stage/alu/shifter/N52 ), 
        .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N247 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N20 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n81 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U54  ( .A1(\dp/ex_stage/alu/shifter/n81 ), 
        .A2(\dp/ex_stage/alu/shifter/n82 ), .ZN(
        \dp/ex_stage/alu/shifter_out [13]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U53  ( .A1(\dp/ex_stage/alu/shifter/N53 ), 
        .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N248 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N21 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n79 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U52  ( .A1(\dp/ex_stage/alu/shifter/n79 ), 
        .A2(\dp/ex_stage/alu/shifter/n80 ), .ZN(
        \dp/ex_stage/alu/shifter_out [14]) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U51  ( .A1(\dp/ex_stage/alu/shifter/N55 ), 
        .A2(\dp/ex_stage/alu/shifter/n7 ), .B1(\dp/ex_stage/alu/shifter/N250 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N23 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n75 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/U50  ( .A1(\dp/ex_stage/alu/shifter/n75 ), 
        .A2(\dp/ex_stage/alu/shifter/n76 ), .ZN(
        \dp/ex_stage/alu/shifter_out [16]) );
  BUF_X1 \dp/ex_stage/alu/shifter/U49  ( .A(\dp/ex_stage/alu/shifter/n25 ), 
        .Z(\dp/ex_stage/alu/shifter/n12 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U48  ( .A(\dp/ex_stage/alu/shifter/n27 ), 
        .Z(\dp/ex_stage/alu/shifter/n6 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U47  ( .A(\dp/ex_stage/alu/shifter/n24 ), 
        .Z(\dp/ex_stage/alu/shifter/n93 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U46  ( .A(\dp/ex_stage/alu/shifter/n25 ), 
        .Z(\dp/ex_stage/alu/shifter/n10 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U45  ( .A(\dp/ex_stage/alu/shifter/n25 ), 
        .Z(\dp/ex_stage/alu/shifter/n11 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U44  ( .A1(\dp/ex_stage/alu/shifter/N218 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N121 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N153 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n76 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U43  ( .A1(\dp/ex_stage/alu/shifter/N219 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N122 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N154 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n74 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U42  ( .A1(\dp/ex_stage/alu/shifter/N220 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N123 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N155 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n72 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U41  ( .A1(\dp/ex_stage/alu/shifter/N221 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N124 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N156 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n70 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U40  ( .A1(\dp/ex_stage/alu/shifter/N222 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N125 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N157 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n66 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U39  ( .A1(\dp/ex_stage/alu/shifter/N223 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N126 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N158 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n64 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U38  ( .A1(\dp/ex_stage/alu/shifter/N224 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N127 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N159 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n62 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U37  ( .A1(\dp/ex_stage/alu/shifter/N225 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N128 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N160 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n60 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U36  ( .A1(\dp/ex_stage/alu/shifter/N226 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N129 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N161 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n58 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U35  ( .A1(\dp/ex_stage/alu/shifter/N227 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N130 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N162 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n56 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U34  ( .A1(\dp/ex_stage/alu/shifter/N228 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N131 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N163 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n54 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U33  ( .A(\dp/ex_stage/alu/shifter/n27 ), 
        .Z(\dp/ex_stage/alu/shifter/n4 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U32  ( .A(\dp/ex_stage/alu/shifter/n24 ), 
        .Z(\dp/ex_stage/alu/shifter/n19 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U31  ( .A(\dp/ex_stage/alu/shifter/n27 ), 
        .Z(\dp/ex_stage/alu/shifter/n5 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U30  ( .A(\dp/ex_stage/alu/shifter/n24 ), 
        .Z(\dp/ex_stage/alu/shifter/n20 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U29  ( .A(\dp/ex_stage/alu/shifter/n23 ), 
        .Z(\dp/ex_stage/alu/shifter/n96 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U28  ( .A(\dp/ex_stage/alu/shifter/n23 ), 
        .Z(\dp/ex_stage/alu/shifter/n94 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/U27  ( .A(\dp/ex_stage/alu/shifter/n23 ), 
        .Z(\dp/ex_stage/alu/shifter/n95 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U26  ( .A1(\dp/ex_stage/alu/shifter/N217 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N120 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N152 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n78 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U25  ( .A1(\dp/ex_stage/alu/shifter/N203 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N106 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N138 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n68 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U24  ( .A1(\dp/ex_stage/alu/shifter/N204 ), .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N107 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N139 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n46 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U23  ( .A1(\dp/ex_stage/alu/shifter/N205 ), .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N108 ), 
        .B2(\dp/ex_stage/alu/shifter/n93 ), .C1(\dp/ex_stage/alu/shifter/N140 ), .C2(\dp/ex_stage/alu/shifter/n12 ), .ZN(\dp/ex_stage/alu/shifter/n40 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U22  ( .A1(\dp/ex_stage/alu/shifter/N231 ), .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N134 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N166 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n48 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U21  ( .A1(\dp/ex_stage/alu/shifter/N232 ), .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N135 ), 
        .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N167 ), .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n44 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U20  ( .A1(\dp/ex_stage/alu/shifter/N213 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N116 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N148 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n86 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U19  ( .A1(\dp/ex_stage/alu/shifter/N40 ), 
        .A2(\dp/ex_stage/alu/shifter/n8 ), .B1(\dp/ex_stage/alu/shifter/N235 ), 
        .B2(\dp/ex_stage/alu/shifter/n4 ), .C1(\dp/ex_stage/alu/shifter/N8 ), 
        .C2(\dp/ex_stage/alu/shifter/n1 ), .ZN(\dp/ex_stage/alu/shifter/n67 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U18  ( .A1(\dp/ex_stage/alu/shifter/N206 ), .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N109 ), 
        .B2(\dp/ex_stage/alu/shifter/n93 ), .C1(\dp/ex_stage/alu/shifter/N141 ), .C2(\dp/ex_stage/alu/shifter/n12 ), .ZN(\dp/ex_stage/alu/shifter/n38 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U17  ( .A1(\dp/ex_stage/alu/shifter/N207 ), .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N110 ), 
        .B2(\dp/ex_stage/alu/shifter/n93 ), .C1(\dp/ex_stage/alu/shifter/N142 ), .C2(\dp/ex_stage/alu/shifter/n12 ), .ZN(\dp/ex_stage/alu/shifter/n36 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U16  ( .A1(\dp/ex_stage/alu/shifter/N208 ), .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N111 ), 
        .B2(\dp/ex_stage/alu/shifter/n93 ), .C1(\dp/ex_stage/alu/shifter/N143 ), .C2(\dp/ex_stage/alu/shifter/n12 ), .ZN(\dp/ex_stage/alu/shifter/n34 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U15  ( .A1(\dp/ex_stage/alu/shifter/N211 ), .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N114 ), 
        .B2(\dp/ex_stage/alu/shifter/n93 ), .C1(\dp/ex_stage/alu/shifter/N146 ), .C2(\dp/ex_stage/alu/shifter/n12 ), .ZN(\dp/ex_stage/alu/shifter/n22 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U14  ( .A1(\dp/ex_stage/alu/shifter/N212 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N115 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N147 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n88 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U13  ( .A1(\dp/ex_stage/alu/shifter/N215 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N118 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N150 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n82 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U10  ( .A1(\dp/ex_stage/alu/shifter/N214 ), .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N117 ), 
        .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N149 ), .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n84 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/U9  ( .A1(\dp/ex_stage/alu/shifter/N216 ), 
        .A2(\dp/ex_stage/alu/shifter/n94 ), .B1(\dp/ex_stage/alu/shifter/N119 ), .B2(\dp/ex_stage/alu/shifter/n19 ), .C1(\dp/ex_stage/alu/shifter/N151 ), 
        .C2(\dp/ex_stage/alu/shifter/n10 ), .ZN(\dp/ex_stage/alu/shifter/n80 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U8  ( .A1(\dp/ex_stage/alu/shifter/N229 ), 
        .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N132 ), .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N164 ), 
        .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n52 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U7  ( .A1(\dp/ex_stage/alu/shifter/N230 ), 
        .A2(\dp/ex_stage/alu/shifter/n95 ), .B1(\dp/ex_stage/alu/shifter/N133 ), .B2(\dp/ex_stage/alu/shifter/n20 ), .C1(\dp/ex_stage/alu/shifter/N165 ), 
        .C2(\dp/ex_stage/alu/shifter/n11 ), .ZN(\dp/ex_stage/alu/shifter/n50 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U6  ( .A1(\dp/ex_stage/alu/shifter/N209 ), 
        .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N112 ), .B2(\dp/ex_stage/alu/shifter/n93 ), .C1(\dp/ex_stage/alu/shifter/N144 ), 
        .C2(\dp/ex_stage/alu/shifter/n12 ), .ZN(\dp/ex_stage/alu/shifter/n32 )
         );
  AOI222_X1 \dp/ex_stage/alu/shifter/U5  ( .A1(\dp/ex_stage/alu/shifter/N210 ), 
        .A2(\dp/ex_stage/alu/shifter/n96 ), .B1(\dp/ex_stage/alu/shifter/N113 ), .B2(\dp/ex_stage/alu/shifter/n93 ), .C1(\dp/ex_stage/alu/shifter/N145 ), 
        .C2(\dp/ex_stage/alu/shifter/n12 ), .ZN(\dp/ex_stage/alu/shifter/n30 )
         );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U54  ( .A1(
        \dp/ex_stage/alu/shifter/N202 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n3 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][0] ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U53  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][0] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n6 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][0] ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U52  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][1] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n6 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][1] ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U51  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][0] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n9 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][0] ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U50  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][1] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n9 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][1] ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U49  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][2] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n9 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][2] ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U48  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][3] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n9 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][3] ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sll_48/U47  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][0] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n29 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sll_48/U46  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][1] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n28 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sll_48/U45  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][2] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n27 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sll_48/U44  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][3] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n26 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sll_48/U43  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][4] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n25 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sll_48/U42  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][5] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n24 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sll_48/U41  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][6] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n23 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sll_48/U40  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][7] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n22 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sll_48/U39  ( .A1(
        \dp/ex_stage/alu/shifter/n97 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n29 ), .ZN(
        \dp/ex_stage/alu/shifter/N234 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U38  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][10] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/N244 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U37  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][11] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/N245 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U36  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][12] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/N246 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U35  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][13] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/N247 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U34  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][14] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/N248 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U33  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][15] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/N249 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sll_48/U32  ( .A1(
        \dp/ex_stage/alu/shifter/n97 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n28 ), .ZN(
        \dp/ex_stage/alu/shifter/N235 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sll_48/U31  ( .A1(
        \dp/ex_stage/alu/shifter/n97 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n27 ), .ZN(
        \dp/ex_stage/alu/shifter/N236 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sll_48/U30  ( .A1(
        \dp/ex_stage/alu/shifter/n97 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n26 ), .ZN(
        \dp/ex_stage/alu/shifter/N237 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sll_48/U29  ( .A1(
        \dp/ex_stage/alu/shifter/n97 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n25 ), .ZN(
        \dp/ex_stage/alu/shifter/N238 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sll_48/U28  ( .A1(
        \dp/ex_stage/alu/shifter/n97 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n24 ), .ZN(
        \dp/ex_stage/alu/shifter/N239 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sll_48/U27  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n23 ), .ZN(
        \dp/ex_stage/alu/shifter/N240 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sll_48/U26  ( .A1(
        \dp/ex_stage/alu/shifter/n97 ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n22 ), .ZN(
        \dp/ex_stage/alu/shifter/N241 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U25  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][8] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/N242 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sll_48/U24  ( .A1(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][9] ), .A2(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/N243 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U23  ( .A(
        \dp/ex_stage/alu/shifter/n97 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n13 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U22  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n10 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U21  ( .A(\dp/ex_stage/alu/n27 ), 
        .ZN(\dp/ex_stage/alu/shifter/sll_48/n9 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U20  ( .A(\dp/ex_stage/muxB_out [0]), 
        .ZN(\dp/ex_stage/alu/shifter/sll_48/n3 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U19  ( .A(\dp/ex_stage/alu/n29 ), 
        .ZN(\dp/ex_stage/alu/shifter/sll_48/n11 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U18  ( .A(\dp/ex_stage/alu/n25 ), 
        .ZN(\dp/ex_stage/alu/shifter/sll_48/n6 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U17  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n3 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n1 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U16  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n3 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n2 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U15  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n9 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n7 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U14  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n9 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n8 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U13  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n6 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n4 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U12  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n6 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n5 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U11  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n29 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n14 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U10  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n28 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n18 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U9  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n27 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n16 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U8  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n26 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n20 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U7  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n25 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n15 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U6  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n24 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n19 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U5  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n23 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n17 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U4  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n22 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n21 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sll_48/U3  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/sll_48/n12 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_1  ( .A(
        \dp/ex_stage/muxA_out [1]), .B(\dp/ex_stage/alu/shifter/N202 ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_2  ( .A(
        \dp/ex_stage/muxA_out [2]), .B(\dp/ex_stage/muxA_out [1]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_3  ( .A(
        \dp/ex_stage/muxA_out [3]), .B(\dp/ex_stage/muxA_out [2]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_4  ( .A(
        \dp/ex_stage/muxA_out [4]), .B(\dp/ex_stage/muxA_out [3]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_5  ( .A(
        \dp/ex_stage/muxA_out [5]), .B(\dp/ex_stage/muxA_out [4]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_6  ( .A(
        \dp/ex_stage/muxA_out [6]), .B(\dp/ex_stage/muxA_out [5]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_7  ( .A(
        \dp/ex_stage/muxA_out [7]), .B(\dp/ex_stage/muxA_out [6]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_8  ( .A(
        \dp/ex_stage/muxA_out [8]), .B(\dp/ex_stage/muxA_out [7]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_9  ( .A(
        \dp/ex_stage/muxA_out [9]), .B(\dp/ex_stage/muxA_out [8]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_10  ( .A(
        \dp/ex_stage/muxA_out [10]), .B(\dp/ex_stage/muxA_out [9]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_11  ( .A(
        \dp/ex_stage/muxA_out [11]), .B(\dp/ex_stage/muxA_out [10]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_12  ( .A(\dp/ex_stage/alu/n34 ), 
        .B(\dp/ex_stage/muxA_out [11]), .S(\dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(\dp/ex_stage/alu/shifter/sll_48/ML_int[1][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_13  ( .A(
        \dp/ex_stage/muxA_out [13]), .B(\dp/ex_stage/alu/n34 ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_14  ( .A(\dp/ex_stage/alu/n37 ), 
        .B(\dp/ex_stage/muxA_out [13]), .S(\dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(\dp/ex_stage/alu/shifter/sll_48/ML_int[1][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_15  ( .A(
        \dp/ex_stage/muxA_out [15]), .B(\dp/ex_stage/alu/n37 ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_16  ( .A(
        \dp/ex_stage/muxA_out [16]), .B(\dp/ex_stage/muxA_out [15]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_17  ( .A(
        \dp/ex_stage/muxA_out [17]), .B(\dp/ex_stage/muxA_out [16]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_18  ( .A(
        \dp/ex_stage/muxA_out [18]), .B(\dp/ex_stage/muxA_out [17]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_19  ( .A(
        \dp/ex_stage/muxA_out [19]), .B(\dp/ex_stage/muxA_out [18]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_20  ( .A(
        \dp/ex_stage/muxA_out [20]), .B(\dp/ex_stage/muxA_out [19]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_21  ( .A(
        \dp/ex_stage/muxA_out [21]), .B(\dp/ex_stage/muxA_out [20]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_22  ( .A(\dp/ex_stage/alu/n43 ), 
        .B(\dp/ex_stage/muxA_out [21]), .S(\dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(\dp/ex_stage/alu/shifter/sll_48/ML_int[1][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_23  ( .A(\dp/ex_stage/alu/n45 ), 
        .B(\dp/ex_stage/alu/n43 ), .S(\dp/ex_stage/alu/shifter/sll_48/n2 ), 
        .Z(\dp/ex_stage/alu/shifter/sll_48/ML_int[1][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_24  ( .A(
        \dp/ex_stage/muxA_out [24]), .B(\dp/ex_stage/alu/n45 ), .S(
        \dp/ex_stage/muxB_out [0]), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_25  ( .A(
        \dp/ex_stage/muxA_out [25]), .B(\dp/ex_stage/muxA_out [24]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_26  ( .A(
        \dp/ex_stage/muxA_out [26]), .B(\dp/ex_stage/muxA_out [25]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_27  ( .A(
        \dp/ex_stage/muxA_out [27]), .B(\dp/ex_stage/muxA_out [26]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_28  ( .A(
        \dp/ex_stage/muxA_out [28]), .B(\dp/ex_stage/muxA_out [27]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_29  ( .A(
        \dp/ex_stage/muxA_out [29]), .B(\dp/ex_stage/muxA_out [28]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_30  ( .A(
        \dp/ex_stage/muxA_out [30]), .B(\dp/ex_stage/muxA_out [29]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n1 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_0_31  ( .A(
        \dp/ex_stage/alu/shifter/N136 ), .B(\dp/ex_stage/muxA_out [30]), .S(
        \dp/ex_stage/alu/shifter/sll_48/n2 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_2  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][2] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][0] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_3  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][3] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][1] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_4  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][4] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][2] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_5  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][5] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][3] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_6  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][6] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][4] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_7  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][7] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][5] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_8  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][8] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][6] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_9  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][9] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][7] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_10  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][10] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][8] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_11  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][11] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][9] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_12  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][12] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][10] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_13  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][13] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][11] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_14  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][14] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][12] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_15  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][15] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][13] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_16  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][16] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][14] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_17  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][17] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][15] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_18  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][18] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][16] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_19  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][19] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][17] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_20  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][20] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][18] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_21  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][21] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][19] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_22  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][22] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][20] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_23  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][23] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][21] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_24  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][24] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][22] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_25  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][25] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][23] ), .S(
        \dp/ex_stage/alu/n25 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_26  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][26] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][24] ), .S(
        \dp/ex_stage/alu/n25 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_27  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][27] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][25] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_28  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][28] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][26] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_29  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][29] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][27] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_30  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][30] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][28] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n4 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_1_31  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][31] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[1][29] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n5 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_4  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][4] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][0] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_5  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][5] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][1] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_6  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][6] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][2] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_7  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][7] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][3] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_8  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][8] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][4] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_9  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][9] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][5] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_10  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][10] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][6] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_11  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][11] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][7] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_12  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][12] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][8] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_13  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][13] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][9] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_14  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][14] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][10] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_15  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][15] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][11] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_16  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][16] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][12] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_17  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][17] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][13] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_18  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][18] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][14] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_19  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][19] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][15] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_20  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][20] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][16] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_21  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][21] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][17] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_22  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][22] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][18] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_23  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][23] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][19] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_24  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][24] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][20] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_25  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][25] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][21] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_26  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][26] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][22] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_27  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][27] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][23] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_28  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][28] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][24] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_29  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][29] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][25] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n7 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_30  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][30] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][26] ), .S(
        \dp/ex_stage/alu/n27 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_2_31  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][31] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[2][27] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n8 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_8  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][8] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][0] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_9  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][9] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][1] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_10  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][10] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][2] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_11  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][11] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][3] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_12  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][12] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][4] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_13  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][13] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][5] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_14  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][14] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][6] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_15  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][15] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][7] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_16  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][16] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][8] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_17  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][17] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][9] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_18  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][18] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][10] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_19  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][19] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][11] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_20  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][20] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][12] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_21  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][21] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][13] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_22  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][22] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][14] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_23  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][23] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][15] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_24  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][24] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][16] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_25  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][25] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][17] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_26  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][26] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][18] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_27  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][27] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][19] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_28  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][28] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][20] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_29  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][29] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][21] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_30  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][30] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][22] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_3_31  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][31] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[3][23] ), .S(
        \dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_16  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][16] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/n14 ), .S(
        \dp/ex_stage/alu/shifter/n97 ), .Z(\dp/ex_stage/alu/shifter/N250 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_17  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][17] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/n18 ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N251 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_18  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][18] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/n16 ), .S(
        \dp/ex_stage/alu/shifter/n97 ), .Z(\dp/ex_stage/alu/shifter/N252 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_19  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][19] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/n20 ), .S(
        \dp/ex_stage/alu/shifter/n97 ), .Z(\dp/ex_stage/alu/shifter/N253 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_20  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][20] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/n15 ), .S(
        \dp/ex_stage/alu/shifter/n97 ), .Z(\dp/ex_stage/alu/shifter/N254 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_21  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][21] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/n19 ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N255 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_22  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][22] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/n17 ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N256 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_23  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][23] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/n21 ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N257 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_24  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][24] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][8] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N258 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_25  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][25] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][9] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N259 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_26  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][26] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][10] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N260 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_27  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][27] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][11] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N261 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_28  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][28] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][12] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N262 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_29  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][29] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][13] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N263 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_30  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][30] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][14] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N264 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sll_48/M1_4_31  ( .A(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][31] ), .B(
        \dp/ex_stage/alu/shifter/sll_48/ML_int[4][15] ), .S(
        \dp/ex_stage/alu/shifter/sll_48/n12 ), .Z(
        \dp/ex_stage/alu/shifter/N265 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sla_46/U221  ( .A1(\dp/ex_stage/alu/n25 ), 
        .A2(\dp/ex_stage/alu/shifter/sla_46/n13 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n91 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sla_46/U220  ( .A1(
        \dp/ex_stage/muxB_out [0]), .A2(\dp/ex_stage/alu/n25 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n92 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sla_46/U219  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n13 ), .A2(\dp/ex_stage/alu/n25 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n94 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sla_46/U218  ( .A1(
        \dp/ex_stage/muxB_out [0]), .A2(\dp/ex_stage/alu/n25 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n95 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U217  ( .A1(
        \dp/ex_stage/muxA_out [5]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/muxA_out [6]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n189 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U216  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n42 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n41 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n189 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n151 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U215  ( .A1(
        \dp/ex_stage/muxA_out [9]), .A2(\dp/ex_stage/alu/shifter/sla_46/n9 ), 
        .B1(\dp/ex_stage/muxA_out [10]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n12 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n188 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U214  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n3 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n47 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n46 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n188 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n150 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sla_46/U213  ( .A1(\dp/ex_stage/alu/n29 ), 
        .A2(\dp/ex_stage/alu/shifter/sla_46/n14 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n133 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U212  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .A2(\dp/ex_stage/muxA_out [2]), 
        .B1(\dp/ex_stage/muxA_out [1]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n9 ), .C1(
        \dp/ex_stage/alu/shifter/N202 ), .C2(\dp/ex_stage/alu/n25 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n187 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sla_46/U211  ( .A1(\dp/ex_stage/alu/n29 ), 
        .A2(\dp/ex_stage/alu/shifter/N202 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n154 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sla_46/U210  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n14 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n154 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n135 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sla_46/U209  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n133 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n32 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n135 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n186 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U208  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n151 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n150 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n30 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n121 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sla_46/U207  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n17 ), .A2(
        \dp/ex_stage/alu/shifter/N202 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n76 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U206  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n17 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n121 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N212 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U205  ( .A1(
        \dp/ex_stage/muxA_out [6]), .A2(\dp/ex_stage/alu/shifter/sla_46/n9 ), 
        .B1(\dp/ex_stage/muxA_out [7]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n12 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n185 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U204  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n3 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n43 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n6 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n42 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n185 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n147 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U203  ( .A1(
        \dp/ex_stage/muxA_out [10]), .A2(\dp/ex_stage/alu/shifter/sla_46/n9 ), 
        .B1(\dp/ex_stage/muxA_out [11]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n12 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n184 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U202  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n3 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n49 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n6 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n47 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n184 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n145 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U201  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n9 ), .A2(\dp/ex_stage/muxA_out [2]), 
        .B1(\dp/ex_stage/muxA_out [3]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n12 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n183 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U200  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n19 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n3 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n39 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n183 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n146 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sla_46/U199  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n133 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n146 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n135 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n182 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U198  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n147 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n145 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n33 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n116 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U197  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n17 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n116 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N213 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U196  ( .A1(
        \dp/ex_stage/muxA_out [7]), .A2(\dp/ex_stage/alu/shifter/sla_46/n9 ), 
        .B1(\dp/ex_stage/muxA_out [8]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n12 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n181 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U195  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n3 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n45 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n6 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n43 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n181 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n141 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U194  ( .A1(
        \dp/ex_stage/muxA_out [11]), .A2(\dp/ex_stage/alu/shifter/sla_46/n9 ), 
        .B1(\dp/ex_stage/alu/n34 ), .B2(\dp/ex_stage/alu/shifter/sla_46/n12 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n180 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U193  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n3 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n50 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n6 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n49 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n180 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n139 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U192  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n9 ), .A2(\dp/ex_stage/muxA_out [3]), 
        .B1(\dp/ex_stage/muxA_out [4]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n12 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n179 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U191  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n3 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n40 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n19 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n179 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n140 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sla_46/U190  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n133 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n140 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n135 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n178 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U189  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n141 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n139 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n34 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n109 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U188  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n17 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n109 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N214 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sla_46/U187  ( .A(
        \dp/ex_stage/alu/shifter/N202 ), .B(\dp/ex_stage/muxA_out [1]), .S(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n134 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sla_46/U186  ( .A1(\dp/ex_stage/alu/n27 ), 
        .A2(\dp/ex_stage/alu/n29 ), .ZN(\dp/ex_stage/alu/shifter/sla_46/n170 )
         );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U185  ( .A1(
        \dp/ex_stage/muxA_out [4]), .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), 
        .B1(\dp/ex_stage/muxA_out [5]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n177 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U184  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n41 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n6 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n40 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n177 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n128 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U183  ( .A1(
        \dp/ex_stage/muxA_out [8]), .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), 
        .B1(\dp/ex_stage/muxA_out [9]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n176 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U182  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n46 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n6 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n45 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n176 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n130 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U181  ( .A1(\dp/ex_stage/alu/n34 ), 
        .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n21 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n175 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U180  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n51 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n6 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n50 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n175 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n127 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U179  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n130 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n127 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n174 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U178  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n134 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n170 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n128 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n133 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n44 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n103 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U177  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n17 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n103 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N215 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U176  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n21 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n8 ), .B1(\dp/ex_stage/alu/n37 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n173 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U175  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n20 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n51 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n173 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n123 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U174  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n170 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n32 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n133 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n151 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n172 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U173  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n150 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n123 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n31 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n96 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U172  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n16 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n96 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N216 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U171  ( .A1(\dp/ex_stage/alu/n37 ), 
        .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), .B1(
        \dp/ex_stage/muxA_out [15]), .B2(\dp/ex_stage/alu/shifter/sla_46/n11 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n171 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U170  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n22 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n20 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n171 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n118 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U169  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n170 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n146 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n133 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n147 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n169 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U168  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n145 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n118 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n38 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n84 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U167  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n16 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n84 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N217 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sla_46/U166  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n83 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U165  ( .A1(
        \dp/ex_stage/muxA_out [15]), .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), 
        .B1(\dp/ex_stage/muxA_out [16]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n168 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U164  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n23 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n22 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n168 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n111 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sla_46/U163  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n115 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sla_46/U162  ( .A1(\dp/ex_stage/alu/n29 ), 
        .A2(\dp/ex_stage/alu/shifter/sla_46/n18 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n167 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sla_46/U161  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n167 ), .A2(\dp/ex_stage/alu/n27 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n86 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U160  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n140 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n141 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n37 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n166 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U159  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n48 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n83 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n52 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n166 ), .ZN(
        \dp/ex_stage/alu/shifter/N218 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U158  ( .A1(
        \dp/ex_stage/muxA_out [16]), .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), 
        .B1(\dp/ex_stage/muxA_out [17]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n165 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U157  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n24 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n23 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n165 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n105 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U156  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n39 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n14 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n154 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n157 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sla_46/U155  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n134 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n157 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n159 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U154  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n127 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n130 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n128 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n164 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U153  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n53 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n159 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n164 ), .ZN(
        \dp/ex_stage/alu/shifter/N219 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U152  ( .A1(
        \dp/ex_stage/muxA_out [17]), .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), 
        .B1(\dp/ex_stage/muxA_out [18]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n163 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U151  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n25 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n24 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n163 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n98 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sla_46/U150  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n32 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n157 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n102 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U149  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n123 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n150 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n151 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n162 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U148  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n54 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n102 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n162 ), .ZN(
        \dp/ex_stage/alu/shifter/N220 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U147  ( .A1(
        \dp/ex_stage/muxA_out [18]), .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), 
        .B1(\dp/ex_stage/muxA_out [19]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n161 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U146  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n26 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n25 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n161 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n87 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sla_46/U145  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n146 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n157 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n82 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U144  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n118 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n145 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n147 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n160 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U143  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n55 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n82 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n160 ), .ZN(
        \dp/ex_stage/alu/shifter/N221 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U142  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n16 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n159 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N203 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U141  ( .A1(
        \dp/ex_stage/muxA_out [19]), .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), 
        .B1(\dp/ex_stage/muxA_out [20]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n158 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U140  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n58 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n26 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n158 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n113 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sla_46/U139  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n140 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n157 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n81 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U138  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n111 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n139 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n141 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n156 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U137  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n56 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n81 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n156 ), .ZN(
        \dp/ex_stage/alu/shifter/N222 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U136  ( .A1(
        \dp/ex_stage/muxA_out [20]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/muxA_out [21]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n155 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U135  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n60 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n58 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n155 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n107 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U134  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n134 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n128 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n36 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n80 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U133  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n105 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n127 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n130 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n153 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U132  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n80 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n153 ), .ZN(
        \dp/ex_stage/alu/shifter/N223 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U131  ( .A1(
        \dp/ex_stage/muxA_out [21]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/alu/n43 ), .B2(\dp/ex_stage/alu/shifter/sla_46/n10 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n152 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U130  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n62 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n60 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n152 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n100 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U129  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n32 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n151 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n36 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n79 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U128  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n98 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n123 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n150 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n149 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U127  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n59 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n79 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n149 ), .ZN(
        \dp/ex_stage/alu/shifter/N224 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U126  ( .A1(\dp/ex_stage/alu/n43 ), 
        .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), .B1(\dp/ex_stage/alu/n45 ), 
        .B2(\dp/ex_stage/alu/shifter/sla_46/n10 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n148 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U125  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n27 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n62 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n148 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n90 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U124  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n146 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n147 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n36 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n78 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U123  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n87 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n118 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n145 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n144 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U122  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n61 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n78 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n144 ), .ZN(
        \dp/ex_stage/alu/shifter/N225 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U121  ( .A1(\dp/ex_stage/alu/n45 ), 
        .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), .B1(
        \dp/ex_stage/muxA_out [24]), .B2(\dp/ex_stage/alu/shifter/sla_46/n10 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n143 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U120  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n28 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n27 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n143 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n142 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U119  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n140 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n141 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n36 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n77 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U118  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n113 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n111 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n139 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n138 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U117  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n63 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n77 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n138 ), .ZN(
        \dp/ex_stage/alu/shifter/N226 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U116  ( .A1(
        \dp/ex_stage/muxA_out [24]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/muxA_out [25]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n137 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U115  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n29 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n28 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n137 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n136 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sla_46/U114  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n133 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n134 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n135 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n132 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sla_46/U113  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n128 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n130 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n131 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n35 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n75 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U112  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n107 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n105 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n127 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n126 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U111  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n75 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n126 ), .ZN(
        \dp/ex_stage/alu/shifter/N227 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U110  ( .A1(
        \dp/ex_stage/muxA_out [25]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/muxA_out [26]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n125 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U109  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n67 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n29 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n125 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n124 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U108  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n100 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n98 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n123 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n122 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U107  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n65 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n121 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n122 ), .ZN(
        \dp/ex_stage/alu/shifter/N228 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U106  ( .A1(
        \dp/ex_stage/muxA_out [26]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/muxA_out [27]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n120 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U105  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n68 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n67 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n120 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n119 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U104  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n74 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n90 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n87 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n118 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n117 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U103  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n66 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n116 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n117 ), .ZN(
        \dp/ex_stage/alu/shifter/N229 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U102  ( .A1(
        \dp/ex_stage/muxA_out [27]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/muxA_out [28]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n114 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U101  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n69 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n68 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n114 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n112 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U100  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n111 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n73 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n113 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n110 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U99  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n63 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n83 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n109 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n110 ), .ZN(
        \dp/ex_stage/alu/shifter/N230 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U98  ( .A1(
        \dp/ex_stage/muxA_out [28]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/muxA_out [29]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n108 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U97  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n70 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n69 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n108 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n106 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U96  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n105 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n73 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n106 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n107 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n104 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U95  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n83 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n103 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n104 ), .ZN(
        \dp/ex_stage/alu/shifter/N231 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U94  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n16 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n102 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N204 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U93  ( .A1(
        \dp/ex_stage/muxA_out [29]), .A2(\dp/ex_stage/alu/shifter/sla_46/n7 ), 
        .B1(\dp/ex_stage/muxA_out [30]), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n10 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n101 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U92  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n1 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n71 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n4 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n70 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n101 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n99 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U91  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n98 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n73 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n99 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n97 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U90  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n65 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n83 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n96 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n97 ), .ZN(
        \dp/ex_stage/alu/shifter/N232 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sla_46/U89  ( .A1(
        \dp/ex_stage/muxA_out [30]), .A2(\dp/ex_stage/alu/shifter/sla_46/n8 ), 
        .B1(\dp/ex_stage/alu/shifter/N136 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n11 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n93 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U88  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n2 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n72 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n5 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n71 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n93 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n88 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sla_46/U87  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n86 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n87 ), .B1(
        \dp/ex_stage/alu/shifter/sla_46/n73 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n88 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n89 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n90 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n85 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sla_46/U86  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n66 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n83 ), .C1(
        \dp/ex_stage/alu/shifter/sla_46/n84 ), .C2(
        \dp/ex_stage/alu/shifter/sla_46/n18 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n85 ), .ZN(
        \dp/ex_stage/alu/shifter/N233 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U85  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n16 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n82 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N205 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U84  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n16 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n81 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N206 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U83  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n16 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n80 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N207 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U82  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n15 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n79 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N208 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U81  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n15 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n78 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N209 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U80  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n15 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n77 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N210 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sla_46/U79  ( .B1(
        \dp/ex_stage/alu/shifter/sla_46/n15 ), .B2(
        \dp/ex_stage/alu/shifter/sla_46/n75 ), .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N211 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U78  ( .A(\dp/ex_stage/alu/n45 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n29 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U77  ( .A(\dp/ex_stage/alu/n43 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n28 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U76  ( .A(\dp/ex_stage/muxA_out [21]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n27 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U75  ( .A(\dp/ex_stage/muxA_out [17]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n26 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U74  ( .A(\dp/ex_stage/muxA_out [16]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n25 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U73  ( .A(\dp/ex_stage/muxA_out [15]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n24 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U72  ( .A(\dp/ex_stage/alu/n37 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n23 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U71  ( .A(\dp/ex_stage/muxA_out [13]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n22 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U70  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n22 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n21 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U69  ( .A(\dp/ex_stage/alu/n34 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n20 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U68  ( .A(\dp/ex_stage/muxA_out [1]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n19 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U67  ( .A(\dp/ex_stage/alu/n27 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n14 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U66  ( .A(\dp/ex_stage/muxB_out [0]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n13 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U65  ( .A(\dp/ex_stage/muxA_out [5]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n43 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U64  ( .A(\dp/ex_stage/muxA_out [20]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n62 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U63  ( .A(\dp/ex_stage/muxA_out [19]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n60 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U62  ( .A(\dp/ex_stage/muxA_out [6]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n45 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U61  ( .A(\dp/ex_stage/muxA_out [4]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n42 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U60  ( .A(\dp/ex_stage/muxA_out [18]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n58 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U59  ( .A(
        \dp/ex_stage/alu/shifter/N202 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n39 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U58  ( .A(\dp/ex_stage/muxA_out [3]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n41 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U57  ( .A(\dp/ex_stage/muxA_out [24]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n67 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U56  ( .A(\dp/ex_stage/muxA_out [25]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n68 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U55  ( .A(\dp/ex_stage/muxA_out [26]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n69 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U54  ( .A(\dp/ex_stage/muxA_out [27]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n70 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U53  ( .A(\dp/ex_stage/muxA_out [28]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n71 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U52  ( .A(\dp/ex_stage/muxA_out [9]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n49 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U51  ( .A(\dp/ex_stage/muxA_out [2]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n40 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U50  ( .A(\dp/ex_stage/muxA_out [8]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n47 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U49  ( .A(\dp/ex_stage/muxA_out [7]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n46 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U48  ( .A(\dp/ex_stage/muxA_out [10]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n50 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U47  ( .A(\dp/ex_stage/muxA_out [11]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n51 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U46  ( .A(\dp/ex_stage/muxA_out [29]), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n72 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U45  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n142 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n63 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U44  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n136 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n64 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U43  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n124 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n65 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U42  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n119 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n66 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U41  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n187 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n32 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U40  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n113 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n56 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U39  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n107 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n57 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U38  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n139 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n48 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U37  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n54 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U36  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n87 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n55 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U35  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n92 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n6 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U34  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n95 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n12 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U33  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n154 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n36 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U32  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n92 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n5 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U31  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n92 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n4 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U30  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n95 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n11 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U29  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n95 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n10 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U28  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n172 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n31 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U27  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n169 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n38 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U26  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n37 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U25  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n174 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n44 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U24  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n132 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n35 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U23  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n186 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n30 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U22  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n182 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n33 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U21  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n178 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n34 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U20  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n90 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n61 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U19  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n59 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U18  ( .A(
        \dp/ex_stage/alu/shifter/n97 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n17 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U17  ( .A(
        \dp/ex_stage/alu/shifter/n97 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n15 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U16  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n91 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n3 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U15  ( .A(
        \dp/ex_stage/alu/shifter/n97 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n16 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U14  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n94 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n9 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U13  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n91 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n1 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U12  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n91 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n2 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U11  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n94 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n7 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sla_46/U10  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n94 ), .Z(
        \dp/ex_stage/alu/shifter/sla_46/n8 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sla_46/U9  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n167 ), .A2(
        \dp/ex_stage/alu/shifter/sla_46/n14 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n89 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U8  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n111 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n52 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U7  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n105 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n53 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U6  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n115 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n73 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U5  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n15 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n18 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sla_46/U4  ( .A(
        \dp/ex_stage/alu/shifter/sla_46/n83 ), .ZN(
        \dp/ex_stage/alu/shifter/sla_46/n74 ) );
  NOR2_X2 \dp/ex_stage/alu/shifter/sla_46/U3  ( .A1(\dp/ex_stage/alu/n27 ), 
        .A2(\dp/ex_stage/alu/n29 ), .ZN(\dp/ex_stage/alu/shifter/sla_46/n131 )
         );
  NOR2_X2 \dp/ex_stage/alu/shifter/sla_46/U2  ( .A1(
        \dp/ex_stage/alu/shifter/sla_46/n14 ), .A2(\dp/ex_stage/alu/n29 ), 
        .ZN(\dp/ex_stage/alu/shifter/sla_46/n129 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/srl_41/U200  ( .A1(\dp/ex_stage/alu/n25 ), 
        .A2(\dp/ex_stage/muxB_out [0]), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n96 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/srl_41/U199  ( .A1(\dp/ex_stage/alu/n25 ), 
        .A2(\dp/ex_stage/alu/shifter/srl_41/n2 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n97 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U198  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n19 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n18 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n167 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U197  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n56 ), .B2(\dp/ex_stage/muxA_out [7]), 
        .C1(\dp/ex_stage/alu/shifter/srl_41/n54 ), .C2(
        \dp/ex_stage/muxA_out [6]), .A(\dp/ex_stage/alu/shifter/srl_41/n167 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n88 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/srl_41/U196  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n91 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U195  ( .A1(\dp/ex_stage/alu/n45 ), 
        .A2(\dp/ex_stage/alu/shifter/srl_41/n56 ), .B1(\dp/ex_stage/alu/n43 ), 
        .B2(\dp/ex_stage/alu/shifter/srl_41/n54 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n166 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U194  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n14 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n40 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n166 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n74 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U193  ( .A1(
        \dp/ex_stage/muxA_out [17]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [16]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n165 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U192  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n38 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n36 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n165 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n73 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/srl_41/U191  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n3 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n4 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n142 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U190  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n3 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n4 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n129 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U189  ( .A1(
        \dp/ex_stage/muxA_out [29]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [28]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n164 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U188  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n52 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n51 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n164 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n111 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U187  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n4 ), .A2(\dp/ex_stage/alu/n27 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n117 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U186  ( .A1(
        \dp/ex_stage/muxA_out [25]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [24]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n163 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U185  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n48 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n46 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n163 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n115 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U184  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n129 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n111 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n117 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n115 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n162 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U183  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n74 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n73 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n42 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n131 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U182  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n4 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n7 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n159 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/srl_41/U181  ( .A1(\dp/ex_stage/alu/n27 ), 
        .A2(\dp/ex_stage/alu/shifter/srl_41/n159 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n67 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U180  ( .A1(
        \dp/ex_stage/muxA_out [13]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/alu/n34 ), .B2(\dp/ex_stage/alu/shifter/srl_41/n100 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n161 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U179  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n11 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n10 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n161 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n72 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/srl_41/U178  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n61 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U177  ( .A1(
        \dp/ex_stage/muxA_out [1]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/alu/shifter/N202 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n160 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U176  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n17 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n16 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n160 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n157 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U175  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n25 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n23 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n158 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U174  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n56 ), .B2(\dp/ex_stage/muxA_out [11]), 
        .C1(\dp/ex_stage/alu/shifter/srl_41/n54 ), .C2(
        \dp/ex_stage/muxA_out [10]), .A(\dp/ex_stage/alu/shifter/srl_41/n158 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n69 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U173  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n72 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n157 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n22 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n156 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U172  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n88 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n131 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n156 ), .ZN(
        \dp/ex_stage/alu/shifter/N137 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U171  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n29 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n27 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n155 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U170  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n56 ), .B2(\dp/ex_stage/muxA_out [13]), 
        .C1(\dp/ex_stage/alu/shifter/srl_41/n54 ), .C2(\dp/ex_stage/alu/n34 ), 
        .A(\dp/ex_stage/alu/shifter/srl_41/n155 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n107 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U169  ( .A1(
        \dp/ex_stage/muxA_out [27]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [26]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n154 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U168  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n50 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n49 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n154 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n119 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U167  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n51 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n52 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n103 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U166  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n119 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n103 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n112 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U165  ( .A1(
        \dp/ex_stage/muxA_out [15]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/alu/n37 ), .B2(\dp/ex_stage/alu/shifter/srl_41/n100 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n153 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U164  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n13 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n12 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n153 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n83 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U163  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n99 ), .A2(\dp/ex_stage/muxA_out [19]), 
        .B1(\dp/ex_stage/alu/shifter/srl_41/n100 ), .B2(
        \dp/ex_stage/muxA_out [18]), .ZN(\dp/ex_stage/alu/shifter/srl_41/n152 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U162  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n14 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n40 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n152 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n84 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U161  ( .A1(\dp/ex_stage/alu/n45 ), 
        .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), .B1(\dp/ex_stage/alu/n43 ), 
        .B2(\dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n151 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U160  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n44 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n41 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n151 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n120 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U159  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n57 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n83 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n84 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n120 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n150 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U158  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n107 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n112 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n150 ), .ZN(
        \dp/ex_stage/alu/shifter/N147 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U157  ( .A1(
        \dp/ex_stage/muxA_out [16]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [15]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n149 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U156  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n36 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n13 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n149 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n78 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U155  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n9 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n29 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n148 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U154  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n56 ), .B2(\dp/ex_stage/alu/n37 ), 
        .C1(\dp/ex_stage/alu/shifter/srl_41/n54 ), .C2(
        \dp/ex_stage/muxA_out [13]), .A(\dp/ex_stage/alu/shifter/srl_41/n148 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n95 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U153  ( .A1(
        \dp/ex_stage/muxA_out [24]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/alu/n45 ), .B2(\dp/ex_stage/alu/shifter/srl_41/n100 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n147 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U152  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n46 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n44 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n147 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n118 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U151  ( .A1(\dp/ex_stage/alu/n43 ), 
        .A2(\dp/ex_stage/alu/shifter/srl_41/n56 ), .B1(
        \dp/ex_stage/muxA_out [21]), .B2(\dp/ex_stage/alu/shifter/srl_41/n54 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n146 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U150  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n40 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n38 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n146 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n79 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U149  ( .A1(
        \dp/ex_stage/muxA_out [28]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [27]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n145 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U148  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n51 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n50 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n145 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n116 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U147  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n52 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n102 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/srl_41/U146  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n116 ), .B(
        \dp/ex_stage/alu/shifter/srl_41/n102 ), .S(\dp/ex_stage/alu/n27 ), .Z(
        \dp/ex_stage/alu/shifter/srl_41/n127 ) );
  NOR3_X1 \dp/ex_stage/alu/shifter/srl_41/U145  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A2(\dp/ex_stage/alu/n29 ), .A3(
        \dp/ex_stage/alu/shifter/srl_41/n47 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n144 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U144  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n118 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n79 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n144 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n143 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U143  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n33 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n95 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n143 ), .ZN(
        \dp/ex_stage/alu/shifter/N148 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U142  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n142 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n133 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U141  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n115 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n133 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n111 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n74 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n141 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U140  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n73 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n57 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n72 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n39 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n140 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U139  ( .A1(
        \dp/ex_stage/muxA_out [18]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [17]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n139 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U138  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n40 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n38 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n139 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n66 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U137  ( .A1(\dp/ex_stage/alu/n37 ), 
        .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), .B1(
        \dp/ex_stage/muxA_out [13]), .B2(\dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(\dp/ex_stage/alu/shifter/srl_41/n138 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U136  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n12 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n11 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n138 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n64 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U135  ( .A1(
        \dp/ex_stage/muxA_out [26]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [25]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n137 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U134  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n49 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n48 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n137 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n113 ) );
  OAI222_X1 \dp/ex_stage/alu/shifter/srl_41/U133  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n51 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n52 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n50 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n110 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U132  ( .A1(\dp/ex_stage/alu/n43 ), 
        .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), .B1(
        \dp/ex_stage/muxA_out [21]), .B2(\dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(\dp/ex_stage/alu/shifter/srl_41/n136 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U131  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n41 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n15 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n136 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n68 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U130  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n113 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n133 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n110 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n68 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n135 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U129  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n34 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n31 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n135 ), .ZN(
        \dp/ex_stage/alu/shifter/N150 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U128  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n119 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n133 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n103 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n120 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n134 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U127  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n35 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n32 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n134 ), .ZN(
        \dp/ex_stage/alu/shifter/N151 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U126  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n116 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n133 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n102 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n118 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n132 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U125  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n37 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n33 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n132 ), .ZN(
        \dp/ex_stage/alu/shifter/N152 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U124  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n6 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n131 ), .ZN(
        \dp/ex_stage/alu/shifter/N153 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U123  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n129 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n110 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n117 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n113 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n130 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U122  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n68 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n66 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n43 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n121 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U121  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n6 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n121 ), .ZN(
        \dp/ex_stage/alu/shifter/N154 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U120  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n129 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n103 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n117 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n119 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n128 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U119  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n120 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n84 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n45 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n104 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U118  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n6 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n104 ), .ZN(
        \dp/ex_stage/alu/shifter/N155 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U117  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n79 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n118 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n127 ), .C2(\dp/ex_stage/alu/n29 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n92 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U116  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n6 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n92 ), .ZN(
        \dp/ex_stage/alu/shifter/N156 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U115  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n20 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n19 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n126 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U114  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n56 ), .B2(\dp/ex_stage/muxA_out [8]), 
        .C1(\dp/ex_stage/alu/shifter/srl_41/n54 ), .C2(
        \dp/ex_stage/muxA_out [7]), .A(\dp/ex_stage/alu/shifter/srl_41/n126 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n85 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U113  ( .A1(
        \dp/ex_stage/muxA_out [2]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [1]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n125 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U112  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n18 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n17 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n125 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n123 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U111  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n27 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n25 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n124 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U110  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n56 ), .B2(\dp/ex_stage/alu/n34 ), 
        .C1(\dp/ex_stage/alu/shifter/srl_41/n54 ), .C2(
        \dp/ex_stage/muxA_out [11]), .A(\dp/ex_stage/alu/shifter/srl_41/n124 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n60 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U109  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n64 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n123 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n24 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n122 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U108  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n85 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n121 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n122 ), .ZN(
        \dp/ex_stage/alu/shifter/N138 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U107  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n115 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n111 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n117 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n74 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n89 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U106  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n6 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n89 ), .ZN(
        \dp/ex_stage/alu/shifter/N157 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U105  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n113 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n110 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n117 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n68 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n86 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U104  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n5 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n86 ), .ZN(
        \dp/ex_stage/alu/shifter/N158 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U103  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n119 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n103 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n117 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n120 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n81 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U102  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n5 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n81 ), .ZN(
        \dp/ex_stage/alu/shifter/N159 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U101  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n116 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n102 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n117 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n118 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n76 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U100  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n5 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/N160 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U99  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n115 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n111 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n70 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U98  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n5 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n70 ), .ZN(
        \dp/ex_stage/alu/shifter/N161 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U97  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n113 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n59 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n110 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n114 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n62 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U96  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n5 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n62 ), .ZN(
        \dp/ex_stage/alu/shifter/N162 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/srl_41/U95  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n5 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n112 ), .ZN(
        \dp/ex_stage/alu/shifter/N163 ) );
  NOR3_X1 \dp/ex_stage/alu/shifter/srl_41/U94  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n47 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n7 ), .A3(\dp/ex_stage/alu/n29 ), .ZN(
        \dp/ex_stage/alu/shifter/N164 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/srl_41/U93  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n111 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .ZN(
        \dp/ex_stage/alu/shifter/N165 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/srl_41/U92  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n110 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .ZN(
        \dp/ex_stage/alu/shifter/N166 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U91  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n21 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n20 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n109 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U90  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n56 ), .B2(\dp/ex_stage/muxA_out [9]), 
        .C1(\dp/ex_stage/alu/shifter/srl_41/n54 ), .C2(
        \dp/ex_stage/muxA_out [8]), .A(\dp/ex_stage/alu/shifter/srl_41/n109 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n80 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U89  ( .A1(
        \dp/ex_stage/muxA_out [3]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [2]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n108 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U88  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n19 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n18 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n108 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n106 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U87  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n83 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n106 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n26 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n105 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U86  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n80 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n104 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n105 ), .ZN(
        \dp/ex_stage/alu/shifter/N139 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/srl_41/U85  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n103 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .ZN(
        \dp/ex_stage/alu/shifter/N167 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/srl_41/U84  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n102 ), .ZN(
        \dp/ex_stage/alu/shifter/N168 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/srl_41/U83  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n23 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n55 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n21 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n101 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/srl_41/U82  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n56 ), .B2(\dp/ex_stage/muxA_out [10]), 
        .C1(\dp/ex_stage/alu/shifter/srl_41/n54 ), .C2(
        \dp/ex_stage/muxA_out [9]), .A(\dp/ex_stage/alu/shifter/srl_41/n101 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n75 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/srl_41/U81  ( .A1(
        \dp/ex_stage/muxA_out [4]), .A2(\dp/ex_stage/alu/shifter/srl_41/n99 ), 
        .B1(\dp/ex_stage/muxA_out [3]), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n98 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U80  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n20 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n1 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n19 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n94 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U79  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n78 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n58 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n94 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n28 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n93 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U78  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n75 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n92 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n93 ), .ZN(
        \dp/ex_stage/alu/shifter/N140 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U77  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n57 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n22 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n72 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n73 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n90 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U76  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n88 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n89 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n90 ), .ZN(
        \dp/ex_stage/alu/shifter/N141 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U75  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n57 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n24 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n64 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n66 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n87 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U74  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n85 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n86 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n87 ), .ZN(
        \dp/ex_stage/alu/shifter/N142 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U73  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n57 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n26 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n83 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n84 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n82 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U72  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n80 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n81 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n82 ), .ZN(
        \dp/ex_stage/alu/shifter/N143 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U71  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n57 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n28 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n78 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n79 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n77 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U70  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n75 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n76 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n77 ), .ZN(
        \dp/ex_stage/alu/shifter/N144 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U69  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n57 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n72 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n73 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n74 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n71 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U68  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n69 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n70 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n71 ), .ZN(
        \dp/ex_stage/alu/shifter/N145 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/srl_41/U67  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n57 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n64 ), .B1(
        \dp/ex_stage/alu/shifter/srl_41/n65 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n66 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n67 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n68 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n63 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/srl_41/U66  ( .B1(
        \dp/ex_stage/alu/shifter/srl_41/n60 ), .B2(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .C1(
        \dp/ex_stage/alu/shifter/srl_41/n62 ), .C2(
        \dp/ex_stage/alu/shifter/srl_41/n8 ), .A(
        \dp/ex_stage/alu/shifter/srl_41/n63 ), .ZN(
        \dp/ex_stage/alu/shifter/N146 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U65  ( .A(\dp/ex_stage/alu/n45 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n15 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U64  ( .A(\dp/ex_stage/muxA_out [21]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n14 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U63  ( .A(\dp/ex_stage/muxA_out [17]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n13 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U62  ( .A(\dp/ex_stage/muxA_out [16]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n12 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U61  ( .A(\dp/ex_stage/muxA_out [15]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n11 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U60  ( .A(\dp/ex_stage/alu/n37 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n10 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U59  ( .A(\dp/ex_stage/alu/n34 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n9 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U58  ( .A(\dp/ex_stage/alu/n29 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n4 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U57  ( .A(\dp/ex_stage/alu/n27 ), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n3 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U56  ( .A(\dp/ex_stage/muxB_out [0]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n2 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U55  ( .A(\dp/ex_stage/muxA_out [18]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n36 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U54  ( .A(\dp/ex_stage/muxA_out [24]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n41 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U53  ( .A(\dp/ex_stage/muxA_out [25]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n44 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U52  ( .A(\dp/ex_stage/muxA_out [28]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n49 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U51  ( .A(\dp/ex_stage/muxA_out [26]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n46 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U50  ( .A(\dp/ex_stage/muxA_out [27]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n48 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U49  ( .A(\dp/ex_stage/muxA_out [3]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n17 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U48  ( .A(\dp/ex_stage/muxA_out [9]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n25 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U47  ( .A(\dp/ex_stage/muxA_out [7]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n21 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U46  ( .A(\dp/ex_stage/muxA_out [8]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n23 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U45  ( .A(\dp/ex_stage/muxA_out [10]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n27 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U44  ( .A(\dp/ex_stage/muxA_out [11]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n29 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U43  ( .A(\dp/ex_stage/muxA_out [19]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n38 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U42  ( .A(\dp/ex_stage/muxA_out [29]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n50 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U41  ( .A(\dp/ex_stage/muxA_out [4]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n18 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U40  ( .A(\dp/ex_stage/muxA_out [6]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n20 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U39  ( .A(\dp/ex_stage/muxA_out [5]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n19 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U38  ( .A(\dp/ex_stage/muxA_out [20]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n40 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U37  ( .A(
        \dp/ex_stage/alu/shifter/N136 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n52 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U36  ( .A(\dp/ex_stage/muxA_out [30]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n51 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U35  ( .A(\dp/ex_stage/muxA_out [2]), 
        .ZN(\dp/ex_stage/alu/shifter/srl_41/n16 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U34  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n66 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n34 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U33  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n84 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n35 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U32  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n69 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n22 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U31  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n60 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n24 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U30  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n130 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n43 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U29  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n162 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n42 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U28  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n96 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n56 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U27  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n140 ), .ZN(
        \dp/ex_stage/alu/shifter/N149 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U26  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n128 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n45 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U25  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n141 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n39 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U24  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n53 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U23  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n127 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n47 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/srl_41/U22  ( .A(
        \dp/ex_stage/alu/shifter/n99 ), .Z(\dp/ex_stage/alu/shifter/srl_41/n7 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U21  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n79 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n37 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/srl_41/U20  ( .A(
        \dp/ex_stage/alu/shifter/n99 ), .Z(\dp/ex_stage/alu/shifter/srl_41/n6 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/srl_41/U19  ( .A(
        \dp/ex_stage/alu/shifter/n99 ), .Z(\dp/ex_stage/alu/shifter/srl_41/n5 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U18  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n64 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n31 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U17  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n83 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n32 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U16  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n95 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n28 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U15  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n107 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n26 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U14  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n78 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n33 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/srl_41/U13  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n97 ), .Z(
        \dp/ex_stage/alu/shifter/srl_41/n1 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/srl_41/U12  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n159 ), .A2(
        \dp/ex_stage/alu/shifter/srl_41/n3 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n65 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U11  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n97 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n54 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U10  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n99 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n55 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U9  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n7 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n8 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U8  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n91 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n57 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U7  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n142 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n59 ) );
  INV_X1 \dp/ex_stage/alu/shifter/srl_41/U6  ( .A(
        \dp/ex_stage/alu/shifter/srl_41/n61 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n58 ) );
  NOR2_X2 \dp/ex_stage/alu/shifter/srl_41/U5  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n2 ), .A2(\dp/ex_stage/alu/n25 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n99 ) );
  NOR2_X2 \dp/ex_stage/alu/shifter/srl_41/U4  ( .A1(
        \dp/ex_stage/alu/shifter/srl_41/n3 ), .A2(\dp/ex_stage/alu/n29 ), .ZN(
        \dp/ex_stage/alu/shifter/srl_41/n114 ) );
  NOR2_X2 \dp/ex_stage/alu/shifter/srl_41/U3  ( .A1(\dp/ex_stage/muxB_out [0]), 
        .A2(\dp/ex_stage/alu/n25 ), .ZN(\dp/ex_stage/alu/shifter/srl_41/n100 )
         );
  NAND2_X1 \dp/ex_stage/alu/shifter/sra_39/U206  ( .A1(
        \dp/ex_stage/muxB_out [0]), .A2(\dp/ex_stage/alu/shifter/sra_39/n2 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n97 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/sra_39/U205  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n15 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n14 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n174 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U204  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [6]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [7]), .A(\dp/ex_stage/alu/shifter/sra_39/n174 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n85 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sra_39/U203  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n88 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U202  ( .A1(\dp/ex_stage/alu/n43 ), 
        .A2(\dp/ex_stage/alu/shifter/sra_39/n94 ), .B1(\dp/ex_stage/alu/n45 ), 
        .B2(\dp/ex_stage/alu/shifter/sra_39/n95 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n173 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U201  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n10 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n37 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n173 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n72 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U200  ( .A1(
        \dp/ex_stage/muxA_out [17]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [16]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n172 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U199  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n34 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n36 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n172 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n71 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sra_39/U198  ( .A1(\dp/ex_stage/alu/n27 ), 
        .A2(\dp/ex_stage/alu/n29 ), .ZN(\dp/ex_stage/alu/shifter/sra_39/n136 )
         );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U197  ( .A1(
        \dp/ex_stage/muxA_out [29]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [28]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n171 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U196  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n50 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n51 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n171 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n115 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sra_39/U195  ( .A1(\dp/ex_stage/alu/n29 ), 
        .A2(\dp/ex_stage/alu/shifter/sra_39/n3 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n122 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U194  ( .A1(
        \dp/ex_stage/muxA_out [25]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [24]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n170 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U193  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n42 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n44 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n170 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n116 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U192  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n136 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n115 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n122 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n116 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n169 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U191  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n72 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n71 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n39 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n139 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sra_39/U190  ( .A1(\dp/ex_stage/alu/n29 ), 
        .A2(\dp/ex_stage/alu/shifter/sra_39/n7 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n166 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sra_39/U189  ( .A1(\dp/ex_stage/alu/n27 ), 
        .A2(\dp/ex_stage/alu/shifter/sra_39/n166 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n66 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U188  ( .A1(
        \dp/ex_stage/muxA_out [13]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/alu/n34 ), .B2(\dp/ex_stage/alu/shifter/sra_39/n56 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n168 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U187  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/alu/n37 ), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [15]), .A(\dp/ex_stage/alu/shifter/sra_39/n27 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n149 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sra_39/U186  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n61 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U185  ( .A1(
        \dp/ex_stage/muxA_out [1]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/alu/shifter/N202 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n167 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U184  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n12 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n13 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n167 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n164 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/sra_39/U183  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n21 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n19 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n165 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U182  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [10]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [11]), .A(\dp/ex_stage/alu/shifter/sra_39/n165 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n68 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U181  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n26 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n58 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n164 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n18 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n163 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U180  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n85 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n88 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n139 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n163 ), .ZN(
        \dp/ex_stage/alu/shifter/N105 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/sra_39/U179  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n25 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n23 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n162 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U178  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/alu/n34 ), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [13]), .A(\dp/ex_stage/alu/shifter/sra_39/n162 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n104 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/sra_39/U177  ( .A(
        \dp/ex_stage/muxA_out [30]), .B(\dp/ex_stage/alu/shifter/N136 ), .S(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .Z(
        \dp/ex_stage/alu/shifter/sra_39/n123 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U176  ( .A1(
        \dp/ex_stage/muxA_out [27]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [26]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n161 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U175  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n45 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n48 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n161 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n119 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sra_39/U174  ( .A1(
        \dp/ex_stage/alu/shifter/N136 ), .A2(\dp/ex_stage/alu/n29 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n135 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U173  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n123 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n119 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n52 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n110 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U172  ( .A1(
        \dp/ex_stage/muxA_out [15]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/alu/n37 ), .B2(\dp/ex_stage/alu/shifter/sra_39/n56 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n160 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U171  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [16]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [17]), .A(\dp/ex_stage/alu/shifter/sra_39/n31 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n141 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U170  ( .A1(
        \dp/ex_stage/muxA_out [20]), .A2(\dp/ex_stage/alu/shifter/sra_39/n94 ), 
        .B1(\dp/ex_stage/muxA_out [21]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n95 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n159 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U169  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n36 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n34 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n159 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n81 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U168  ( .A1(\dp/ex_stage/alu/n45 ), 
        .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), .B1(\dp/ex_stage/alu/n43 ), 
        .B2(\dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n158 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U167  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n38 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n41 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n158 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n120 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U166  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n30 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n81 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n120 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n157 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U165  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n104 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n110 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n157 ), .ZN(
        \dp/ex_stage/alu/shifter/N115 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/sra_39/U164  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n8 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n25 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n156 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U163  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [13]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(\dp/ex_stage/alu/n37 ), 
        .A(\dp/ex_stage/alu/shifter/sra_39/n156 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n92 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U162  ( .A1(
        \dp/ex_stage/muxA_out [28]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [27]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n155 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U161  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n48 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n50 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n155 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n117 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U160  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n3 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n51 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n135 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n143 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sra_39/U159  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n117 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n143 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n109 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U158  ( .A1(
        \dp/ex_stage/muxA_out [16]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [15]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n154 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U157  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n9 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n34 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n154 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n76 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U156  ( .A1(
        \dp/ex_stage/muxA_out [21]), .A2(\dp/ex_stage/alu/shifter/sra_39/n94 ), 
        .B1(\dp/ex_stage/alu/n43 ), .B2(\dp/ex_stage/alu/shifter/sra_39/n95 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n153 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U155  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n37 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n36 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n153 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n77 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U154  ( .A1(
        \dp/ex_stage/muxA_out [24]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/alu/n45 ), .B2(\dp/ex_stage/alu/shifter/sra_39/n56 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n152 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U153  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n41 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n42 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n152 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n118 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U152  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n76 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n77 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n118 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n151 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U151  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n92 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n109 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n151 ), .ZN(
        \dp/ex_stage/alu/shifter/N116 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sra_39/U150  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n115 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n143 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n108 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U149  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n71 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n72 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n116 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n150 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U148  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n149 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n108 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n150 ), .ZN(
        \dp/ex_stage/alu/shifter/N117 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U147  ( .A1(\dp/ex_stage/alu/n37 ), 
        .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), .B1(
        \dp/ex_stage/muxA_out [13]), .B2(\dp/ex_stage/alu/shifter/sra_39/n56 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n148 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U146  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [15]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [16]), .A(\dp/ex_stage/alu/shifter/sra_39/n29 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n132 ) );
  OAI222_X1 \dp/ex_stage/alu/shifter/sra_39/U145  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n48 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n50 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n2 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n51 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n111 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sra_39/U144  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n111 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n143 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n107 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U143  ( .A1(
        \dp/ex_stage/muxA_out [18]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [17]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n147 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U142  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n36 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n37 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n147 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n65 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U141  ( .A1(\dp/ex_stage/alu/n43 ), 
        .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), .B1(
        \dp/ex_stage/muxA_out [21]), .B2(\dp/ex_stage/alu/shifter/sra_39/n56 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n146 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U140  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n11 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n38 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n146 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n67 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U139  ( .A1(
        \dp/ex_stage/muxA_out [26]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [25]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n145 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U138  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n44 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n45 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n145 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n113 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U137  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n65 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n67 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n113 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n144 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U136  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n132 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n107 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n144 ), .ZN(
        \dp/ex_stage/alu/shifter/N118 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sra_39/U135  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n123 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n143 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n99 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U134  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n81 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n120 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n119 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n142 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U133  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n141 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n99 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n142 ), .ZN(
        \dp/ex_stage/alu/shifter/N119 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sra_39/U132  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n6 ), .A2(
        \dp/ex_stage/alu/shifter/N136 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n100 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U131  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n117 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n118 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n53 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n140 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U130  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n35 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n88 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n32 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n140 ), .ZN(
        \dp/ex_stage/alu/shifter/N120 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U129  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n6 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n139 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N121 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U128  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n136 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n111 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n122 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n113 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n138 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U127  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n67 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n65 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n40 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n127 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U126  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n6 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n127 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N122 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U125  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n120 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n81 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n137 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U124  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n123 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n136 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n119 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n122 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n33 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n101 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U123  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n6 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n101 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N123 ) );
  NOR2_X1 \dp/ex_stage/alu/shifter/sra_39/U122  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n135 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n3 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n124 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sra_39/U121  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n122 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n117 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n124 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n134 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U120  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n118 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n77 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n43 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n89 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U119  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n6 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n89 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N124 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/sra_39/U118  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n16 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n15 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n133 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U117  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [7]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [8]), .A(\dp/ex_stage/alu/shifter/sra_39/n133 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n82 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U116  ( .A1(
        \dp/ex_stage/muxA_out [2]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [1]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n131 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U115  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n13 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n14 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n131 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n129 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/sra_39/U114  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n23 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n21 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n130 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U113  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [11]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(\dp/ex_stage/alu/n34 ), 
        .A(\dp/ex_stage/alu/shifter/sra_39/n130 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n60 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U112  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n28 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n58 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n129 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n20 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n128 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U111  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n82 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n88 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n127 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n128 ), .ZN(
        \dp/ex_stage/alu/shifter/N106 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sra_39/U110  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n122 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n115 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n124 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n126 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U109  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n116 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n72 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n46 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n86 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U108  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n5 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n86 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N125 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sra_39/U107  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n122 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n111 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n124 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n125 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U106  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n113 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n67 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n47 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n83 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U105  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n5 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n83 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N126 ) );
  AOI21_X1 \dp/ex_stage/alu/shifter/sra_39/U104  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n122 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n123 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n124 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n121 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U103  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n119 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n120 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n49 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n79 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U102  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n5 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n79 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N127 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U101  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n117 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n118 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n52 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n74 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U100  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n5 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n74 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N128 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U99  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n115 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n116 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n52 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n69 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U98  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n5 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n69 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N129 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U97  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n111 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n112 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n113 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n114 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n52 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n62 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U96  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n5 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n62 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N130 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U95  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n5 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n110 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N131 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U94  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n4 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n109 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N132 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U93  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n4 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n108 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N133 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U92  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n4 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n107 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N134 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/sra_39/U91  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n17 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n16 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n106 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U90  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [8]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [9]), .A(\dp/ex_stage/alu/shifter/sra_39/n106 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n78 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U89  ( .A1(
        \dp/ex_stage/muxA_out [3]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [2]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n105 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U88  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n14 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n15 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n105 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n103 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U87  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n30 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n58 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n103 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n22 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n102 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U86  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n78 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n88 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n101 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n102 ), .ZN(
        \dp/ex_stage/alu/shifter/N107 ) );
  OAI21_X1 \dp/ex_stage/alu/shifter/sra_39/U85  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n4 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n99 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/N135 ) );
  OAI22_X1 \dp/ex_stage/alu/shifter/sra_39/U84  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n19 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n17 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n96 ) );
  AOI221_X1 \dp/ex_stage/alu/shifter/sra_39/U83  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .B2(\dp/ex_stage/muxA_out [9]), 
        .C1(\dp/ex_stage/alu/shifter/sra_39/n95 ), .C2(
        \dp/ex_stage/muxA_out [10]), .A(\dp/ex_stage/alu/shifter/sra_39/n96 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n73 ) );
  AOI22_X1 \dp/ex_stage/alu/shifter/sra_39/U82  ( .A1(
        \dp/ex_stage/muxA_out [4]), .A2(\dp/ex_stage/alu/shifter/sra_39/n54 ), 
        .B1(\dp/ex_stage/muxA_out [3]), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n56 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n93 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U81  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n57 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n15 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n55 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n16 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n93 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n91 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U80  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n76 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n58 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n91 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n24 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n90 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U79  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n73 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n88 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n89 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n90 ), .ZN(
        \dp/ex_stage/alu/shifter/N108 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U78  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n18 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n26 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n71 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n87 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U77  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n85 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n86 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n87 ), .ZN(
        \dp/ex_stage/alu/shifter/N109 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U76  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n20 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n28 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n65 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n84 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U75  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n82 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n83 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n84 ), .ZN(
        \dp/ex_stage/alu/shifter/N110 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U74  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n22 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n30 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n81 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n80 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U73  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n78 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n79 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n80 ), .ZN(
        \dp/ex_stage/alu/shifter/N111 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U72  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n24 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n76 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n77 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n75 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U71  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n73 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n74 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n75 ), .ZN(
        \dp/ex_stage/alu/shifter/N112 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U70  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n26 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n71 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n72 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n70 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U69  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n68 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n69 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n70 ), .ZN(
        \dp/ex_stage/alu/shifter/N113 ) );
  AOI222_X1 \dp/ex_stage/alu/shifter/sra_39/U68  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n59 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n28 ), .B1(
        \dp/ex_stage/alu/shifter/sra_39/n64 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n65 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n66 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n67 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n63 ) );
  OAI221_X1 \dp/ex_stage/alu/shifter/sra_39/U67  ( .B1(
        \dp/ex_stage/alu/shifter/sra_39/n60 ), .B2(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .C1(
        \dp/ex_stage/alu/shifter/sra_39/n62 ), .C2(
        \dp/ex_stage/alu/shifter/sra_39/n7 ), .A(
        \dp/ex_stage/alu/shifter/sra_39/n63 ), .ZN(
        \dp/ex_stage/alu/shifter/N114 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U66  ( .A(\dp/ex_stage/alu/n45 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n11 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U65  ( .A(\dp/ex_stage/muxA_out [21]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n10 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U64  ( .A(\dp/ex_stage/muxA_out [17]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n9 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U63  ( .A(\dp/ex_stage/alu/n34 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n8 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U62  ( .A(\dp/ex_stage/alu/n27 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n3 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U61  ( .A(\dp/ex_stage/alu/n25 ), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n2 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U60  ( .A(\dp/ex_stage/muxB_out [0]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n1 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U59  ( .A(\dp/ex_stage/muxA_out [24]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n38 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U58  ( .A(\dp/ex_stage/muxA_out [28]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n45 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U57  ( .A(\dp/ex_stage/muxA_out [25]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n41 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U56  ( .A(\dp/ex_stage/muxA_out [27]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n44 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U55  ( .A(\dp/ex_stage/muxA_out [26]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n42 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U54  ( .A(\dp/ex_stage/muxA_out [3]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n13 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U53  ( .A(
        \dp/ex_stage/alu/shifter/N136 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n51 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U52  ( .A(\dp/ex_stage/muxA_out [9]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n21 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U51  ( .A(\dp/ex_stage/muxA_out [7]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n17 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U50  ( .A(\dp/ex_stage/muxA_out [8]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n19 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U49  ( .A(\dp/ex_stage/muxA_out [10]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n23 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U48  ( .A(\dp/ex_stage/muxA_out [11]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n25 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U47  ( .A(\dp/ex_stage/muxA_out [20]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n37 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U46  ( .A(\dp/ex_stage/muxA_out [30]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n50 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U45  ( .A(\dp/ex_stage/muxA_out [29]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n48 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U44  ( .A(\dp/ex_stage/muxA_out [4]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n14 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U43  ( .A(\dp/ex_stage/muxA_out [6]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n16 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U42  ( .A(\dp/ex_stage/muxA_out [18]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n34 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U41  ( .A(\dp/ex_stage/muxA_out [5]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n15 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U40  ( .A(\dp/ex_stage/muxA_out [19]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n36 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U39  ( .A(\dp/ex_stage/muxA_out [2]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n12 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U38  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n135 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n52 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U37  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n68 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n18 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U36  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n60 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n20 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U35  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n134 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n43 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U34  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n126 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n46 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U33  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n100 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n53 ) );
  NAND2_X1 \dp/ex_stage/alu/shifter/sra_39/U32  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n1 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n2 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n98 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U31  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n137 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n33 ) );
  NOR2_X2 \dp/ex_stage/alu/shifter/sra_39/U30  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n1 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n2 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n95 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U29  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n94 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n57 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U28  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n97 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n54 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U27  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n169 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n39 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U26  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n138 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n40 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U25  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n125 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n47 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U24  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n121 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n49 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U23  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n168 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n27 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U22  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n148 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n29 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U21  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n160 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n31 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sra_39/U20  ( .A(
        \dp/ex_stage/alu/shifter/n98 ), .Z(\dp/ex_stage/alu/shifter/sra_39/n6 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U19  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n77 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n35 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U18  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n76 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n32 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sra_39/U17  ( .A(
        \dp/ex_stage/alu/shifter/n98 ), .Z(\dp/ex_stage/alu/shifter/sra_39/n4 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/sra_39/U16  ( .A(
        \dp/ex_stage/alu/shifter/n98 ), .Z(\dp/ex_stage/alu/shifter/sra_39/n5 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U15  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n104 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n22 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U14  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n92 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n24 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U13  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n149 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n26 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U12  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n132 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n28 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U11  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n141 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n30 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U10  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n95 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n55 ) );
  AND2_X1 \dp/ex_stage/alu/shifter/sra_39/U9  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n166 ), .A2(
        \dp/ex_stage/alu/shifter/sra_39/n3 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n64 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U8  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n98 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n56 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U7  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n61 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n58 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U6  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n4 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n7 ) );
  INV_X1 \dp/ex_stage/alu/shifter/sra_39/U5  ( .A(
        \dp/ex_stage/alu/shifter/sra_39/n88 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n59 ) );
  NOR2_X2 \dp/ex_stage/alu/shifter/sra_39/U4  ( .A1(\dp/ex_stage/alu/n27 ), 
        .A2(\dp/ex_stage/alu/n29 ), .ZN(\dp/ex_stage/alu/shifter/sra_39/n114 )
         );
  NOR2_X2 \dp/ex_stage/alu/shifter/sra_39/U3  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n2 ), .A2(\dp/ex_stage/muxB_out [0]), 
        .ZN(\dp/ex_stage/alu/shifter/sra_39/n94 ) );
  NOR2_X2 \dp/ex_stage/alu/shifter/sra_39/U2  ( .A1(
        \dp/ex_stage/alu/shifter/sra_39/n3 ), .A2(\dp/ex_stage/alu/n29 ), .ZN(
        \dp/ex_stage/alu/shifter/sra_39/n112 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U16  ( .A(\dp/ex_stage/muxB_out [0]), 
        .Z(\dp/ex_stage/alu/shifter/rol_32/n3 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U15  ( .A(\dp/ex_stage/muxB_out [0]), 
        .Z(\dp/ex_stage/alu/shifter/rol_32/n2 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U14  ( .A(\dp/ex_stage/muxB_out [0]), 
        .Z(\dp/ex_stage/alu/shifter/rol_32/n1 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U13  ( .A(\dp/ex_stage/alu/n27 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n9 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U12  ( .A(\dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n12 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U11  ( .A(\dp/ex_stage/alu/n25 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n6 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U10  ( .A(\dp/ex_stage/alu/n27 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n7 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U9  ( .A(\dp/ex_stage/alu/n27 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n8 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U8  ( .A(\dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n10 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U7  ( .A(\dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n11 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U6  ( .A(\dp/ex_stage/alu/n25 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n5 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U5  ( .A(\dp/ex_stage/alu/n25 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n4 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U4  ( .A(
        \dp/ex_stage/alu/shifter/n98 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n15 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U3  ( .A(
        \dp/ex_stage/alu/shifter/n98 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n13 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/rol_32/U2  ( .A(
        \dp/ex_stage/alu/shifter/n98 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/n14 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_0_0  ( .A(
        \dp/ex_stage/alu/shifter/N202 ), .B(\dp/ex_stage/alu/shifter/N136 ), 
        .S(\dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][0] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_1  ( .A(
        \dp/ex_stage/muxA_out [1]), .B(\dp/ex_stage/alu/shifter/N202 ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_2  ( .A(
        \dp/ex_stage/muxA_out [2]), .B(\dp/ex_stage/muxA_out [1]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_3  ( .A(
        \dp/ex_stage/muxA_out [3]), .B(\dp/ex_stage/muxA_out [2]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_4  ( .A(
        \dp/ex_stage/muxA_out [4]), .B(\dp/ex_stage/muxA_out [3]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_5  ( .A(
        \dp/ex_stage/muxA_out [5]), .B(\dp/ex_stage/muxA_out [4]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_6  ( .A(
        \dp/ex_stage/muxA_out [6]), .B(\dp/ex_stage/muxA_out [5]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_7  ( .A(
        \dp/ex_stage/muxA_out [7]), .B(\dp/ex_stage/muxA_out [6]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_8  ( .A(
        \dp/ex_stage/muxA_out [8]), .B(\dp/ex_stage/muxA_out [7]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_9  ( .A(
        \dp/ex_stage/muxA_out [9]), .B(\dp/ex_stage/muxA_out [8]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_10  ( .A(
        \dp/ex_stage/muxA_out [10]), .B(\dp/ex_stage/muxA_out [9]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n1 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_11  ( .A(
        \dp/ex_stage/muxA_out [11]), .B(\dp/ex_stage/muxA_out [10]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_12  ( .A(\dp/ex_stage/alu/n34 ), 
        .B(\dp/ex_stage/muxA_out [11]), .S(\dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(\dp/ex_stage/alu/shifter/rol_32/ML_int[1][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_13  ( .A(
        \dp/ex_stage/muxA_out [13]), .B(\dp/ex_stage/alu/n34 ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_14  ( .A(\dp/ex_stage/alu/n37 ), 
        .B(\dp/ex_stage/muxA_out [13]), .S(\dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(\dp/ex_stage/alu/shifter/rol_32/ML_int[1][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_15  ( .A(
        \dp/ex_stage/muxA_out [15]), .B(\dp/ex_stage/alu/n37 ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_16  ( .A(
        \dp/ex_stage/muxA_out [16]), .B(\dp/ex_stage/muxA_out [15]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_17  ( .A(
        \dp/ex_stage/muxA_out [17]), .B(\dp/ex_stage/muxA_out [16]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_18  ( .A(
        \dp/ex_stage/muxA_out [18]), .B(\dp/ex_stage/muxA_out [17]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_19  ( .A(
        \dp/ex_stage/muxA_out [19]), .B(\dp/ex_stage/muxA_out [18]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_20  ( .A(
        \dp/ex_stage/muxA_out [20]), .B(\dp/ex_stage/muxA_out [19]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_21  ( .A(
        \dp/ex_stage/muxA_out [21]), .B(\dp/ex_stage/muxA_out [20]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n2 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_22  ( .A(\dp/ex_stage/alu/n43 ), 
        .B(\dp/ex_stage/muxA_out [21]), .S(\dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(\dp/ex_stage/alu/shifter/rol_32/ML_int[1][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_23  ( .A(\dp/ex_stage/alu/n45 ), 
        .B(\dp/ex_stage/alu/n43 ), .S(\dp/ex_stage/alu/shifter/rol_32/n3 ), 
        .Z(\dp/ex_stage/alu/shifter/rol_32/ML_int[1][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_24  ( .A(
        \dp/ex_stage/muxA_out [24]), .B(\dp/ex_stage/alu/n45 ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_25  ( .A(
        \dp/ex_stage/muxA_out [25]), .B(\dp/ex_stage/muxA_out [24]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_26  ( .A(
        \dp/ex_stage/muxA_out [26]), .B(\dp/ex_stage/muxA_out [25]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_27  ( .A(
        \dp/ex_stage/muxA_out [27]), .B(\dp/ex_stage/muxA_out [26]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_28  ( .A(
        \dp/ex_stage/muxA_out [28]), .B(\dp/ex_stage/muxA_out [27]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_29  ( .A(
        \dp/ex_stage/muxA_out [29]), .B(\dp/ex_stage/muxA_out [28]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_30  ( .A(
        \dp/ex_stage/muxA_out [30]), .B(\dp/ex_stage/muxA_out [29]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_0_31  ( .A(
        \dp/ex_stage/alu/shifter/N136 ), .B(\dp/ex_stage/muxA_out [30]), .S(
        \dp/ex_stage/alu/shifter/rol_32/n3 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_1_0  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][0] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][30] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][0] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_1_1  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][1] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][31] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_2  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][2] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][0] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_3  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][3] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][1] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_4  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][4] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][2] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_5  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][5] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][3] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_6  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][6] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][4] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_7  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][7] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][5] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_8  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][8] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][6] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_9  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][9] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][7] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_10  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][10] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][8] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n4 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_11  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][11] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][9] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_12  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][12] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][10] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_13  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][13] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][11] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_14  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][14] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][12] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_15  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][15] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][13] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_16  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][16] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][14] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_17  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][17] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][15] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_18  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][18] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][16] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_19  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][19] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][17] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_20  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][20] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][18] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_21  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][21] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][19] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n5 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_22  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][22] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][20] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_23  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][23] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][21] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_24  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][24] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][22] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_25  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][25] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][23] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_26  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][26] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][24] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_27  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][27] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][25] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_28  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][28] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][26] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_29  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][29] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][27] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_30  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][30] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][28] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_1_31  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][31] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[1][29] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n6 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_2_0  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][0] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][28] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][0] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_2_1  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][1] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][29] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_2_2  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][2] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][30] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_2_3  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][3] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][31] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_4  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][4] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][0] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_5  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][5] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][1] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_6  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][6] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][2] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_7  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][7] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][3] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_8  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][8] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][4] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_9  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][9] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][5] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_10  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][10] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][6] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n7 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_11  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][11] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][7] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_12  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][12] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][8] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_13  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][13] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][9] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_14  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][14] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][10] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_15  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][15] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][11] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_16  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][16] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][12] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_17  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][17] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][13] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_18  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][18] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][14] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_19  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][19] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][15] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_20  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][20] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][16] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_21  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][21] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][17] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n8 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_22  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][22] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][18] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_23  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][23] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][19] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_24  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][24] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][20] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_25  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][25] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][21] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_26  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][26] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][22] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_27  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][27] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][23] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_28  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][28] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][24] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_29  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][29] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][25] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_30  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][30] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][26] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_2_31  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][31] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[2][27] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n9 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_3_0  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][0] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][24] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][0] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_3_1  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][1] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][25] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_3_2  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][2] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][26] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_3_3  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][3] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][27] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_3_4  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][4] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][28] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_3_5  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][5] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][29] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_3_6  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][6] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][30] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_3_7  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][7] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][31] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_8  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][8] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][0] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_9  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][9] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][1] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_10  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][10] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][2] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n10 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_11  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][11] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][3] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_12  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][12] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][4] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_13  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][13] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][5] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_14  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][14] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][6] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_15  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][15] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][7] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_16  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][16] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][8] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_17  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][17] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][9] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_18  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][18] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][10] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_19  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][19] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][11] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_20  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][20] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][12] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_21  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][21] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][13] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n11 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_22  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][22] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][14] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_23  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][23] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][15] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_24  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][24] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][16] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_25  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][25] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][17] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_26  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][26] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][18] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_27  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][27] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][19] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_28  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][28] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][20] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_29  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][29] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][21] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_30  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][30] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][22] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_3_31  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][31] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[3][23] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n12 ), .Z(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_0  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][0] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][16] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N39 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_1  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][1] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][17] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N40 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_2  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][2] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][18] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N41 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_3  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][3] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][19] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N42 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_4  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][4] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][20] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N43 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_5  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][5] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][21] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N44 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_6  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][6] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][22] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N45 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_7  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][7] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][23] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N46 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_8  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][8] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][24] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N47 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_9  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][9] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][25] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N48 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_10  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][10] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][26] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N49 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_11  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][11] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][27] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N50 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_12  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][12] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][28] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N51 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_13  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][13] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][29] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N52 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_14  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][14] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][30] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N53 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M0_4_15  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][15] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][31] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N54 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_16  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][16] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][0] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N55 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_17  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][17] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][1] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N56 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_18  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][18] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][2] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N57 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_19  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][19] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][3] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N58 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_20  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][20] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][4] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N59 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_21  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][21] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][5] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N60 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_22  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][22] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][6] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N61 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_23  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][23] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][7] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N62 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_24  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][24] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][8] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N63 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_25  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][25] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][9] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N64 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_26  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][26] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][10] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N65 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_27  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][27] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][11] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N66 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_28  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][28] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][12] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N67 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_29  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][29] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][13] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N68 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_30  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][30] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][14] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N69 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/rol_32/M1_4_31  ( .A(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][31] ), .B(
        \dp/ex_stage/alu/shifter/rol_32/ML_int[4][15] ), .S(
        \dp/ex_stage/alu/shifter/rol_32/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N70 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U16  ( .A(\dp/ex_stage/muxB_out [0]), 
        .Z(\dp/ex_stage/alu/shifter/ror_30/n3 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U15  ( .A(\dp/ex_stage/muxB_out [0]), 
        .Z(\dp/ex_stage/alu/shifter/ror_30/n1 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U14  ( .A(\dp/ex_stage/muxB_out [0]), 
        .Z(\dp/ex_stage/alu/shifter/ror_30/n2 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U13  ( .A(\dp/ex_stage/alu/n27 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n9 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U12  ( .A(\dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n12 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U11  ( .A(\dp/ex_stage/alu/n25 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n6 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U10  ( .A(\dp/ex_stage/alu/n27 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n7 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U9  ( .A(\dp/ex_stage/alu/n27 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n8 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U8  ( .A(\dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n10 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U7  ( .A(\dp/ex_stage/alu/n29 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n11 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U6  ( .A(\dp/ex_stage/alu/n25 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n4 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U5  ( .A(\dp/ex_stage/alu/n25 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n5 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U4  ( .A(
        \dp/ex_stage/alu/shifter/n99 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n15 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U3  ( .A(
        \dp/ex_stage/alu/shifter/n99 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n13 ) );
  BUF_X1 \dp/ex_stage/alu/shifter/ror_30/U2  ( .A(
        \dp/ex_stage/alu/shifter/n99 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/n14 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_0  ( .A(
        \dp/ex_stage/alu/shifter/N202 ), .B(\dp/ex_stage/muxA_out [1]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][0] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_1_0  ( .A(
        \dp/ex_stage/muxA_out [1]), .B(\dp/ex_stage/muxA_out [2]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_2_0  ( .A(
        \dp/ex_stage/muxA_out [2]), .B(\dp/ex_stage/muxA_out [3]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_3_0  ( .A(
        \dp/ex_stage/muxA_out [3]), .B(\dp/ex_stage/muxA_out [4]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_4_0  ( .A(
        \dp/ex_stage/muxA_out [4]), .B(\dp/ex_stage/muxA_out [5]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_5_0  ( .A(
        \dp/ex_stage/muxA_out [5]), .B(\dp/ex_stage/muxA_out [6]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_6_0  ( .A(
        \dp/ex_stage/muxA_out [6]), .B(\dp/ex_stage/muxA_out [7]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_7_0  ( .A(
        \dp/ex_stage/muxA_out [7]), .B(\dp/ex_stage/muxA_out [8]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_8_0  ( .A(
        \dp/ex_stage/muxA_out [8]), .B(\dp/ex_stage/muxA_out [9]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_9_0  ( .A(
        \dp/ex_stage/muxA_out [9]), .B(\dp/ex_stage/muxA_out [10]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_10_0  ( .A(
        \dp/ex_stage/muxA_out [10]), .B(\dp/ex_stage/muxA_out [11]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n1 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_11_0  ( .A(
        \dp/ex_stage/muxA_out [11]), .B(\dp/ex_stage/alu/n34 ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_12_0  ( .A(
        \dp/ex_stage/alu/n34 ), .B(\dp/ex_stage/muxA_out [13]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_13_0  ( .A(
        \dp/ex_stage/muxA_out [13]), .B(\dp/ex_stage/alu/n37 ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_14_0  ( .A(
        \dp/ex_stage/alu/n37 ), .B(\dp/ex_stage/muxA_out [15]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_15_0  ( .A(
        \dp/ex_stage/muxA_out [15]), .B(\dp/ex_stage/muxA_out [16]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_16_0  ( .A(
        \dp/ex_stage/muxA_out [16]), .B(\dp/ex_stage/muxA_out [17]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_17_0  ( .A(
        \dp/ex_stage/muxA_out [17]), .B(\dp/ex_stage/muxA_out [18]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_18_0  ( .A(
        \dp/ex_stage/muxA_out [18]), .B(\dp/ex_stage/muxA_out [19]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_19_0  ( .A(
        \dp/ex_stage/muxA_out [19]), .B(\dp/ex_stage/muxA_out [20]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_20_0  ( .A(
        \dp/ex_stage/muxA_out [20]), .B(\dp/ex_stage/muxA_out [21]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_21_0  ( .A(
        \dp/ex_stage/muxA_out [21]), .B(\dp/ex_stage/alu/n43 ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n2 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_22_0  ( .A(
        \dp/ex_stage/alu/n43 ), .B(\dp/ex_stage/alu/n45 ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_23_0  ( .A(
        \dp/ex_stage/alu/n45 ), .B(\dp/ex_stage/muxA_out [24]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_24_0  ( .A(
        \dp/ex_stage/muxA_out [24]), .B(\dp/ex_stage/muxA_out [25]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_25_0  ( .A(
        \dp/ex_stage/muxA_out [25]), .B(\dp/ex_stage/muxA_out [26]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_26_0  ( .A(
        \dp/ex_stage/muxA_out [26]), .B(\dp/ex_stage/muxA_out [27]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_27_0  ( .A(
        \dp/ex_stage/muxA_out [27]), .B(\dp/ex_stage/muxA_out [28]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_28_0  ( .A(
        \dp/ex_stage/muxA_out [28]), .B(\dp/ex_stage/muxA_out [29]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_29_0  ( .A(
        \dp/ex_stage/muxA_out [29]), .B(\dp/ex_stage/muxA_out [30]), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_30_0  ( .A(
        \dp/ex_stage/muxA_out [30]), .B(\dp/ex_stage/alu/shifter/N136 ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_0_31_0  ( .A(
        \dp/ex_stage/alu/shifter/N136 ), .B(\dp/ex_stage/alu/shifter/N202 ), 
        .S(\dp/ex_stage/alu/shifter/ror_30/n3 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][0] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][2] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][0] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_1  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][1] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][3] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_2_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][2] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][4] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_3_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][3] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][5] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_4_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][4] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][6] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_5_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][5] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][7] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_6_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][6] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][8] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_7_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][7] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][9] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_8_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][8] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][10] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_9_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][9] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][11] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_10_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][10] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][12] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n4 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_11_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][11] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][13] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_12_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][12] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][14] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_13_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][13] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][15] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_14_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][14] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][16] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_15_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][15] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][17] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_16_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][16] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][18] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_17_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][17] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][19] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_18_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][18] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][20] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_19_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][19] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][21] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_20_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][20] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][22] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_21_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][21] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][23] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n5 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_22_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][22] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][24] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_23_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][23] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][25] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_24_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][24] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][26] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_25_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][25] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][27] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_26_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][26] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][28] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_27_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][27] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][29] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_28_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][28] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][30] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_29_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][29] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][31] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_30_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][30] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][0] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_1_31_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][31] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[1][1] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n6 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][0] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][4] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][0] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_1  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][1] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][5] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_2  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][2] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][6] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_3  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][3] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][7] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_4_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][4] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][8] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_5_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][5] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][9] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_6_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][6] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][10] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_7_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][7] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][11] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_8_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][8] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][12] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_9_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][9] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][13] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_10_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][10] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][14] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n7 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_11_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][11] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][15] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_12_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][12] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][16] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_13_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][13] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][17] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_14_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][14] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][18] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_15_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][15] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][19] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_16_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][16] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][20] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_17_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][17] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][21] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_18_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][18] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][22] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_19_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][19] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][23] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_20_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][20] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][24] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_21_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][21] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][25] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n8 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_22_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][22] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][26] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_23_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][23] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][27] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_24_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][24] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][28] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_25_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][25] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][29] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_26_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][26] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][30] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_27_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][27] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][31] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_28_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][28] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][0] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_29_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][29] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][1] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_30_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][30] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][2] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_2_31_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][31] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[2][3] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n9 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][0] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][8] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][0] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_1  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][1] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][9] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][1] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_2  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][2] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][10] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][2] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_3  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][3] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][11] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][3] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_4  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][4] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][12] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][4] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_5  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][5] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][13] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][5] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_6  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][6] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][14] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][6] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_7  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][7] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][15] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][7] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_8_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][8] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][16] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][8] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_9_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][9] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][17] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][9] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_10_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][10] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][18] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n10 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][10] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_11_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][11] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][19] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][11] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_12_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][12] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][20] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][12] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_13_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][13] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][21] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][13] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_14_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][14] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][22] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][14] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_15_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][15] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][23] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][15] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_16_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][16] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][24] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][16] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_17_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][17] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][25] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][17] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_18_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][18] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][26] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][18] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_19_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][19] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][27] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][19] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_20_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][20] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][28] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][20] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_21_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][21] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][29] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n11 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][21] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_22_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][22] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][30] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][22] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_23_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][23] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][31] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][23] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_24_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][24] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][0] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][24] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_25_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][25] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][1] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][25] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_26_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][26] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][2] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][26] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_27_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][27] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][3] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][27] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_28_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][28] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][4] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][28] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_29_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][29] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][5] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][29] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_30_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][30] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][6] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][30] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_3_31_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][31] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[3][7] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n12 ), .Z(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][31] ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_0  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][0] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][16] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(\dp/ex_stage/alu/shifter/N7 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_1  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][1] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][17] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(\dp/ex_stage/alu/shifter/N8 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_2  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][2] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][18] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(\dp/ex_stage/alu/shifter/N9 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_3  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][3] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][19] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N10 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_4  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][4] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][20] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N11 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_5  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][5] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][21] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N12 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_6  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][6] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][22] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N13 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_7  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][7] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][23] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N14 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_8  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][8] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][24] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N15 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_9  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][9] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][25] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N16 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_10  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][10] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][26] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n13 ), .Z(
        \dp/ex_stage/alu/shifter/N17 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_11  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][11] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][27] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N18 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_12  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][12] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][28] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N19 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_13  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][13] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][29] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N20 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_14  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][14] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][30] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N21 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_15  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][15] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][31] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N22 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_16  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][16] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][0] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N23 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_17  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][17] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][1] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N24 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_18  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][18] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][2] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N25 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_19  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][19] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][3] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N26 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_20  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][20] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][4] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N27 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_21  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][21] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][5] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n14 ), .Z(
        \dp/ex_stage/alu/shifter/N28 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_22  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][22] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][6] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N29 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_23  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][23] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][7] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N30 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_24  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][24] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][8] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N31 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_25  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][25] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][9] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N32 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_26  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][26] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][10] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N33 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_27  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][27] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][11] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N34 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_28  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][28] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][12] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N35 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_29  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][29] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][13] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N36 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_30  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][30] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][14] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N37 ) );
  MUX2_X1 \dp/ex_stage/alu/shifter/ror_30/M1_4_31  ( .A(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][31] ), .B(
        \dp/ex_stage/alu/shifter/ror_30/MR_int[4][15] ), .S(
        \dp/ex_stage/alu/shifter/ror_30/n15 ), .Z(
        \dp/ex_stage/alu/shifter/N38 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U112  ( .A1(\dp/ex_stage/alu/n29 ), .A2(
        \dp/ex_stage/alu/r61/n16 ), .ZN(\dp/ex_stage/alu/r61/n106 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U111  ( .A1(\dp/ex_stage/muxB_out [6]), .A2(
        \dp/ex_stage/alu/r61/n20 ), .ZN(\dp/ex_stage/alu/r61/n103 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U110  ( .A1(\dp/ex_stage/muxB_out [5]), .A2(
        \dp/ex_stage/alu/r61/n19 ), .ZN(\dp/ex_stage/alu/r61/n102 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U109  ( .A1(\dp/ex_stage/muxB_out [8]), .A2(
        \dp/ex_stage/alu/r61/n22 ), .ZN(\dp/ex_stage/alu/r61/n99 ) );
  AND4_X1 \dp/ex_stage/alu/r61/U108  ( .A1(\dp/ex_stage/alu/r61/n106 ), .A2(
        \dp/ex_stage/alu/r61/n103 ), .A3(\dp/ex_stage/alu/r61/n102 ), .A4(
        \dp/ex_stage/alu/r61/n99 ), .ZN(\dp/ex_stage/alu/r61/n37 ) );
  AND2_X1 \dp/ex_stage/alu/r61/U107  ( .A1(\dp/ex_stage/muxB_out [31]), .A2(
        \dp/ex_stage/alu/r61/n35 ), .ZN(\dp/ex_stage/alu/r61/n72 ) );
  OR2_X1 \dp/ex_stage/alu/r61/U106  ( .A1(\dp/ex_stage/alu/r61/n36 ), .A2(
        \dp/ex_stage/muxA_out [30]), .ZN(\dp/ex_stage/alu/r61/n47 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U105  ( .A1(\dp/ex_stage/muxB_out [29]), .A2(
        \dp/ex_stage/alu/r61/n34 ), .ZN(\dp/ex_stage/alu/r61/n46 ) );
  AND2_X1 \dp/ex_stage/alu/r61/U104  ( .A1(\dp/ex_stage/alu/r61/n47 ), .A2(
        \dp/ex_stage/alu/r61/n46 ), .ZN(\dp/ex_stage/alu/r61/n76 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U103  ( .A1(\dp/ex_stage/muxB_out [27]), .A2(
        \dp/ex_stage/alu/r61/n32 ), .ZN(\dp/ex_stage/alu/r61/n48 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U102  ( .A1(\dp/ex_stage/muxB_out [28]), .A2(
        \dp/ex_stage/alu/r61/n33 ), .ZN(\dp/ex_stage/alu/r61/n50 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U101  ( .A1(\dp/ex_stage/muxB_out [25]), .A2(
        \dp/ex_stage/alu/r61/n30 ), .ZN(\dp/ex_stage/alu/r61/n51 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U100  ( .A1(\dp/ex_stage/muxB_out [26]), .A2(
        \dp/ex_stage/alu/r61/n31 ), .ZN(\dp/ex_stage/alu/r61/n52 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U99  ( .A1(\dp/ex_stage/muxB_out [23]), .A2(
        \dp/ex_stage/alu/r61/n11 ), .ZN(\dp/ex_stage/alu/r61/n53 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U98  ( .A1(\dp/ex_stage/muxB_out [24]), .A2(
        \dp/ex_stage/alu/r61/n29 ), .ZN(\dp/ex_stage/alu/r61/n54 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U97  ( .A1(\dp/ex_stage/muxB_out [21]), .A2(
        \dp/ex_stage/alu/r61/n9 ), .ZN(\dp/ex_stage/alu/r61/n55 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U96  ( .A1(\dp/ex_stage/muxB_out [22]), .A2(
        \dp/ex_stage/alu/r61/n10 ), .ZN(\dp/ex_stage/alu/r61/n56 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U95  ( .A1(\dp/ex_stage/muxB_out [19]), .A2(
        \dp/ex_stage/alu/r61/n27 ), .ZN(\dp/ex_stage/alu/r61/n57 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U94  ( .A1(\dp/ex_stage/muxB_out [20]), .A2(
        \dp/ex_stage/alu/r61/n28 ), .ZN(\dp/ex_stage/alu/r61/n58 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U93  ( .A1(\dp/ex_stage/muxB_out [17]), .A2(
        \dp/ex_stage/alu/r61/n8 ), .ZN(\dp/ex_stage/alu/r61/n59 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U92  ( .A1(\dp/ex_stage/muxB_out [18]), .A2(
        \dp/ex_stage/alu/r61/n26 ), .ZN(\dp/ex_stage/alu/r61/n60 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U91  ( .A1(\dp/ex_stage/muxB_out [15]), .A2(
        \dp/ex_stage/alu/r61/n6 ), .ZN(\dp/ex_stage/alu/r61/n61 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U90  ( .A1(\dp/ex_stage/muxB_out [16]), .A2(
        \dp/ex_stage/alu/r61/n7 ), .ZN(\dp/ex_stage/alu/r61/n64 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U89  ( .A1(\dp/ex_stage/muxB_out [13]), .A2(
        \dp/ex_stage/alu/r61/n4 ), .ZN(\dp/ex_stage/alu/r61/n65 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U88  ( .A1(\dp/ex_stage/muxB_out [14]), .A2(
        \dp/ex_stage/alu/r61/n5 ), .ZN(\dp/ex_stage/alu/r61/n66 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U87  ( .A1(\dp/ex_stage/muxB_out [11]), .A2(
        \dp/ex_stage/alu/r61/n25 ), .ZN(\dp/ex_stage/alu/r61/n67 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U86  ( .A1(\dp/ex_stage/muxB_out [12]), .A2(
        \dp/ex_stage/alu/r61/n3 ), .ZN(\dp/ex_stage/alu/r61/n68 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U85  ( .A1(\dp/ex_stage/muxB_out [9]), .A2(
        \dp/ex_stage/alu/r61/n23 ), .ZN(\dp/ex_stage/alu/r61/n69 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U84  ( .A1(\dp/ex_stage/muxB_out [10]), .A2(
        \dp/ex_stage/alu/r61/n24 ), .ZN(\dp/ex_stage/alu/r61/n70 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U83  ( .A1(\dp/ex_stage/muxB_out [7]), .A2(
        \dp/ex_stage/alu/r61/n21 ), .ZN(\dp/ex_stage/alu/r61/n71 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U82  ( .A1(\dp/ex_stage/alu/n31 ), .A2(
        \dp/ex_stage/alu/r61/n18 ), .ZN(\dp/ex_stage/alu/r61/n73 ) );
  NOR2_X1 \dp/ex_stage/alu/r61/U81  ( .A1(\dp/ex_stage/alu/r61/n13 ), .A2(
        \dp/ex_stage/muxB_out [0]), .ZN(\dp/ex_stage/alu/r61/n110 ) );
  AND2_X1 \dp/ex_stage/alu/r61/U80  ( .A1(\dp/ex_stage/alu/r61/n110 ), .A2(
        \dp/ex_stage/muxA_out [1]), .ZN(\dp/ex_stage/alu/r61/n109 ) );
  NAND2_X1 \dp/ex_stage/alu/r61/U79  ( .A1(\dp/ex_stage/alu/n27 ), .A2(
        \dp/ex_stage/alu/r61/n15 ), .ZN(\dp/ex_stage/alu/r61/n74 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U78  ( .B1(\dp/ex_stage/alu/r61/n109 ), .B2(
        \dp/ex_stage/alu/r61/n1 ), .C1(\dp/ex_stage/muxA_out [1]), .C2(
        \dp/ex_stage/alu/r61/n110 ), .A(\dp/ex_stage/alu/r61/n74 ), .ZN(
        \dp/ex_stage/alu/r61/n108 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U77  ( .B1(\dp/ex_stage/alu/n27 ), .B2(
        \dp/ex_stage/alu/r61/n15 ), .C1(\dp/ex_stage/alu/n29 ), .C2(
        \dp/ex_stage/alu/r61/n16 ), .A(\dp/ex_stage/alu/r61/n108 ), .ZN(
        \dp/ex_stage/alu/r61/n107 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U76  ( .A1(\dp/ex_stage/alu/r61/n106 ), .A2(
        \dp/ex_stage/alu/r61/n73 ), .A3(\dp/ex_stage/alu/r61/n107 ), .ZN(
        \dp/ex_stage/alu/r61/n105 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U75  ( .B1(\dp/ex_stage/alu/n31 ), .B2(
        \dp/ex_stage/alu/r61/n18 ), .C1(\dp/ex_stage/muxB_out [5]), .C2(
        \dp/ex_stage/alu/r61/n19 ), .A(\dp/ex_stage/alu/r61/n105 ), .ZN(
        \dp/ex_stage/alu/r61/n104 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U74  ( .A1(\dp/ex_stage/alu/r61/n102 ), .A2(
        \dp/ex_stage/alu/r61/n103 ), .A3(\dp/ex_stage/alu/r61/n104 ), .ZN(
        \dp/ex_stage/alu/r61/n101 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U73  ( .B1(\dp/ex_stage/muxB_out [6]), .B2(
        \dp/ex_stage/alu/r61/n20 ), .C1(\dp/ex_stage/muxB_out [7]), .C2(
        \dp/ex_stage/alu/r61/n21 ), .A(\dp/ex_stage/alu/r61/n101 ), .ZN(
        \dp/ex_stage/alu/r61/n100 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U72  ( .A1(\dp/ex_stage/alu/r61/n71 ), .A2(
        \dp/ex_stage/alu/r61/n99 ), .A3(\dp/ex_stage/alu/r61/n100 ), .ZN(
        \dp/ex_stage/alu/r61/n98 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U71  ( .B1(\dp/ex_stage/muxB_out [8]), .B2(
        \dp/ex_stage/alu/r61/n22 ), .C1(\dp/ex_stage/muxB_out [9]), .C2(
        \dp/ex_stage/alu/r61/n23 ), .A(\dp/ex_stage/alu/r61/n98 ), .ZN(
        \dp/ex_stage/alu/r61/n97 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U70  ( .A1(\dp/ex_stage/alu/r61/n69 ), .A2(
        \dp/ex_stage/alu/r61/n70 ), .A3(\dp/ex_stage/alu/r61/n97 ), .ZN(
        \dp/ex_stage/alu/r61/n96 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U69  ( .B1(\dp/ex_stage/muxB_out [10]), .B2(
        \dp/ex_stage/alu/r61/n24 ), .C1(\dp/ex_stage/muxB_out [11]), .C2(
        \dp/ex_stage/alu/r61/n25 ), .A(\dp/ex_stage/alu/r61/n96 ), .ZN(
        \dp/ex_stage/alu/r61/n95 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U68  ( .A1(\dp/ex_stage/alu/r61/n67 ), .A2(
        \dp/ex_stage/alu/r61/n68 ), .A3(\dp/ex_stage/alu/r61/n95 ), .ZN(
        \dp/ex_stage/alu/r61/n94 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U67  ( .B1(\dp/ex_stage/muxB_out [12]), .B2(
        \dp/ex_stage/alu/r61/n3 ), .C1(\dp/ex_stage/muxB_out [13]), .C2(
        \dp/ex_stage/alu/r61/n4 ), .A(\dp/ex_stage/alu/r61/n94 ), .ZN(
        \dp/ex_stage/alu/r61/n93 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U66  ( .A1(\dp/ex_stage/alu/r61/n65 ), .A2(
        \dp/ex_stage/alu/r61/n66 ), .A3(\dp/ex_stage/alu/r61/n93 ), .ZN(
        \dp/ex_stage/alu/r61/n92 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U65  ( .B1(\dp/ex_stage/muxB_out [14]), .B2(
        \dp/ex_stage/alu/r61/n5 ), .C1(\dp/ex_stage/muxB_out [15]), .C2(
        \dp/ex_stage/alu/r61/n6 ), .A(\dp/ex_stage/alu/r61/n92 ), .ZN(
        \dp/ex_stage/alu/r61/n91 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U64  ( .A1(\dp/ex_stage/alu/r61/n61 ), .A2(
        \dp/ex_stage/alu/r61/n64 ), .A3(\dp/ex_stage/alu/r61/n91 ), .ZN(
        \dp/ex_stage/alu/r61/n90 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U63  ( .B1(\dp/ex_stage/muxB_out [16]), .B2(
        \dp/ex_stage/alu/r61/n7 ), .C1(\dp/ex_stage/muxB_out [17]), .C2(
        \dp/ex_stage/alu/r61/n8 ), .A(\dp/ex_stage/alu/r61/n90 ), .ZN(
        \dp/ex_stage/alu/r61/n89 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U62  ( .A1(\dp/ex_stage/alu/r61/n59 ), .A2(
        \dp/ex_stage/alu/r61/n60 ), .A3(\dp/ex_stage/alu/r61/n89 ), .ZN(
        \dp/ex_stage/alu/r61/n88 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U61  ( .B1(\dp/ex_stage/muxB_out [18]), .B2(
        \dp/ex_stage/alu/r61/n26 ), .C1(\dp/ex_stage/muxB_out [19]), .C2(
        \dp/ex_stage/alu/r61/n27 ), .A(\dp/ex_stage/alu/r61/n88 ), .ZN(
        \dp/ex_stage/alu/r61/n87 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U60  ( .A1(\dp/ex_stage/alu/r61/n57 ), .A2(
        \dp/ex_stage/alu/r61/n58 ), .A3(\dp/ex_stage/alu/r61/n87 ), .ZN(
        \dp/ex_stage/alu/r61/n86 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U59  ( .B1(\dp/ex_stage/muxB_out [20]), .B2(
        \dp/ex_stage/alu/r61/n28 ), .C1(\dp/ex_stage/muxB_out [21]), .C2(
        \dp/ex_stage/alu/r61/n9 ), .A(\dp/ex_stage/alu/r61/n86 ), .ZN(
        \dp/ex_stage/alu/r61/n85 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U58  ( .A1(\dp/ex_stage/alu/r61/n55 ), .A2(
        \dp/ex_stage/alu/r61/n56 ), .A3(\dp/ex_stage/alu/r61/n85 ), .ZN(
        \dp/ex_stage/alu/r61/n84 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U57  ( .B1(\dp/ex_stage/muxB_out [22]), .B2(
        \dp/ex_stage/alu/r61/n10 ), .C1(\dp/ex_stage/muxB_out [23]), .C2(
        \dp/ex_stage/alu/r61/n11 ), .A(\dp/ex_stage/alu/r61/n84 ), .ZN(
        \dp/ex_stage/alu/r61/n83 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U56  ( .A1(\dp/ex_stage/alu/r61/n53 ), .A2(
        \dp/ex_stage/alu/r61/n54 ), .A3(\dp/ex_stage/alu/r61/n83 ), .ZN(
        \dp/ex_stage/alu/r61/n82 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U55  ( .B1(\dp/ex_stage/muxB_out [24]), .B2(
        \dp/ex_stage/alu/r61/n29 ), .C1(\dp/ex_stage/muxB_out [25]), .C2(
        \dp/ex_stage/alu/r61/n30 ), .A(\dp/ex_stage/alu/r61/n82 ), .ZN(
        \dp/ex_stage/alu/r61/n81 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U54  ( .A1(\dp/ex_stage/alu/r61/n51 ), .A2(
        \dp/ex_stage/alu/r61/n52 ), .A3(\dp/ex_stage/alu/r61/n81 ), .ZN(
        \dp/ex_stage/alu/r61/n80 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U53  ( .B1(\dp/ex_stage/muxB_out [26]), .B2(
        \dp/ex_stage/alu/r61/n31 ), .C1(\dp/ex_stage/muxB_out [27]), .C2(
        \dp/ex_stage/alu/r61/n32 ), .A(\dp/ex_stage/alu/r61/n80 ), .ZN(
        \dp/ex_stage/alu/r61/n79 ) );
  NAND3_X1 \dp/ex_stage/alu/r61/U52  ( .A1(\dp/ex_stage/alu/r61/n48 ), .A2(
        \dp/ex_stage/alu/r61/n50 ), .A3(\dp/ex_stage/alu/r61/n79 ), .ZN(
        \dp/ex_stage/alu/r61/n78 ) );
  OAI221_X1 \dp/ex_stage/alu/r61/U51  ( .B1(\dp/ex_stage/muxB_out [28]), .B2(
        \dp/ex_stage/alu/r61/n33 ), .C1(\dp/ex_stage/muxB_out [29]), .C2(
        \dp/ex_stage/alu/r61/n34 ), .A(\dp/ex_stage/alu/r61/n78 ), .ZN(
        \dp/ex_stage/alu/r61/n77 ) );
  AOI22_X1 \dp/ex_stage/alu/r61/U50  ( .A1(\dp/ex_stage/muxA_out [30]), .A2(
        \dp/ex_stage/alu/r61/n36 ), .B1(\dp/ex_stage/alu/r61/n76 ), .B2(
        \dp/ex_stage/alu/r61/n77 ), .ZN(\dp/ex_stage/alu/r61/n75 ) );
  OAI22_X1 \dp/ex_stage/alu/r61/U49  ( .A1(\dp/ex_stage/muxB_out [31]), .A2(
        \dp/ex_stage/alu/r61/n35 ), .B1(\dp/ex_stage/alu/r61/n72 ), .B2(
        \dp/ex_stage/alu/r61/n75 ), .ZN(\dp/ex_stage/alu/N21 ) );
  NOR4_X1 \dp/ex_stage/alu/r61/U48  ( .A1(\dp/ex_stage/alu/N21 ), .A2(
        \dp/ex_stage/alu/r61/n72 ), .A3(\dp/ex_stage/alu/r61/n14 ), .A4(
        \dp/ex_stage/alu/r61/n17 ), .ZN(\dp/ex_stage/alu/r61/n38 ) );
  NAND4_X1 \dp/ex_stage/alu/r61/U47  ( .A1(\dp/ex_stage/alu/r61/n68 ), .A2(
        \dp/ex_stage/alu/r61/n69 ), .A3(\dp/ex_stage/alu/r61/n70 ), .A4(
        \dp/ex_stage/alu/r61/n71 ), .ZN(\dp/ex_stage/alu/r61/n62 ) );
  NAND4_X1 \dp/ex_stage/alu/r61/U46  ( .A1(\dp/ex_stage/alu/r61/n64 ), .A2(
        \dp/ex_stage/alu/r61/n65 ), .A3(\dp/ex_stage/alu/r61/n66 ), .A4(
        \dp/ex_stage/alu/r61/n67 ), .ZN(\dp/ex_stage/alu/r61/n63 ) );
  NOR2_X1 \dp/ex_stage/alu/r61/U45  ( .A1(\dp/ex_stage/alu/r61/n62 ), .A2(
        \dp/ex_stage/alu/r61/n63 ), .ZN(\dp/ex_stage/alu/r61/n39 ) );
  NAND4_X1 \dp/ex_stage/alu/r61/U44  ( .A1(\dp/ex_stage/alu/r61/n58 ), .A2(
        \dp/ex_stage/alu/r61/n59 ), .A3(\dp/ex_stage/alu/r61/n60 ), .A4(
        \dp/ex_stage/alu/r61/n61 ), .ZN(\dp/ex_stage/alu/r61/n41 ) );
  NAND4_X1 \dp/ex_stage/alu/r61/U43  ( .A1(\dp/ex_stage/alu/r61/n54 ), .A2(
        \dp/ex_stage/alu/r61/n55 ), .A3(\dp/ex_stage/alu/r61/n56 ), .A4(
        \dp/ex_stage/alu/r61/n57 ), .ZN(\dp/ex_stage/alu/r61/n42 ) );
  NAND4_X1 \dp/ex_stage/alu/r61/U42  ( .A1(\dp/ex_stage/alu/r61/n50 ), .A2(
        \dp/ex_stage/alu/r61/n51 ), .A3(\dp/ex_stage/alu/r61/n52 ), .A4(
        \dp/ex_stage/alu/r61/n53 ), .ZN(\dp/ex_stage/alu/r61/n43 ) );
  AND2_X1 \dp/ex_stage/alu/r61/U41  ( .A1(\dp/ex_stage/muxB_out [0]), .A2(
        \dp/ex_stage/alu/r61/n13 ), .ZN(\dp/ex_stage/alu/r61/n49 ) );
  OAI22_X1 \dp/ex_stage/alu/r61/U40  ( .A1(\dp/ex_stage/alu/r61/n49 ), .A2(
        \dp/ex_stage/alu/r61/n2 ), .B1(\dp/ex_stage/alu/n25 ), .B2(
        \dp/ex_stage/alu/r61/n49 ), .ZN(\dp/ex_stage/alu/r61/n45 ) );
  NAND4_X1 \dp/ex_stage/alu/r61/U39  ( .A1(\dp/ex_stage/alu/r61/n45 ), .A2(
        \dp/ex_stage/alu/r61/n46 ), .A3(\dp/ex_stage/alu/r61/n47 ), .A4(
        \dp/ex_stage/alu/r61/n48 ), .ZN(\dp/ex_stage/alu/r61/n44 ) );
  NOR4_X1 \dp/ex_stage/alu/r61/U38  ( .A1(\dp/ex_stage/alu/r61/n41 ), .A2(
        \dp/ex_stage/alu/r61/n42 ), .A3(\dp/ex_stage/alu/r61/n43 ), .A4(
        \dp/ex_stage/alu/r61/n44 ), .ZN(\dp/ex_stage/alu/r61/n40 ) );
  NAND4_X1 \dp/ex_stage/alu/r61/U37  ( .A1(\dp/ex_stage/alu/r61/n37 ), .A2(
        \dp/ex_stage/alu/r61/n38 ), .A3(\dp/ex_stage/alu/r61/n39 ), .A4(
        \dp/ex_stage/alu/r61/n40 ), .ZN(\dp/ex_stage/alu/N18 ) );
  INV_X1 \dp/ex_stage/alu/r61/U36  ( .A(\dp/ex_stage/alu/n45 ), .ZN(
        \dp/ex_stage/alu/r61/n11 ) );
  INV_X1 \dp/ex_stage/alu/r61/U35  ( .A(\dp/ex_stage/alu/n43 ), .ZN(
        \dp/ex_stage/alu/r61/n10 ) );
  INV_X1 \dp/ex_stage/alu/r61/U34  ( .A(\dp/ex_stage/muxA_out [21]), .ZN(
        \dp/ex_stage/alu/r61/n9 ) );
  INV_X1 \dp/ex_stage/alu/r61/U33  ( .A(\dp/ex_stage/muxA_out [17]), .ZN(
        \dp/ex_stage/alu/r61/n8 ) );
  INV_X1 \dp/ex_stage/alu/r61/U32  ( .A(\dp/ex_stage/muxA_out [16]), .ZN(
        \dp/ex_stage/alu/r61/n7 ) );
  INV_X1 \dp/ex_stage/alu/r61/U31  ( .A(\dp/ex_stage/muxA_out [15]), .ZN(
        \dp/ex_stage/alu/r61/n6 ) );
  INV_X1 \dp/ex_stage/alu/r61/U30  ( .A(\dp/ex_stage/alu/n37 ), .ZN(
        \dp/ex_stage/alu/r61/n5 ) );
  INV_X1 \dp/ex_stage/alu/r61/U29  ( .A(\dp/ex_stage/muxA_out [13]), .ZN(
        \dp/ex_stage/alu/r61/n4 ) );
  INV_X1 \dp/ex_stage/alu/r61/U28  ( .A(\dp/ex_stage/alu/n34 ), .ZN(
        \dp/ex_stage/alu/r61/n3 ) );
  INV_X1 \dp/ex_stage/alu/r61/U27  ( .A(\dp/ex_stage/muxA_out [1]), .ZN(
        \dp/ex_stage/alu/r61/n2 ) );
  INV_X1 \dp/ex_stage/alu/r61/U26  ( .A(\dp/ex_stage/alu/n25 ), .ZN(
        \dp/ex_stage/alu/r61/n1 ) );
  INV_X1 \dp/ex_stage/alu/r61/U25  ( .A(\dp/ex_stage/muxB_out [30]), .ZN(
        \dp/ex_stage/alu/r61/n36 ) );
  INV_X1 \dp/ex_stage/alu/r61/U24  ( .A(\dp/ex_stage/alu/shifter/N136 ), .ZN(
        \dp/ex_stage/alu/r61/n35 ) );
  INV_X1 \dp/ex_stage/alu/r61/U23  ( .A(\dp/ex_stage/muxA_out [19]), .ZN(
        \dp/ex_stage/alu/r61/n27 ) );
  INV_X1 \dp/ex_stage/alu/r61/U22  ( .A(\dp/ex_stage/muxA_out [20]), .ZN(
        \dp/ex_stage/alu/r61/n28 ) );
  INV_X1 \dp/ex_stage/alu/r61/U21  ( .A(\dp/ex_stage/muxA_out [29]), .ZN(
        \dp/ex_stage/alu/r61/n34 ) );
  INV_X1 \dp/ex_stage/alu/r61/U20  ( .A(\dp/ex_stage/muxA_out [18]), .ZN(
        \dp/ex_stage/alu/r61/n26 ) );
  INV_X1 \dp/ex_stage/alu/r61/U19  ( .A(\dp/ex_stage/muxA_out [27]), .ZN(
        \dp/ex_stage/alu/r61/n32 ) );
  INV_X1 \dp/ex_stage/alu/r61/U18  ( .A(\dp/ex_stage/muxA_out [25]), .ZN(
        \dp/ex_stage/alu/r61/n30 ) );
  INV_X1 \dp/ex_stage/alu/r61/U17  ( .A(\dp/ex_stage/muxA_out [28]), .ZN(
        \dp/ex_stage/alu/r61/n33 ) );
  INV_X1 \dp/ex_stage/alu/r61/U16  ( .A(\dp/ex_stage/muxA_out [26]), .ZN(
        \dp/ex_stage/alu/r61/n31 ) );
  INV_X1 \dp/ex_stage/alu/r61/U15  ( .A(\dp/ex_stage/muxA_out [24]), .ZN(
        \dp/ex_stage/alu/r61/n29 ) );
  INV_X1 \dp/ex_stage/alu/r61/U14  ( .A(\dp/ex_stage/alu/N18 ), .ZN(
        \dp/ex_stage/alu/N19 ) );
  INV_X1 \dp/ex_stage/alu/r61/U13  ( .A(\dp/ex_stage/muxA_out [5]), .ZN(
        \dp/ex_stage/alu/r61/n19 ) );
  INV_X1 \dp/ex_stage/alu/r61/U12  ( .A(\dp/ex_stage/muxA_out [6]), .ZN(
        \dp/ex_stage/alu/r61/n20 ) );
  INV_X1 \dp/ex_stage/alu/r61/U11  ( .A(\dp/ex_stage/muxA_out [4]), .ZN(
        \dp/ex_stage/alu/r61/n18 ) );
  INV_X1 \dp/ex_stage/alu/r61/U10  ( .A(\dp/ex_stage/alu/shifter/N202 ), .ZN(
        \dp/ex_stage/alu/r61/n13 ) );
  INV_X1 \dp/ex_stage/alu/r61/U9  ( .A(\dp/ex_stage/muxA_out [3]), .ZN(
        \dp/ex_stage/alu/r61/n16 ) );
  INV_X1 \dp/ex_stage/alu/r61/U8  ( .A(\dp/ex_stage/muxA_out [9]), .ZN(
        \dp/ex_stage/alu/r61/n23 ) );
  INV_X1 \dp/ex_stage/alu/r61/U7  ( .A(\dp/ex_stage/muxA_out [11]), .ZN(
        \dp/ex_stage/alu/r61/n25 ) );
  INV_X1 \dp/ex_stage/alu/r61/U6  ( .A(\dp/ex_stage/muxA_out [7]), .ZN(
        \dp/ex_stage/alu/r61/n21 ) );
  INV_X1 \dp/ex_stage/alu/r61/U5  ( .A(\dp/ex_stage/muxA_out [2]), .ZN(
        \dp/ex_stage/alu/r61/n15 ) );
  INV_X1 \dp/ex_stage/alu/r61/U4  ( .A(\dp/ex_stage/muxA_out [10]), .ZN(
        \dp/ex_stage/alu/r61/n24 ) );
  INV_X1 \dp/ex_stage/alu/r61/U3  ( .A(\dp/ex_stage/muxA_out [8]), .ZN(
        \dp/ex_stage/alu/r61/n22 ) );
  INV_X1 \dp/ex_stage/alu/r61/U2  ( .A(\dp/ex_stage/alu/r61/n74 ), .ZN(
        \dp/ex_stage/alu/r61/n14 ) );
  INV_X1 \dp/ex_stage/alu/r61/U1  ( .A(\dp/ex_stage/alu/r61/n73 ), .ZN(
        \dp/ex_stage/alu/r61/n17 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U204  ( .A1(\dp/ex_stage/alu/r60/n64 ), .A2(
        \dp/ex_stage/muxB_out [31]), .ZN(\dp/ex_stage/alu/r60/n67 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U203  ( .A1(\dp/ex_stage/alu/r60/n16 ), .A2(
        \dp/ex_stage/muxB_out [0]), .ZN(\dp/ex_stage/alu/r60/n202 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U202  ( .A1(\dp/ex_stage/alu/r60/n202 ), .A2(
        \dp/ex_stage/alu/r60/n1 ), .ZN(\dp/ex_stage/alu/r60/n201 ) );
  OAI22_X1 \dp/ex_stage/alu/r60/U201  ( .A1(\dp/ex_stage/alu/r60/n201 ), .A2(
        \dp/ex_stage/muxA_out [1]), .B1(\dp/ex_stage/alu/r60/n1 ), .B2(
        \dp/ex_stage/alu/r60/n202 ), .ZN(\dp/ex_stage/alu/r60/n200 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U200  ( .A1(\dp/ex_stage/alu/r60/n18 ), .A2(
        \dp/ex_stage/alu/n27 ), .ZN(\dp/ex_stage/alu/r60/n199 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U199  ( .A1(\dp/ex_stage/alu/n27 ), .A2(
        \dp/ex_stage/alu/r60/n18 ), .ZN(\dp/ex_stage/alu/r60/n138 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U198  ( .A1(\dp/ex_stage/alu/r60/n199 ), .A2(
        \dp/ex_stage/alu/r60/n17 ), .ZN(\dp/ex_stage/alu/r60/n141 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U197  ( .B1(\dp/ex_stage/alu/r60/n12 ), .B2(
        \dp/ex_stage/alu/r60/n141 ), .A(\dp/ex_stage/alu/r60/n199 ), .ZN(
        \dp/ex_stage/alu/r60/n198 ) );
  OR2_X1 \dp/ex_stage/alu/r60/U196  ( .A1(\dp/ex_stage/alu/r60/n20 ), .A2(
        \dp/ex_stage/alu/n29 ), .ZN(\dp/ex_stage/alu/r60/n135 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U195  ( .A1(\dp/ex_stage/alu/n29 ), .A2(
        \dp/ex_stage/alu/r60/n20 ), .ZN(\dp/ex_stage/alu/r60/n137 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U194  ( .B1(\dp/ex_stage/alu/r60/n198 ), .B2(
        \dp/ex_stage/alu/r60/n135 ), .A(\dp/ex_stage/alu/r60/n19 ), .ZN(
        \dp/ex_stage/alu/r60/n196 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U193  ( .A1(\dp/ex_stage/alu/r60/n21 ), .A2(
        \dp/ex_stage/alu/n31 ), .ZN(\dp/ex_stage/alu/r60/n197 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U192  ( .A1(\dp/ex_stage/alu/n31 ), .A2(
        \dp/ex_stage/alu/r60/n21 ), .ZN(\dp/ex_stage/alu/r60/n143 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U191  ( .A1(\dp/ex_stage/alu/r60/n197 ), .A2(
        \dp/ex_stage/alu/r60/n143 ), .ZN(\dp/ex_stage/alu/r60/n136 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U190  ( .B1(\dp/ex_stage/alu/r60/n196 ), .B2(
        \dp/ex_stage/alu/r60/n136 ), .A(\dp/ex_stage/alu/r60/n197 ), .ZN(
        \dp/ex_stage/alu/r60/n195 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U189  ( .A1(\dp/ex_stage/alu/r60/n23 ), .A2(
        \dp/ex_stage/muxB_out [5]), .ZN(\dp/ex_stage/alu/r60/n133 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U188  ( .A1(\dp/ex_stage/muxB_out [5]), .A2(
        \dp/ex_stage/alu/r60/n23 ), .ZN(\dp/ex_stage/alu/r60/n144 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U187  ( .B1(\dp/ex_stage/alu/r60/n195 ), .B2(
        \dp/ex_stage/alu/r60/n22 ), .A(\dp/ex_stage/alu/r60/n144 ), .ZN(
        \dp/ex_stage/alu/r60/n193 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U186  ( .A1(\dp/ex_stage/alu/r60/n26 ), .A2(
        \dp/ex_stage/muxB_out [6]), .ZN(\dp/ex_stage/alu/r60/n194 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U185  ( .A1(\dp/ex_stage/muxB_out [6]), .A2(
        \dp/ex_stage/alu/r60/n26 ), .ZN(\dp/ex_stage/alu/r60/n129 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U184  ( .A1(\dp/ex_stage/alu/r60/n25 ), .A2(
        \dp/ex_stage/alu/r60/n129 ), .ZN(\dp/ex_stage/alu/r60/n132 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U183  ( .B1(\dp/ex_stage/alu/r60/n193 ), .B2(
        \dp/ex_stage/alu/r60/n24 ), .A(\dp/ex_stage/alu/r60/n194 ), .ZN(
        \dp/ex_stage/alu/r60/n192 ) );
  OR2_X1 \dp/ex_stage/alu/r60/U182  ( .A1(\dp/ex_stage/alu/r60/n28 ), .A2(
        \dp/ex_stage/muxB_out [7]), .ZN(\dp/ex_stage/alu/r60/n126 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U181  ( .A1(\dp/ex_stage/muxB_out [7]), .A2(
        \dp/ex_stage/alu/r60/n28 ), .ZN(\dp/ex_stage/alu/r60/n128 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U180  ( .B1(\dp/ex_stage/alu/r60/n192 ), .B2(
        \dp/ex_stage/alu/r60/n126 ), .A(\dp/ex_stage/alu/r60/n27 ), .ZN(
        \dp/ex_stage/alu/r60/n190 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U179  ( .A1(\dp/ex_stage/alu/r60/n29 ), .A2(
        \dp/ex_stage/muxB_out [8]), .ZN(\dp/ex_stage/alu/r60/n191 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U178  ( .A1(\dp/ex_stage/muxB_out [8]), .A2(
        \dp/ex_stage/alu/r60/n29 ), .ZN(\dp/ex_stage/alu/r60/n145 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U177  ( .A1(\dp/ex_stage/alu/r60/n191 ), .A2(
        \dp/ex_stage/alu/r60/n145 ), .ZN(\dp/ex_stage/alu/r60/n127 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U176  ( .B1(\dp/ex_stage/alu/r60/n190 ), .B2(
        \dp/ex_stage/alu/r60/n127 ), .A(\dp/ex_stage/alu/r60/n191 ), .ZN(
        \dp/ex_stage/alu/r60/n189 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U175  ( .A1(\dp/ex_stage/alu/r60/n31 ), .A2(
        \dp/ex_stage/muxB_out [9]), .ZN(\dp/ex_stage/alu/r60/n123 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U174  ( .A1(\dp/ex_stage/muxB_out [9]), .A2(
        \dp/ex_stage/alu/r60/n31 ), .ZN(\dp/ex_stage/alu/r60/n146 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U173  ( .B1(\dp/ex_stage/alu/r60/n189 ), .B2(
        \dp/ex_stage/alu/r60/n30 ), .A(\dp/ex_stage/alu/r60/n146 ), .ZN(
        \dp/ex_stage/alu/r60/n187 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U172  ( .A1(\dp/ex_stage/alu/r60/n34 ), .A2(
        \dp/ex_stage/muxB_out [10]), .ZN(\dp/ex_stage/alu/r60/n188 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U171  ( .A1(\dp/ex_stage/muxB_out [10]), .A2(
        \dp/ex_stage/alu/r60/n34 ), .ZN(\dp/ex_stage/alu/r60/n119 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U170  ( .A1(\dp/ex_stage/alu/r60/n33 ), .A2(
        \dp/ex_stage/alu/r60/n119 ), .ZN(\dp/ex_stage/alu/r60/n122 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U169  ( .B1(\dp/ex_stage/alu/r60/n187 ), .B2(
        \dp/ex_stage/alu/r60/n32 ), .A(\dp/ex_stage/alu/r60/n188 ), .ZN(
        \dp/ex_stage/alu/r60/n186 ) );
  OR2_X1 \dp/ex_stage/alu/r60/U168  ( .A1(\dp/ex_stage/alu/r60/n36 ), .A2(
        \dp/ex_stage/muxB_out [11]), .ZN(\dp/ex_stage/alu/r60/n116 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U167  ( .A1(\dp/ex_stage/muxB_out [11]), .A2(
        \dp/ex_stage/alu/r60/n36 ), .ZN(\dp/ex_stage/alu/r60/n118 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U166  ( .B1(\dp/ex_stage/alu/r60/n186 ), .B2(
        \dp/ex_stage/alu/r60/n116 ), .A(\dp/ex_stage/alu/r60/n35 ), .ZN(
        \dp/ex_stage/alu/r60/n184 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U165  ( .A1(\dp/ex_stage/alu/r60/n2 ), .A2(
        \dp/ex_stage/muxB_out [12]), .ZN(\dp/ex_stage/alu/r60/n185 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U164  ( .A1(\dp/ex_stage/muxB_out [12]), .A2(
        \dp/ex_stage/alu/r60/n2 ), .ZN(\dp/ex_stage/alu/r60/n147 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U163  ( .A1(\dp/ex_stage/alu/r60/n185 ), .A2(
        \dp/ex_stage/alu/r60/n147 ), .ZN(\dp/ex_stage/alu/r60/n117 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U162  ( .B1(\dp/ex_stage/alu/r60/n184 ), .B2(
        \dp/ex_stage/alu/r60/n117 ), .A(\dp/ex_stage/alu/r60/n185 ), .ZN(
        \dp/ex_stage/alu/r60/n183 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U161  ( .A1(\dp/ex_stage/alu/r60/n3 ), .A2(
        \dp/ex_stage/muxB_out [13]), .ZN(\dp/ex_stage/alu/r60/n113 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U160  ( .A1(\dp/ex_stage/muxB_out [13]), .A2(
        \dp/ex_stage/alu/r60/n3 ), .ZN(\dp/ex_stage/alu/r60/n148 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U159  ( .B1(\dp/ex_stage/alu/r60/n183 ), .B2(
        \dp/ex_stage/alu/r60/n37 ), .A(\dp/ex_stage/alu/r60/n148 ), .ZN(
        \dp/ex_stage/alu/r60/n181 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U158  ( .A1(\dp/ex_stage/alu/r60/n4 ), .A2(
        \dp/ex_stage/muxB_out [14]), .ZN(\dp/ex_stage/alu/r60/n182 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U157  ( .A1(\dp/ex_stage/muxB_out [14]), .A2(
        \dp/ex_stage/alu/r60/n4 ), .ZN(\dp/ex_stage/alu/r60/n109 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U156  ( .A1(\dp/ex_stage/alu/r60/n39 ), .A2(
        \dp/ex_stage/alu/r60/n109 ), .ZN(\dp/ex_stage/alu/r60/n112 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U155  ( .B1(\dp/ex_stage/alu/r60/n181 ), .B2(
        \dp/ex_stage/alu/r60/n38 ), .A(\dp/ex_stage/alu/r60/n182 ), .ZN(
        \dp/ex_stage/alu/r60/n180 ) );
  OR2_X1 \dp/ex_stage/alu/r60/U154  ( .A1(\dp/ex_stage/alu/r60/n5 ), .A2(
        \dp/ex_stage/muxB_out [15]), .ZN(\dp/ex_stage/alu/r60/n106 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U153  ( .A1(\dp/ex_stage/muxB_out [15]), .A2(
        \dp/ex_stage/alu/r60/n5 ), .ZN(\dp/ex_stage/alu/r60/n108 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U152  ( .B1(\dp/ex_stage/alu/r60/n180 ), .B2(
        \dp/ex_stage/alu/r60/n106 ), .A(\dp/ex_stage/alu/r60/n40 ), .ZN(
        \dp/ex_stage/alu/r60/n178 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U151  ( .A1(\dp/ex_stage/alu/r60/n6 ), .A2(
        \dp/ex_stage/muxB_out [16]), .ZN(\dp/ex_stage/alu/r60/n179 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U150  ( .A1(\dp/ex_stage/muxB_out [16]), .A2(
        \dp/ex_stage/alu/r60/n6 ), .ZN(\dp/ex_stage/alu/r60/n149 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U149  ( .A1(\dp/ex_stage/alu/r60/n179 ), .A2(
        \dp/ex_stage/alu/r60/n149 ), .ZN(\dp/ex_stage/alu/r60/n107 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U148  ( .B1(\dp/ex_stage/alu/r60/n178 ), .B2(
        \dp/ex_stage/alu/r60/n107 ), .A(\dp/ex_stage/alu/r60/n179 ), .ZN(
        \dp/ex_stage/alu/r60/n177 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U147  ( .A1(\dp/ex_stage/alu/r60/n7 ), .A2(
        \dp/ex_stage/muxB_out [17]), .ZN(\dp/ex_stage/alu/r60/n103 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U146  ( .A1(\dp/ex_stage/muxB_out [17]), .A2(
        \dp/ex_stage/alu/r60/n7 ), .ZN(\dp/ex_stage/alu/r60/n150 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U145  ( .B1(\dp/ex_stage/alu/r60/n177 ), .B2(
        \dp/ex_stage/alu/r60/n41 ), .A(\dp/ex_stage/alu/r60/n150 ), .ZN(
        \dp/ex_stage/alu/r60/n175 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U144  ( .A1(\dp/ex_stage/alu/r60/n44 ), .A2(
        \dp/ex_stage/muxB_out [18]), .ZN(\dp/ex_stage/alu/r60/n176 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U143  ( .A1(\dp/ex_stage/muxB_out [18]), .A2(
        \dp/ex_stage/alu/r60/n44 ), .ZN(\dp/ex_stage/alu/r60/n99 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U142  ( .A1(\dp/ex_stage/alu/r60/n43 ), .A2(
        \dp/ex_stage/alu/r60/n99 ), .ZN(\dp/ex_stage/alu/r60/n102 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U141  ( .B1(\dp/ex_stage/alu/r60/n175 ), .B2(
        \dp/ex_stage/alu/r60/n42 ), .A(\dp/ex_stage/alu/r60/n176 ), .ZN(
        \dp/ex_stage/alu/r60/n174 ) );
  OR2_X1 \dp/ex_stage/alu/r60/U140  ( .A1(\dp/ex_stage/alu/r60/n46 ), .A2(
        \dp/ex_stage/muxB_out [19]), .ZN(\dp/ex_stage/alu/r60/n96 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U139  ( .A1(\dp/ex_stage/muxB_out [19]), .A2(
        \dp/ex_stage/alu/r60/n46 ), .ZN(\dp/ex_stage/alu/r60/n98 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U138  ( .B1(\dp/ex_stage/alu/r60/n174 ), .B2(
        \dp/ex_stage/alu/r60/n96 ), .A(\dp/ex_stage/alu/r60/n45 ), .ZN(
        \dp/ex_stage/alu/r60/n172 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U137  ( .A1(\dp/ex_stage/alu/r60/n47 ), .A2(
        \dp/ex_stage/muxB_out [20]), .ZN(\dp/ex_stage/alu/r60/n173 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U136  ( .A1(\dp/ex_stage/muxB_out [20]), .A2(
        \dp/ex_stage/alu/r60/n47 ), .ZN(\dp/ex_stage/alu/r60/n151 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U135  ( .A1(\dp/ex_stage/alu/r60/n173 ), .A2(
        \dp/ex_stage/alu/r60/n151 ), .ZN(\dp/ex_stage/alu/r60/n97 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U134  ( .B1(\dp/ex_stage/alu/r60/n172 ), .B2(
        \dp/ex_stage/alu/r60/n97 ), .A(\dp/ex_stage/alu/r60/n173 ), .ZN(
        \dp/ex_stage/alu/r60/n171 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U133  ( .A1(\dp/ex_stage/alu/r60/n8 ), .A2(
        \dp/ex_stage/muxB_out [21]), .ZN(\dp/ex_stage/alu/r60/n93 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U132  ( .A1(\dp/ex_stage/muxB_out [21]), .A2(
        \dp/ex_stage/alu/r60/n8 ), .ZN(\dp/ex_stage/alu/r60/n152 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U131  ( .B1(\dp/ex_stage/alu/r60/n171 ), .B2(
        \dp/ex_stage/alu/r60/n48 ), .A(\dp/ex_stage/alu/r60/n152 ), .ZN(
        \dp/ex_stage/alu/r60/n169 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U130  ( .A1(\dp/ex_stage/alu/r60/n9 ), .A2(
        \dp/ex_stage/muxB_out [22]), .ZN(\dp/ex_stage/alu/r60/n170 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U129  ( .A1(\dp/ex_stage/muxB_out [22]), .A2(
        \dp/ex_stage/alu/r60/n9 ), .ZN(\dp/ex_stage/alu/r60/n89 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U128  ( .A1(\dp/ex_stage/alu/r60/n50 ), .A2(
        \dp/ex_stage/alu/r60/n89 ), .ZN(\dp/ex_stage/alu/r60/n92 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U127  ( .B1(\dp/ex_stage/alu/r60/n169 ), .B2(
        \dp/ex_stage/alu/r60/n49 ), .A(\dp/ex_stage/alu/r60/n170 ), .ZN(
        \dp/ex_stage/alu/r60/n168 ) );
  OR2_X1 \dp/ex_stage/alu/r60/U126  ( .A1(\dp/ex_stage/alu/r60/n10 ), .A2(
        \dp/ex_stage/muxB_out [23]), .ZN(\dp/ex_stage/alu/r60/n86 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U125  ( .A1(\dp/ex_stage/muxB_out [23]), .A2(
        \dp/ex_stage/alu/r60/n10 ), .ZN(\dp/ex_stage/alu/r60/n88 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U124  ( .B1(\dp/ex_stage/alu/r60/n168 ), .B2(
        \dp/ex_stage/alu/r60/n86 ), .A(\dp/ex_stage/alu/r60/n51 ), .ZN(
        \dp/ex_stage/alu/r60/n166 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U123  ( .A1(\dp/ex_stage/alu/r60/n52 ), .A2(
        \dp/ex_stage/muxB_out [24]), .ZN(\dp/ex_stage/alu/r60/n167 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U122  ( .A1(\dp/ex_stage/muxB_out [24]), .A2(
        \dp/ex_stage/alu/r60/n52 ), .ZN(\dp/ex_stage/alu/r60/n153 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U121  ( .A1(\dp/ex_stage/alu/r60/n167 ), .A2(
        \dp/ex_stage/alu/r60/n153 ), .ZN(\dp/ex_stage/alu/r60/n87 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U120  ( .B1(\dp/ex_stage/alu/r60/n166 ), .B2(
        \dp/ex_stage/alu/r60/n87 ), .A(\dp/ex_stage/alu/r60/n167 ), .ZN(
        \dp/ex_stage/alu/r60/n165 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U119  ( .A1(\dp/ex_stage/alu/r60/n54 ), .A2(
        \dp/ex_stage/muxB_out [25]), .ZN(\dp/ex_stage/alu/r60/n83 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U118  ( .A1(\dp/ex_stage/muxB_out [25]), .A2(
        \dp/ex_stage/alu/r60/n54 ), .ZN(\dp/ex_stage/alu/r60/n154 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U117  ( .B1(\dp/ex_stage/alu/r60/n165 ), .B2(
        \dp/ex_stage/alu/r60/n53 ), .A(\dp/ex_stage/alu/r60/n154 ), .ZN(
        \dp/ex_stage/alu/r60/n163 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U116  ( .A1(\dp/ex_stage/alu/r60/n57 ), .A2(
        \dp/ex_stage/muxB_out [26]), .ZN(\dp/ex_stage/alu/r60/n164 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U115  ( .A1(\dp/ex_stage/muxB_out [26]), .A2(
        \dp/ex_stage/alu/r60/n57 ), .ZN(\dp/ex_stage/alu/r60/n79 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U114  ( .A1(\dp/ex_stage/alu/r60/n56 ), .A2(
        \dp/ex_stage/alu/r60/n79 ), .ZN(\dp/ex_stage/alu/r60/n82 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U113  ( .B1(\dp/ex_stage/alu/r60/n163 ), .B2(
        \dp/ex_stage/alu/r60/n55 ), .A(\dp/ex_stage/alu/r60/n164 ), .ZN(
        \dp/ex_stage/alu/r60/n162 ) );
  OR2_X1 \dp/ex_stage/alu/r60/U112  ( .A1(\dp/ex_stage/alu/r60/n59 ), .A2(
        \dp/ex_stage/muxB_out [27]), .ZN(\dp/ex_stage/alu/r60/n76 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U111  ( .A1(\dp/ex_stage/muxB_out [27]), .A2(
        \dp/ex_stage/alu/r60/n59 ), .ZN(\dp/ex_stage/alu/r60/n78 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U110  ( .B1(\dp/ex_stage/alu/r60/n162 ), .B2(
        \dp/ex_stage/alu/r60/n76 ), .A(\dp/ex_stage/alu/r60/n58 ), .ZN(
        \dp/ex_stage/alu/r60/n160 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U109  ( .A1(\dp/ex_stage/alu/r60/n60 ), .A2(
        \dp/ex_stage/muxB_out [28]), .ZN(\dp/ex_stage/alu/r60/n161 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U108  ( .A1(\dp/ex_stage/muxB_out [28]), .A2(
        \dp/ex_stage/alu/r60/n60 ), .ZN(\dp/ex_stage/alu/r60/n155 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U107  ( .A1(\dp/ex_stage/alu/r60/n161 ), .A2(
        \dp/ex_stage/alu/r60/n155 ), .ZN(\dp/ex_stage/alu/r60/n77 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U106  ( .B1(\dp/ex_stage/alu/r60/n160 ), .B2(
        \dp/ex_stage/alu/r60/n77 ), .A(\dp/ex_stage/alu/r60/n161 ), .ZN(
        \dp/ex_stage/alu/r60/n159 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U105  ( .A1(\dp/ex_stage/alu/r60/n62 ), .A2(
        \dp/ex_stage/muxB_out [29]), .ZN(\dp/ex_stage/alu/r60/n73 ) );
  AND2_X1 \dp/ex_stage/alu/r60/U104  ( .A1(\dp/ex_stage/muxB_out [29]), .A2(
        \dp/ex_stage/alu/r60/n62 ), .ZN(\dp/ex_stage/alu/r60/n156 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U103  ( .B1(\dp/ex_stage/alu/r60/n159 ), .B2(
        \dp/ex_stage/alu/r60/n61 ), .A(\dp/ex_stage/alu/r60/n156 ), .ZN(
        \dp/ex_stage/alu/r60/n158 ) );
  XOR2_X1 \dp/ex_stage/alu/r60/U102  ( .A(\dp/ex_stage/alu/r60/n65 ), .B(
        \dp/ex_stage/muxA_out [30]), .Z(\dp/ex_stage/alu/r60/n70 ) );
  AOI22_X1 \dp/ex_stage/alu/r60/U101  ( .A1(\dp/ex_stage/muxA_out [30]), .A2(
        \dp/ex_stage/alu/r60/n65 ), .B1(\dp/ex_stage/alu/r60/n158 ), .B2(
        \dp/ex_stage/alu/r60/n70 ), .ZN(\dp/ex_stage/alu/r60/n157 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U100  ( .A1(\dp/ex_stage/muxB_out [31]), .A2(
        \dp/ex_stage/alu/r60/n64 ), .ZN(\dp/ex_stage/alu/r60/n66 ) );
  OAI21_X1 \dp/ex_stage/alu/r60/U99  ( .B1(\dp/ex_stage/alu/r60/n67 ), .B2(
        \dp/ex_stage/alu/r60/n157 ), .A(\dp/ex_stage/alu/r60/n66 ), .ZN(
        \dp/ex_stage/alu/N20 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U98  ( .A1(\dp/ex_stage/alu/r60/n155 ), .A2(
        \dp/ex_stage/alu/r60/n156 ), .ZN(\dp/ex_stage/alu/r60/n71 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U97  ( .A1(\dp/ex_stage/alu/r60/n153 ), .A2(
        \dp/ex_stage/alu/r60/n154 ), .ZN(\dp/ex_stage/alu/r60/n80 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U96  ( .A1(\dp/ex_stage/alu/r60/n151 ), .A2(
        \dp/ex_stage/alu/r60/n152 ), .ZN(\dp/ex_stage/alu/r60/n90 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U95  ( .A1(\dp/ex_stage/alu/r60/n149 ), .A2(
        \dp/ex_stage/alu/r60/n150 ), .ZN(\dp/ex_stage/alu/r60/n100 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U94  ( .A1(\dp/ex_stage/alu/r60/n147 ), .A2(
        \dp/ex_stage/alu/r60/n148 ), .ZN(\dp/ex_stage/alu/r60/n110 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U93  ( .A1(\dp/ex_stage/alu/r60/n145 ), .A2(
        \dp/ex_stage/alu/r60/n146 ), .ZN(\dp/ex_stage/alu/r60/n120 ) );
  NOR2_X1 \dp/ex_stage/alu/r60/U92  ( .A1(\dp/ex_stage/alu/r60/n143 ), .A2(
        \dp/ex_stage/alu/r60/n144 ), .ZN(\dp/ex_stage/alu/r60/n130 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U91  ( .A1(\dp/ex_stage/muxB_out [0]), .A2(
        \dp/ex_stage/alu/r60/n16 ), .ZN(\dp/ex_stage/alu/r60/n142 ) );
  OAI21_X1 \dp/ex_stage/alu/r60/U90  ( .B1(\dp/ex_stage/alu/r60/n1 ), .B2(
        \dp/ex_stage/alu/r60/n142 ), .A(\dp/ex_stage/muxA_out [1]), .ZN(
        \dp/ex_stage/alu/r60/n140 ) );
  OAI211_X1 \dp/ex_stage/alu/r60/U89  ( .C1(\dp/ex_stage/alu/n25 ), .C2(
        \dp/ex_stage/alu/r60/n15 ), .A(\dp/ex_stage/alu/r60/n140 ), .B(
        \dp/ex_stage/alu/r60/n141 ), .ZN(\dp/ex_stage/alu/r60/n139 ) );
  NAND3_X1 \dp/ex_stage/alu/r60/U88  ( .A1(\dp/ex_stage/alu/r60/n137 ), .A2(
        \dp/ex_stage/alu/r60/n138 ), .A3(\dp/ex_stage/alu/r60/n139 ), .ZN(
        \dp/ex_stage/alu/r60/n134 ) );
  NAND3_X1 \dp/ex_stage/alu/r60/U87  ( .A1(\dp/ex_stage/alu/r60/n134 ), .A2(
        \dp/ex_stage/alu/r60/n135 ), .A3(\dp/ex_stage/alu/r60/n136 ), .ZN(
        \dp/ex_stage/alu/r60/n131 ) );
  AOI211_X1 \dp/ex_stage/alu/r60/U86  ( .C1(\dp/ex_stage/alu/r60/n130 ), .C2(
        \dp/ex_stage/alu/r60/n131 ), .A(\dp/ex_stage/alu/r60/n132 ), .B(
        \dp/ex_stage/alu/r60/n133 ), .ZN(\dp/ex_stage/alu/r60/n124 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U85  ( .A1(\dp/ex_stage/alu/r60/n128 ), .A2(
        \dp/ex_stage/alu/r60/n129 ), .ZN(\dp/ex_stage/alu/r60/n125 ) );
  OAI211_X1 \dp/ex_stage/alu/r60/U84  ( .C1(\dp/ex_stage/alu/r60/n124 ), .C2(
        \dp/ex_stage/alu/r60/n125 ), .A(\dp/ex_stage/alu/r60/n126 ), .B(
        \dp/ex_stage/alu/r60/n127 ), .ZN(\dp/ex_stage/alu/r60/n121 ) );
  AOI211_X1 \dp/ex_stage/alu/r60/U83  ( .C1(\dp/ex_stage/alu/r60/n120 ), .C2(
        \dp/ex_stage/alu/r60/n121 ), .A(\dp/ex_stage/alu/r60/n122 ), .B(
        \dp/ex_stage/alu/r60/n123 ), .ZN(\dp/ex_stage/alu/r60/n114 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U82  ( .A1(\dp/ex_stage/alu/r60/n118 ), .A2(
        \dp/ex_stage/alu/r60/n119 ), .ZN(\dp/ex_stage/alu/r60/n115 ) );
  OAI211_X1 \dp/ex_stage/alu/r60/U81  ( .C1(\dp/ex_stage/alu/r60/n114 ), .C2(
        \dp/ex_stage/alu/r60/n115 ), .A(\dp/ex_stage/alu/r60/n116 ), .B(
        \dp/ex_stage/alu/r60/n117 ), .ZN(\dp/ex_stage/alu/r60/n111 ) );
  AOI211_X1 \dp/ex_stage/alu/r60/U80  ( .C1(\dp/ex_stage/alu/r60/n110 ), .C2(
        \dp/ex_stage/alu/r60/n111 ), .A(\dp/ex_stage/alu/r60/n112 ), .B(
        \dp/ex_stage/alu/r60/n113 ), .ZN(\dp/ex_stage/alu/r60/n104 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U79  ( .A1(\dp/ex_stage/alu/r60/n108 ), .A2(
        \dp/ex_stage/alu/r60/n109 ), .ZN(\dp/ex_stage/alu/r60/n105 ) );
  OAI211_X1 \dp/ex_stage/alu/r60/U78  ( .C1(\dp/ex_stage/alu/r60/n104 ), .C2(
        \dp/ex_stage/alu/r60/n105 ), .A(\dp/ex_stage/alu/r60/n106 ), .B(
        \dp/ex_stage/alu/r60/n107 ), .ZN(\dp/ex_stage/alu/r60/n101 ) );
  AOI211_X1 \dp/ex_stage/alu/r60/U77  ( .C1(\dp/ex_stage/alu/r60/n100 ), .C2(
        \dp/ex_stage/alu/r60/n101 ), .A(\dp/ex_stage/alu/r60/n102 ), .B(
        \dp/ex_stage/alu/r60/n103 ), .ZN(\dp/ex_stage/alu/r60/n94 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U76  ( .A1(\dp/ex_stage/alu/r60/n98 ), .A2(
        \dp/ex_stage/alu/r60/n99 ), .ZN(\dp/ex_stage/alu/r60/n95 ) );
  OAI211_X1 \dp/ex_stage/alu/r60/U75  ( .C1(\dp/ex_stage/alu/r60/n94 ), .C2(
        \dp/ex_stage/alu/r60/n95 ), .A(\dp/ex_stage/alu/r60/n96 ), .B(
        \dp/ex_stage/alu/r60/n97 ), .ZN(\dp/ex_stage/alu/r60/n91 ) );
  AOI211_X1 \dp/ex_stage/alu/r60/U74  ( .C1(\dp/ex_stage/alu/r60/n90 ), .C2(
        \dp/ex_stage/alu/r60/n91 ), .A(\dp/ex_stage/alu/r60/n92 ), .B(
        \dp/ex_stage/alu/r60/n93 ), .ZN(\dp/ex_stage/alu/r60/n84 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U73  ( .A1(\dp/ex_stage/alu/r60/n88 ), .A2(
        \dp/ex_stage/alu/r60/n89 ), .ZN(\dp/ex_stage/alu/r60/n85 ) );
  OAI211_X1 \dp/ex_stage/alu/r60/U72  ( .C1(\dp/ex_stage/alu/r60/n84 ), .C2(
        \dp/ex_stage/alu/r60/n85 ), .A(\dp/ex_stage/alu/r60/n86 ), .B(
        \dp/ex_stage/alu/r60/n87 ), .ZN(\dp/ex_stage/alu/r60/n81 ) );
  AOI211_X1 \dp/ex_stage/alu/r60/U71  ( .C1(\dp/ex_stage/alu/r60/n80 ), .C2(
        \dp/ex_stage/alu/r60/n81 ), .A(\dp/ex_stage/alu/r60/n82 ), .B(
        \dp/ex_stage/alu/r60/n83 ), .ZN(\dp/ex_stage/alu/r60/n74 ) );
  NAND2_X1 \dp/ex_stage/alu/r60/U70  ( .A1(\dp/ex_stage/alu/r60/n78 ), .A2(
        \dp/ex_stage/alu/r60/n79 ), .ZN(\dp/ex_stage/alu/r60/n75 ) );
  OAI211_X1 \dp/ex_stage/alu/r60/U69  ( .C1(\dp/ex_stage/alu/r60/n74 ), .C2(
        \dp/ex_stage/alu/r60/n75 ), .A(\dp/ex_stage/alu/r60/n76 ), .B(
        \dp/ex_stage/alu/r60/n77 ), .ZN(\dp/ex_stage/alu/r60/n72 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U68  ( .B1(\dp/ex_stage/alu/r60/n71 ), .B2(
        \dp/ex_stage/alu/r60/n72 ), .A(\dp/ex_stage/alu/r60/n73 ), .ZN(
        \dp/ex_stage/alu/r60/n69 ) );
  AOI22_X1 \dp/ex_stage/alu/r60/U67  ( .A1(\dp/ex_stage/muxB_out [30]), .A2(
        \dp/ex_stage/alu/r60/n63 ), .B1(\dp/ex_stage/alu/r60/n69 ), .B2(
        \dp/ex_stage/alu/r60/n70 ), .ZN(\dp/ex_stage/alu/r60/n68 ) );
  AOI21_X1 \dp/ex_stage/alu/r60/U66  ( .B1(\dp/ex_stage/alu/r60/n66 ), .B2(
        \dp/ex_stage/alu/r60/n14 ), .A(\dp/ex_stage/alu/r60/n67 ), .ZN(
        \dp/ex_stage/alu/N16 ) );
  INV_X1 \dp/ex_stage/alu/r60/U65  ( .A(\dp/ex_stage/alu/n45 ), .ZN(
        \dp/ex_stage/alu/r60/n10 ) );
  INV_X1 \dp/ex_stage/alu/r60/U64  ( .A(\dp/ex_stage/alu/n43 ), .ZN(
        \dp/ex_stage/alu/r60/n9 ) );
  INV_X1 \dp/ex_stage/alu/r60/U63  ( .A(\dp/ex_stage/muxA_out [21]), .ZN(
        \dp/ex_stage/alu/r60/n8 ) );
  INV_X1 \dp/ex_stage/alu/r60/U62  ( .A(\dp/ex_stage/muxA_out [17]), .ZN(
        \dp/ex_stage/alu/r60/n7 ) );
  INV_X1 \dp/ex_stage/alu/r60/U61  ( .A(\dp/ex_stage/muxA_out [16]), .ZN(
        \dp/ex_stage/alu/r60/n6 ) );
  INV_X1 \dp/ex_stage/alu/r60/U60  ( .A(\dp/ex_stage/muxA_out [15]), .ZN(
        \dp/ex_stage/alu/r60/n5 ) );
  INV_X1 \dp/ex_stage/alu/r60/U59  ( .A(\dp/ex_stage/alu/n37 ), .ZN(
        \dp/ex_stage/alu/r60/n4 ) );
  INV_X1 \dp/ex_stage/alu/r60/U58  ( .A(\dp/ex_stage/muxA_out [13]), .ZN(
        \dp/ex_stage/alu/r60/n3 ) );
  INV_X1 \dp/ex_stage/alu/r60/U57  ( .A(\dp/ex_stage/alu/n34 ), .ZN(
        \dp/ex_stage/alu/r60/n2 ) );
  INV_X1 \dp/ex_stage/alu/r60/U56  ( .A(\dp/ex_stage/alu/n25 ), .ZN(
        \dp/ex_stage/alu/r60/n1 ) );
  INV_X1 \dp/ex_stage/alu/r60/U55  ( .A(\dp/ex_stage/alu/N16 ), .ZN(
        \dp/ex_stage/alu/N22 ) );
  INV_X1 \dp/ex_stage/alu/r60/U54  ( .A(\dp/ex_stage/alu/N20 ), .ZN(
        \dp/ex_stage/alu/N17 ) );
  INV_X1 \dp/ex_stage/alu/r60/U53  ( .A(\dp/ex_stage/muxB_out [30]), .ZN(
        \dp/ex_stage/alu/r60/n65 ) );
  INV_X1 \dp/ex_stage/alu/r60/U52  ( .A(\dp/ex_stage/muxA_out [19]), .ZN(
        \dp/ex_stage/alu/r60/n46 ) );
  INV_X1 \dp/ex_stage/alu/r60/U51  ( .A(\dp/ex_stage/muxA_out [20]), .ZN(
        \dp/ex_stage/alu/r60/n47 ) );
  INV_X1 \dp/ex_stage/alu/r60/U50  ( .A(\dp/ex_stage/muxA_out [29]), .ZN(
        \dp/ex_stage/alu/r60/n62 ) );
  INV_X1 \dp/ex_stage/alu/r60/U49  ( .A(\dp/ex_stage/alu/shifter/N136 ), .ZN(
        \dp/ex_stage/alu/r60/n64 ) );
  INV_X1 \dp/ex_stage/alu/r60/U48  ( .A(\dp/ex_stage/muxA_out [27]), .ZN(
        \dp/ex_stage/alu/r60/n59 ) );
  INV_X1 \dp/ex_stage/alu/r60/U47  ( .A(\dp/ex_stage/muxA_out [28]), .ZN(
        \dp/ex_stage/alu/r60/n60 ) );
  INV_X1 \dp/ex_stage/alu/r60/U46  ( .A(\dp/ex_stage/muxA_out [25]), .ZN(
        \dp/ex_stage/alu/r60/n54 ) );
  INV_X1 \dp/ex_stage/alu/r60/U45  ( .A(\dp/ex_stage/muxA_out [24]), .ZN(
        \dp/ex_stage/alu/r60/n52 ) );
  INV_X1 \dp/ex_stage/alu/r60/U44  ( .A(\dp/ex_stage/muxA_out [18]), .ZN(
        \dp/ex_stage/alu/r60/n44 ) );
  INV_X1 \dp/ex_stage/alu/r60/U43  ( .A(\dp/ex_stage/muxA_out [26]), .ZN(
        \dp/ex_stage/alu/r60/n57 ) );
  INV_X1 \dp/ex_stage/alu/r60/U42  ( .A(\dp/ex_stage/muxA_out [30]), .ZN(
        \dp/ex_stage/alu/r60/n63 ) );
  INV_X1 \dp/ex_stage/alu/r60/U41  ( .A(\dp/ex_stage/alu/r60/n68 ), .ZN(
        \dp/ex_stage/alu/r60/n14 ) );
  INV_X1 \dp/ex_stage/alu/r60/U40  ( .A(\dp/ex_stage/alu/r60/n200 ), .ZN(
        \dp/ex_stage/alu/r60/n12 ) );
  INV_X1 \dp/ex_stage/alu/r60/U39  ( .A(\dp/ex_stage/muxA_out [5]), .ZN(
        \dp/ex_stage/alu/r60/n23 ) );
  INV_X1 \dp/ex_stage/alu/r60/U38  ( .A(\dp/ex_stage/muxA_out [4]), .ZN(
        \dp/ex_stage/alu/r60/n21 ) );
  INV_X1 \dp/ex_stage/alu/r60/U37  ( .A(\dp/ex_stage/muxA_out [6]), .ZN(
        \dp/ex_stage/alu/r60/n26 ) );
  INV_X1 \dp/ex_stage/alu/r60/U36  ( .A(\dp/ex_stage/muxA_out [3]), .ZN(
        \dp/ex_stage/alu/r60/n20 ) );
  INV_X1 \dp/ex_stage/alu/r60/U35  ( .A(\dp/ex_stage/muxA_out [11]), .ZN(
        \dp/ex_stage/alu/r60/n36 ) );
  INV_X1 \dp/ex_stage/alu/r60/U34  ( .A(\dp/ex_stage/muxA_out [7]), .ZN(
        \dp/ex_stage/alu/r60/n28 ) );
  INV_X1 \dp/ex_stage/alu/r60/U33  ( .A(\dp/ex_stage/muxA_out [9]), .ZN(
        \dp/ex_stage/alu/r60/n31 ) );
  INV_X1 \dp/ex_stage/alu/r60/U32  ( .A(\dp/ex_stage/muxA_out [8]), .ZN(
        \dp/ex_stage/alu/r60/n29 ) );
  INV_X1 \dp/ex_stage/alu/r60/U31  ( .A(\dp/ex_stage/alu/shifter/N202 ), .ZN(
        \dp/ex_stage/alu/r60/n16 ) );
  INV_X1 \dp/ex_stage/alu/r60/U30  ( .A(\dp/ex_stage/muxA_out [2]), .ZN(
        \dp/ex_stage/alu/r60/n18 ) );
  INV_X1 \dp/ex_stage/alu/r60/U29  ( .A(\dp/ex_stage/muxA_out [10]), .ZN(
        \dp/ex_stage/alu/r60/n34 ) );
  INV_X1 \dp/ex_stage/alu/r60/U28  ( .A(\dp/ex_stage/alu/r60/n142 ), .ZN(
        \dp/ex_stage/alu/r60/n15 ) );
  INV_X1 \dp/ex_stage/alu/r60/U27  ( .A(\dp/ex_stage/alu/r60/n73 ), .ZN(
        \dp/ex_stage/alu/r60/n61 ) );
  INV_X1 \dp/ex_stage/alu/r60/U26  ( .A(\dp/ex_stage/alu/r60/n88 ), .ZN(
        \dp/ex_stage/alu/r60/n51 ) );
  INV_X1 \dp/ex_stage/alu/r60/U25  ( .A(\dp/ex_stage/alu/r60/n108 ), .ZN(
        \dp/ex_stage/alu/r60/n40 ) );
  INV_X1 \dp/ex_stage/alu/r60/U24  ( .A(\dp/ex_stage/alu/r60/n164 ), .ZN(
        \dp/ex_stage/alu/r60/n56 ) );
  INV_X1 \dp/ex_stage/alu/r60/U23  ( .A(\dp/ex_stage/alu/r60/n170 ), .ZN(
        \dp/ex_stage/alu/r60/n50 ) );
  INV_X1 \dp/ex_stage/alu/r60/U22  ( .A(\dp/ex_stage/alu/r60/n176 ), .ZN(
        \dp/ex_stage/alu/r60/n43 ) );
  INV_X1 \dp/ex_stage/alu/r60/U21  ( .A(\dp/ex_stage/alu/r60/n128 ), .ZN(
        \dp/ex_stage/alu/r60/n27 ) );
  INV_X1 \dp/ex_stage/alu/r60/U20  ( .A(\dp/ex_stage/alu/r60/n182 ), .ZN(
        \dp/ex_stage/alu/r60/n39 ) );
  INV_X1 \dp/ex_stage/alu/r60/U19  ( .A(\dp/ex_stage/alu/r60/n188 ), .ZN(
        \dp/ex_stage/alu/r60/n33 ) );
  INV_X1 \dp/ex_stage/alu/r60/U18  ( .A(\dp/ex_stage/alu/r60/n194 ), .ZN(
        \dp/ex_stage/alu/r60/n25 ) );
  INV_X1 \dp/ex_stage/alu/r60/U17  ( .A(\dp/ex_stage/alu/r60/n83 ), .ZN(
        \dp/ex_stage/alu/r60/n53 ) );
  INV_X1 \dp/ex_stage/alu/r60/U16  ( .A(\dp/ex_stage/alu/r60/n98 ), .ZN(
        \dp/ex_stage/alu/r60/n45 ) );
  INV_X1 \dp/ex_stage/alu/r60/U15  ( .A(\dp/ex_stage/alu/r60/n103 ), .ZN(
        \dp/ex_stage/alu/r60/n41 ) );
  INV_X1 \dp/ex_stage/alu/r60/U14  ( .A(\dp/ex_stage/alu/r60/n137 ), .ZN(
        \dp/ex_stage/alu/r60/n19 ) );
  INV_X1 \dp/ex_stage/alu/r60/U13  ( .A(\dp/ex_stage/alu/r60/n113 ), .ZN(
        \dp/ex_stage/alu/r60/n37 ) );
  INV_X1 \dp/ex_stage/alu/r60/U12  ( .A(\dp/ex_stage/alu/r60/n112 ), .ZN(
        \dp/ex_stage/alu/r60/n38 ) );
  INV_X1 \dp/ex_stage/alu/r60/U11  ( .A(\dp/ex_stage/alu/r60/n118 ), .ZN(
        \dp/ex_stage/alu/r60/n35 ) );
  INV_X1 \dp/ex_stage/alu/r60/U10  ( .A(\dp/ex_stage/alu/r60/n123 ), .ZN(
        \dp/ex_stage/alu/r60/n30 ) );
  INV_X1 \dp/ex_stage/alu/r60/U9  ( .A(\dp/ex_stage/alu/r60/n78 ), .ZN(
        \dp/ex_stage/alu/r60/n58 ) );
  INV_X1 \dp/ex_stage/alu/r60/U8  ( .A(\dp/ex_stage/alu/r60/n93 ), .ZN(
        \dp/ex_stage/alu/r60/n48 ) );
  INV_X1 \dp/ex_stage/alu/r60/U7  ( .A(\dp/ex_stage/alu/r60/n92 ), .ZN(
        \dp/ex_stage/alu/r60/n49 ) );
  INV_X1 \dp/ex_stage/alu/r60/U6  ( .A(\dp/ex_stage/alu/r60/n133 ), .ZN(
        \dp/ex_stage/alu/r60/n22 ) );
  INV_X1 \dp/ex_stage/alu/r60/U5  ( .A(\dp/ex_stage/alu/r60/n132 ), .ZN(
        \dp/ex_stage/alu/r60/n24 ) );
  INV_X1 \dp/ex_stage/alu/r60/U4  ( .A(\dp/ex_stage/alu/r60/n82 ), .ZN(
        \dp/ex_stage/alu/r60/n55 ) );
  INV_X1 \dp/ex_stage/alu/r60/U3  ( .A(\dp/ex_stage/alu/r60/n102 ), .ZN(
        \dp/ex_stage/alu/r60/n42 ) );
  INV_X1 \dp/ex_stage/alu/r60/U2  ( .A(\dp/ex_stage/alu/r60/n122 ), .ZN(
        \dp/ex_stage/alu/r60/n32 ) );
  INV_X1 \dp/ex_stage/alu/r60/U1  ( .A(\dp/ex_stage/alu/r60/n138 ), .ZN(
        \dp/ex_stage/alu/r60/n17 ) );
endmodule

