
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX.all;

entity DLX is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ISSUE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ISSUE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA : inout 
         std_logic_vector (31 downto 0));

end DLX;

architecture SYN_dlx_rtl of DLX is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X2
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component TBUF_X1
      port( A, EN : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X4
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ISSUE_port, DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, DRAM_ADDRESS_0_port, 
      DRAM_ISSUE_port, DRAM_READNOTWRITE_port, pipe_if_id_en_i, 
      pipe_ex_mem_en_i, pipe_clear_n_i, rf_call_i, rf_ret_i, rf_spill_i, 
      rf_fill_i, rf_en_i, rf_rs1_en_i, rf_rs2_en_i, imm_isoff_i, imm_uns_i, 
      reg31_sel_i, regrd_sel_i, muxA_sel_i, muxB_sel_i, is_zero_i, 
      alu_op_i_4_port, alu_op_i_3_port, alu_op_i_2_port, alu_op_i_1_port, 
      alu_op_i_0_port, mem_in_en_i, npc_wb_en_i, jump_en_i, wb_mux_sel_i, 
      rf_we_i, CU_I_n291, CU_I_n290, CU_I_n289, CU_I_n288, CU_I_n287, CU_I_n286
      , CU_I_n285, CU_I_n284, CU_I_n283, CU_I_n282, CU_I_n281, CU_I_n280, 
      CU_I_n279, CU_I_n278, CU_I_n277, CU_I_n276, CU_I_n275, CU_I_n274, 
      CU_I_n273, CU_I_n272, CU_I_n271, CU_I_n270, CU_I_n269, CU_I_n268, 
      CU_I_n267, CU_I_n266, CU_I_n265, CU_I_n264, CU_I_n263, CU_I_n262, 
      CU_I_n261, CU_I_n260, CU_I_n259, CU_I_n258, CU_I_n257, CU_I_n256, 
      CU_I_n76, CU_I_n75, CU_I_n74, CU_I_n73, CU_I_n72, CU_I_n71, CU_I_n70, 
      CU_I_n69, CU_I_n68, CU_I_n67, CU_I_n66, CU_I_n65, CU_I_n64, CU_I_n63, 
      CU_I_n60, CU_I_n59, CU_I_n58, CU_I_n57, CU_I_n56, CU_I_n55, CU_I_n54, 
      CU_I_n53, CU_I_n52, CU_I_n51, CU_I_n50, CU_I_n49, CU_I_n48, CU_I_n47, 
      CU_I_n45, CU_I_n43, CU_I_n42, CU_I_n41, CU_I_n39, CU_I_n38, CU_I_n29, 
      CU_I_n28, CU_I_n26, CU_I_n25, CU_I_n24, CU_I_n20, CU_I_n18, CU_I_n14, 
      CU_I_n1, CU_I_n254, CU_I_n253, CU_I_n252, CU_I_n251, CU_I_n250, CU_I_n249
      , CU_I_n248, CU_I_n247, CU_I_n246, CU_I_n245, CU_I_n244, CU_I_n243, 
      CU_I_n242, CU_I_n241, CU_I_n240, CU_I_n239, CU_I_n238, CU_I_n237, 
      CU_I_n236, CU_I_n235, CU_I_n234, CU_I_n233, CU_I_n232, CU_I_n231, 
      CU_I_n230, CU_I_n229, CU_I_n228, CU_I_n227, CU_I_n226, CU_I_n225, 
      CU_I_n224, CU_I_n223, CU_I_n222, CU_I_n221, CU_I_n220, CU_I_n219, 
      CU_I_n218, CU_I_n217, CU_I_n216, CU_I_n215, CU_I_n214, CU_I_n213, 
      CU_I_n212, CU_I_n211, CU_I_n210, CU_I_n209, CU_I_n208, CU_I_n207, 
      CU_I_n206, CU_I_n205, CU_I_n204, CU_I_n203, CU_I_n202, CU_I_n201, 
      CU_I_n200, CU_I_n199, CU_I_n198, CU_I_n197, CU_I_n196, CU_I_n195, 
      CU_I_n194, CU_I_n193, CU_I_n192, CU_I_n191, CU_I_n190, CU_I_n189, 
      CU_I_n188, CU_I_n187, CU_I_n186, CU_I_n185, CU_I_n184, CU_I_n183, 
      CU_I_n182, CU_I_n181, CU_I_n180, CU_I_n179, CU_I_n178, CU_I_n177, 
      CU_I_n176, CU_I_n175, CU_I_n174, CU_I_n173, CU_I_n172, CU_I_n171, 
      CU_I_n170, CU_I_n169, CU_I_n168, CU_I_n167, CU_I_n166, CU_I_n165, 
      CU_I_n164, CU_I_n163, CU_I_n162, CU_I_n161, CU_I_n160, CU_I_n159, 
      CU_I_n158, CU_I_n157, CU_I_n156, CU_I_n155, CU_I_n154, CU_I_n153, 
      CU_I_n152, CU_I_n151, CU_I_n150, CU_I_n149, CU_I_n148, CU_I_n147, 
      CU_I_n146, CU_I_n145, CU_I_n144, CU_I_n143, CU_I_n142, CU_I_n141, 
      CU_I_n140, CU_I_n139, CU_I_n138, CU_I_n137, CU_I_n136, CU_I_n135, 
      CU_I_n134, CU_I_n133, CU_I_n132, CU_I_n131, CU_I_n130, CU_I_n129, 
      CU_I_n128, CU_I_n127, CU_I_n126, CU_I_n125, CU_I_n124, CU_I_n123, 
      CU_I_n122, CU_I_n121, CU_I_n120, CU_I_n119, CU_I_n118, CU_I_n117, 
      CU_I_n116, CU_I_n115, CU_I_n114, CU_I_n113, CU_I_n112, CU_I_n111, 
      CU_I_n110, CU_I_n109, CU_I_n108, CU_I_n107, CU_I_n106, CU_I_n105, 
      CU_I_n104, CU_I_n103, CU_I_n102, CU_I_n101, CU_I_n100, CU_I_n99, CU_I_n98
      , CU_I_n97, CU_I_n96, CU_I_n95, CU_I_n94, CU_I_n93, CU_I_n92, CU_I_n91, 
      CU_I_n90, CU_I_n89, CU_I_n88, CU_I_n87, CU_I_n86, CU_I_n85, CU_I_n84, 
      CU_I_n83, CU_I_n82, CU_I_n81, CU_I_n80, CU_I_n79, CU_I_n78, CU_I_n77, 
      CU_I_n37, CU_I_n36, CU_I_n35, CU_I_n34, CU_I_n33, CU_I_n32, CU_I_n31, 
      CU_I_n30, CU_I_n27, CU_I_n23, CU_I_n22, CU_I_n21, CU_I_n19, CU_I_n17, 
      CU_I_n16, CU_I_n15, CU_I_n13, CU_I_n12, CU_I_n11, CU_I_n10, CU_I_n9, 
      CU_I_n8, CU_I_n7, CU_I_n6, CU_I_n5, CU_I_n4, CU_I_n3, CU_I_n2, 
      CU_I_cw3_4_port, CU_I_cw3_5_port, CU_I_cw2_4_port, CU_I_cw2_5_port, 
      CU_I_cw1_1_port, CU_I_n294, CU_I_n293, CU_I_n292, CU_I_Logic0_port, 
      CU_I_Logic1_port, dp_n1055, dp_n1054, dp_n1053, dp_n1052, dp_n1051, 
      dp_n1050, dp_n1049, dp_n1048, dp_n1047, dp_n1046, dp_n1045, dp_n1044, 
      dp_n1043, dp_n1042, dp_n1041, dp_n1040, dp_n1039, dp_n1038, dp_n1037, 
      dp_n1036, dp_n1035, dp_n1034, dp_n1033, dp_n1032, dp_n1031, dp_n1030, 
      dp_n1029, dp_n1028, dp_n1027, dp_n1026, dp_n1025, dp_n1024, dp_n1023, 
      dp_n1022, dp_n1021, dp_n1020, dp_n1019, dp_n1018, dp_n1017, dp_n1016, 
      dp_n648, dp_n647, dp_n646, dp_n645, dp_n644, dp_n643, dp_n642, dp_n641, 
      dp_n640, dp_n639, dp_n638, dp_n637, dp_n636, dp_n635, dp_n634, dp_n633, 
      dp_n632, dp_n631, dp_n630, dp_n629, dp_n628, dp_n627, dp_n626, dp_n625, 
      dp_n624, dp_n623, dp_n622, dp_n621, dp_n620, dp_n619, dp_n618, dp_n617, 
      dp_n616, dp_n615, dp_n614, dp_n613, dp_n612, dp_n611, dp_n610, dp_n609, 
      dp_n608, dp_n607, dp_n606, dp_n605, dp_n604, dp_n603, dp_n602, dp_n601, 
      dp_n600, dp_n599, dp_n598, dp_n597, dp_n596, dp_n595, dp_n594, dp_n593, 
      dp_n592, dp_n591, dp_n590, dp_n589, dp_n588, dp_n587, dp_n586, dp_n585, 
      dp_n584, dp_n525, dp_n523, dp_n521, dp_n519, dp_n517, dp_n413, dp_n412, 
      dp_n411, dp_n410, dp_n409, dp_n408, dp_n407, dp_n406, dp_n405, dp_n404, 
      dp_n403, dp_n402, dp_n334, dp_n333, dp_n332, dp_n331, dp_n330, dp_n329, 
      dp_n328, dp_n327, dp_n326, dp_n325, dp_n324, dp_n323, dp_n322, dp_n321, 
      dp_n320, dp_n319, dp_n318, dp_n317, dp_n316, dp_n315, dp_n314, dp_n313, 
      dp_n312, dp_n311, dp_n310, dp_n309, dp_n308, dp_n307, dp_n306, dp_n305, 
      dp_n304, dp_n303, dp_n300, dp_n299, dp_n298, dp_n297, dp_n296, dp_n295, 
      dp_n294, dp_n293, dp_n292, dp_n291, dp_n290, dp_n289, dp_n288, dp_n287, 
      dp_n286, dp_n285, dp_n284, dp_n283, dp_n282, dp_n281, dp_n280, dp_n279, 
      dp_n278, dp_n277, dp_n276, dp_n275, dp_n274, dp_n273, dp_n272, dp_n271, 
      dp_n270, dp_n269, dp_n268, dp_n267, dp_n266, dp_n265, dp_n264, dp_n263, 
      dp_n262, dp_n261, dp_n260, dp_n259, dp_n258, dp_n257, dp_n256, dp_n255, 
      dp_n254, dp_n253, dp_n252, dp_n251, dp_n250, dp_n249, dp_n248, dp_n247, 
      dp_n246, dp_n245, dp_n244, dp_n243, dp_n242, dp_n241, dp_n240, dp_n239, 
      dp_n238, dp_n237, dp_n236, dp_n235, dp_n234, dp_n233, dp_n232, dp_n231, 
      dp_n230, dp_n229, dp_n228, dp_n227, dp_n226, dp_n225, dp_n224, dp_n223, 
      dp_n222, dp_n221, dp_n220, dp_n219, dp_n218, dp_n217, dp_n216, dp_n215, 
      dp_n214, dp_n213, dp_n212, dp_n211, dp_n210, dp_n209, dp_n208, dp_n207, 
      dp_n206, dp_n205, dp_n204, dp_n203, dp_n202, dp_n201, dp_n200, dp_n199, 
      dp_n198, dp_n197, dp_n196, dp_n195, dp_n194, dp_n193, dp_n192, dp_n191, 
      dp_n190, dp_n189, dp_n188, dp_n187, dp_n186, dp_n185, dp_n184, dp_n183, 
      dp_n182, dp_n181, dp_n180, dp_n179, dp_n178, dp_n177, dp_n176, dp_n175, 
      dp_n174, dp_n173, dp_n172, dp_n171, dp_n170, dp_n169, dp_n168, dp_n167, 
      dp_n166, dp_n165, dp_n164, dp_n163, dp_n162, dp_n161, dp_n160, dp_n159, 
      dp_n158, dp_n157, dp_n156, dp_n155, dp_n154, dp_n153, dp_n152, dp_n151, 
      dp_n150, dp_n149, dp_n148, dp_n147, dp_n146, dp_n145, dp_n144, dp_n143, 
      dp_n142, dp_n141, dp_n140, dp_n139, dp_n138, dp_n137, dp_n136, dp_n135, 
      dp_n134, dp_n133, dp_n130, dp_n129, dp_n128, dp_n127, dp_n126, dp_n125, 
      dp_n124, dp_n123, dp_n122, dp_n121, dp_n120, dp_n119, dp_n118, dp_n117, 
      dp_n116, dp_n115, dp_n114, dp_n113, dp_n112, dp_n111, dp_n110, dp_n109, 
      dp_n108, dp_n107, dp_n106, dp_n105, dp_n104, dp_n103, dp_n102, dp_n101, 
      dp_n100, dp_n99, dp_n98, dp_n97, dp_n96, dp_n95, dp_n94, dp_n93, dp_n92, 
      dp_n91, dp_n90, dp_n89, dp_n88, dp_n87, dp_n86, dp_n85, dp_n84, dp_n83, 
      dp_n82, dp_n81, dp_n80, dp_n79, dp_n78, dp_n77, dp_n76, dp_n75, dp_n74, 
      dp_n73, dp_n72, dp_n71, dp_n70, dp_n67, dp_n66, dp_n65, dp_n64, dp_n63, 
      dp_n62, dp_n61, dp_n60, dp_n59, dp_n58, dp_n57, dp_n56, dp_n55, dp_n54, 
      dp_n53, dp_n52, dp_n51, dp_n50, dp_n49, dp_n48, dp_n47, dp_n46, dp_n45, 
      dp_n44, dp_n43, dp_n42, dp_n41, dp_n40, dp_n39, dp_n38, dp_n37, dp_n36, 
      dp_n35, dp_n34, dp_n33, dp_n32, dp_n31, dp_n30, dp_n29, dp_n28, dp_n27, 
      dp_n26, dp_n25, dp_n24, dp_n23, dp_n22, dp_n21, dp_n20, dp_n19, dp_n18, 
      dp_n17, dp_n16, dp_n15, dp_n14, dp_n13, dp_n12, dp_n11, dp_n10, dp_n9, 
      dp_n8, dp_n7, dp_n6, dp_n5, dp_n4, dp_n3, dp_n1015, dp_n1014, dp_n1013, 
      dp_n1012, dp_n1011, dp_n1010, dp_n1009, dp_n1008, dp_n1007, dp_n1006, 
      dp_n1005, dp_n1004, dp_n1003, dp_n1002, dp_n1001, dp_n1000, dp_n999, 
      dp_n998, dp_n997, dp_n996, dp_n995, dp_n994, dp_n993, dp_n992, dp_n991, 
      dp_n990, dp_n989, dp_n988, dp_n987, dp_n986, dp_n985, dp_n984, dp_n983, 
      dp_n982, dp_n981, dp_n980, dp_n979, dp_n978, dp_n977, dp_n976, dp_n975, 
      dp_n974, dp_n973, dp_n972, dp_n971, dp_n970, dp_n969, dp_n968, dp_n967, 
      dp_n966, dp_n965, dp_n964, dp_n963, dp_n962, dp_n961, dp_n960, dp_n959, 
      dp_n958, dp_n957, dp_n956, dp_n955, dp_n954, dp_n953, dp_n952, dp_n951, 
      dp_n950, dp_n949, dp_n948, dp_n947, dp_n946, dp_n945, dp_n944, dp_n943, 
      dp_n942, dp_n941, dp_n940, dp_n939, dp_n938, dp_n937, dp_n936, dp_n935, 
      dp_n934, dp_n933, dp_n932, dp_n931, dp_n930, dp_n929, dp_n928, dp_n927, 
      dp_n926, dp_n925, dp_n924, dp_n923, dp_n922, dp_n921, dp_n920, dp_n919, 
      dp_n918, dp_n917, dp_n916, dp_n915, dp_n914, dp_n913, dp_n912, dp_n911, 
      dp_n910, dp_n909, dp_n908, dp_n907, dp_n906, dp_n905, dp_n904, dp_n903, 
      dp_n902, dp_n901, dp_n900, dp_n899, dp_n898, dp_n897, dp_n896, dp_n895, 
      dp_n894, dp_n893, dp_n892, dp_n891, dp_n890, dp_n889, dp_n888, dp_n887, 
      dp_n886, dp_n885, dp_n884, dp_n883, dp_n882, dp_n881, dp_n880, dp_n879, 
      dp_n878, dp_n877, dp_n876, dp_n875, dp_n874, dp_n873, dp_n872, dp_n871, 
      dp_n870, dp_n869, dp_n868, dp_n867, dp_n866, dp_n865, dp_n864, dp_n863, 
      dp_n862, dp_n861, dp_n860, dp_n859, dp_n858, dp_n857, dp_n856, dp_n855, 
      dp_n854, dp_n853, dp_n852, dp_n851, dp_n850, dp_n849, dp_n848, dp_n847, 
      dp_n846, dp_n845, dp_n844, dp_n843, dp_n842, dp_n841, dp_n840, dp_n839, 
      dp_n838, dp_n837, dp_n836, dp_n835, dp_n834, dp_n833, dp_n832, dp_n831, 
      dp_n830, dp_n829, dp_n828, dp_n827, dp_n826, dp_n825, dp_n824, dp_n823, 
      dp_n822, dp_n821, dp_n820, dp_n819, dp_n818, dp_n817, dp_n816, dp_n815, 
      dp_n814, dp_n813, dp_n812, dp_n811, dp_n810, dp_n809, dp_n808, dp_n807, 
      dp_n806, dp_n805, dp_n804, dp_n803, dp_n802, dp_n801, dp_n800, dp_n799, 
      dp_n798, dp_n797, dp_n796, dp_n795, dp_n794, dp_n793, dp_n792, dp_n791, 
      dp_n790, dp_n789, dp_n788, dp_n787, dp_n786, dp_n785, dp_n784, dp_n783, 
      dp_n782, dp_n781, dp_n780, dp_n779, dp_n778, dp_n777, dp_n776, dp_n775, 
      dp_n774, dp_n773, dp_n772, dp_n771, dp_n770, dp_n769, dp_n768, dp_n767, 
      dp_n766, dp_n765, dp_n764, dp_n763, dp_n762, dp_n761, dp_n760, dp_n759, 
      dp_n758, dp_n757, dp_n756, dp_n755, dp_n754, dp_n753, dp_n752, dp_n751, 
      dp_n750, dp_n749, dp_n748, dp_n747, dp_n746, dp_n745, dp_n744, dp_n743, 
      dp_n742, dp_n741, dp_n740, dp_n739, dp_n738, dp_n737, dp_n736, dp_n735, 
      dp_n734, dp_n733, dp_n732, dp_n731, dp_n730, dp_n729, dp_n728, dp_n727, 
      dp_n726, dp_n725, dp_n724, dp_n723, dp_n722, dp_n721, dp_n720, dp_n719, 
      dp_n718, dp_n717, dp_n716, dp_n715, dp_n714, dp_n713, dp_n712, dp_n706, 
      dp_n705, dp_n704, dp_n703, dp_n702, dp_n701, dp_n700, dp_n699, dp_n698, 
      dp_n697, dp_n696, dp_n695, dp_n694, dp_n693, dp_n692, dp_n691, dp_n690, 
      dp_n689, dp_n688, dp_n687, dp_n686, dp_n685, dp_n684, dp_n683, dp_n682, 
      dp_n681, dp_n680, dp_n679, dp_n678, dp_n677, dp_n676, dp_n675, dp_n674, 
      dp_n673, dp_n672, dp_n671, dp_n670, dp_n669, dp_n668, dp_n667, dp_n666, 
      dp_n665, dp_n664, dp_n663, dp_n662, dp_n661, dp_n660, dp_n659, dp_n658, 
      dp_n657, dp_n656, dp_n655, dp_n654, dp_n653, dp_n652, dp_n651, dp_n650, 
      dp_n649, dp_n583, dp_n582, dp_n581, dp_n580, dp_n579, dp_n578, dp_n577, 
      dp_n576, dp_n575, dp_n574, dp_n573, dp_n572, dp_n571, dp_n570, dp_n569, 
      dp_n568, dp_n567, dp_n566, dp_n565, dp_n564, dp_n563, dp_n562, dp_n561, 
      dp_n560, dp_n559, dp_n558, dp_n557, dp_n556, dp_n555, dp_n554, dp_n553, 
      dp_n552, dp_n551, dp_n550, dp_n549, dp_n548, dp_n547, dp_n546, dp_n545, 
      dp_n544, dp_n543, dp_n542, dp_n541, dp_n540, dp_n539, dp_n538, dp_n537, 
      dp_n536, dp_n535, dp_n534, dp_n533, dp_n532, dp_n531, dp_n530, dp_n529, 
      dp_n528, dp_n527, dp_n526, dp_n524, dp_n522, dp_n520, dp_n518, dp_n516, 
      dp_n515, dp_n514, dp_n513, dp_n512, dp_n511, dp_n510, dp_n509, dp_n508, 
      dp_n507, dp_n506, dp_n505, dp_n504, dp_n503, dp_n502, dp_n501, dp_n500, 
      dp_n499, dp_n498, dp_n497, dp_n496, dp_n495, dp_n494, dp_n493, dp_n492, 
      dp_n491, dp_n490, dp_n489, dp_n488, dp_n487, dp_n486, dp_n485, dp_n484, 
      dp_n483, dp_n482, dp_n481, dp_n480, dp_n479, dp_n478, dp_n477, dp_n476, 
      dp_n475, dp_n474, dp_n473, dp_n472, dp_n471, dp_n470, dp_n469, dp_n468, 
      dp_n467, dp_n466, dp_n465, dp_n464, dp_n463, dp_n462, dp_n461, dp_n460, 
      dp_n459, dp_n458, dp_n457, dp_n456, dp_n455, dp_n454, dp_n453, dp_n452, 
      dp_n451, dp_n450, dp_n449, dp_n448, dp_n447, dp_n446, dp_n445, dp_n444, 
      dp_n443, dp_n442, dp_n441, dp_n440, dp_n439, dp_n438, dp_n437, dp_n436, 
      dp_n435, dp_n434, dp_n433, dp_n432, dp_n431, dp_n430, dp_n429, dp_n428, 
      dp_n427, dp_n426, dp_n425, dp_n424, dp_n423, dp_n422, dp_n421, dp_n420, 
      dp_n419, dp_n418, dp_n417, dp_n416, dp_n415, dp_n414, dp_n401, dp_n400, 
      dp_n399, dp_n398, dp_n397, dp_n396, dp_n395, dp_n394, dp_n393, dp_n392, 
      dp_n391, dp_n390, dp_n389, dp_n388, dp_n387, dp_n386, dp_n385, dp_n384, 
      dp_n383, dp_n382, dp_n381, dp_n380, dp_n379, dp_n378, dp_n377, dp_n376, 
      dp_n375, dp_n374, dp_n373, dp_n372, dp_n371, dp_n370, dp_n369, dp_n368, 
      dp_n367, dp_n366, dp_n365, dp_n364, dp_n363, dp_n362, dp_n361, dp_n360, 
      dp_n359, dp_n358, dp_n357, dp_n356, dp_n355, dp_n354, dp_n353, dp_n352, 
      dp_n351, dp_n350, dp_n349, dp_n348, dp_n347, dp_n346, dp_n345, dp_n344, 
      dp_n343, dp_n342, dp_n341, dp_n340, dp_n339, dp_n338, dp_n337, dp_n336, 
      dp_n335, dp_n302, dp_n301, dp_n132, dp_n131, dp_n69, dp_n68, dp_n2, dp_n1
      , dp_z_word_0_port, dp_z_word_1_port, dp_z_word_2_port, dp_z_word_3_port,
      dp_z_word_4_port, dp_z_word_5_port, dp_z_word_6_port, dp_z_word_7_port, 
      dp_z_word_8_port, dp_z_word_9_port, dp_z_word_10_port, dp_z_word_11_port,
      dp_z_word_12_port, dp_z_word_13_port, dp_z_word_14_port, 
      dp_z_word_15_port, dp_z_word_16_port, dp_z_word_17_port, 
      dp_z_word_18_port, dp_z_word_19_port, dp_z_word_20_port, 
      dp_z_word_21_port, dp_z_word_22_port, dp_z_word_23_port, 
      dp_z_word_24_port, dp_z_word_25_port, dp_z_word_26_port, 
      dp_z_word_27_port, dp_z_word_28_port, dp_z_word_29_port, 
      dp_z_word_30_port, dp_z_word_31_port, dp_branch_t_ex_o, 
      dp_rd_fwd_ex_o_0_port, dp_rd_fwd_ex_o_1_port, dp_rd_fwd_ex_o_2_port, 
      dp_rd_fwd_ex_o_3_port, dp_rd_fwd_ex_o_4_port, dp_data_mem_ex_o_0_port, 
      dp_data_mem_ex_o_1_port, dp_data_mem_ex_o_2_port, dp_data_mem_ex_o_3_port
      , dp_data_mem_ex_o_4_port, dp_data_mem_ex_o_5_port, 
      dp_data_mem_ex_o_6_port, dp_data_mem_ex_o_7_port, dp_data_mem_ex_o_8_port
      , dp_data_mem_ex_o_9_port, dp_data_mem_ex_o_10_port, 
      dp_data_mem_ex_o_11_port, dp_data_mem_ex_o_12_port, 
      dp_data_mem_ex_o_13_port, dp_data_mem_ex_o_14_port, 
      dp_data_mem_ex_o_15_port, dp_data_mem_ex_o_16_port, 
      dp_data_mem_ex_o_17_port, dp_data_mem_ex_o_18_port, 
      dp_data_mem_ex_o_19_port, dp_data_mem_ex_o_20_port, 
      dp_data_mem_ex_o_21_port, dp_data_mem_ex_o_22_port, 
      dp_data_mem_ex_o_23_port, dp_data_mem_ex_o_24_port, 
      dp_data_mem_ex_o_25_port, dp_data_mem_ex_o_26_port, 
      dp_data_mem_ex_o_27_port, dp_data_mem_ex_o_28_port, 
      dp_data_mem_ex_o_29_port, dp_data_mem_ex_o_30_port, 
      dp_data_mem_ex_o_31_port, dp_alu_out_ex_o_0_port, dp_alu_out_ex_o_1_port,
      dp_alu_out_ex_o_2_port, dp_alu_out_ex_o_3_port, dp_alu_out_ex_o_4_port, 
      dp_alu_out_ex_o_5_port, dp_alu_out_ex_o_6_port, dp_alu_out_ex_o_7_port, 
      dp_alu_out_ex_o_8_port, dp_alu_out_ex_o_9_port, dp_alu_out_ex_o_10_port, 
      dp_alu_out_ex_o_11_port, dp_alu_out_ex_o_12_port, dp_alu_out_ex_o_13_port
      , dp_alu_out_ex_o_14_port, dp_alu_out_ex_o_15_port, 
      dp_alu_out_ex_o_16_port, dp_alu_out_ex_o_17_port, dp_alu_out_ex_o_18_port
      , dp_alu_out_ex_o_19_port, dp_alu_out_ex_o_20_port, 
      dp_alu_out_ex_o_21_port, dp_alu_out_ex_o_22_port, dp_alu_out_ex_o_23_port
      , dp_alu_out_ex_o_24_port, dp_alu_out_ex_o_25_port, 
      dp_alu_out_ex_o_26_port, dp_alu_out_ex_o_27_port, dp_alu_out_ex_o_28_port
      , dp_alu_out_ex_o_29_port, dp_alu_out_ex_o_30_port, 
      dp_alu_out_ex_o_31_port, dp_npc_ex_i_0_port, dp_npc_ex_i_1_port, 
      dp_npc_ex_i_2_port, dp_npc_ex_i_3_port, dp_npc_ex_i_4_port, 
      dp_npc_ex_i_5_port, dp_npc_ex_i_6_port, dp_npc_ex_i_7_port, 
      dp_npc_ex_i_8_port, dp_npc_ex_i_9_port, dp_npc_ex_i_10_port, 
      dp_npc_ex_i_11_port, dp_npc_ex_i_12_port, dp_npc_ex_i_13_port, 
      dp_npc_ex_i_14_port, dp_npc_ex_i_15_port, dp_npc_ex_i_16_port, 
      dp_npc_ex_i_17_port, dp_npc_ex_i_18_port, dp_npc_ex_i_19_port, 
      dp_npc_ex_i_20_port, dp_npc_ex_i_21_port, dp_npc_ex_i_22_port, 
      dp_npc_ex_i_23_port, dp_npc_ex_i_24_port, dp_npc_ex_i_25_port, 
      dp_npc_ex_i_26_port, dp_npc_ex_i_27_port, dp_npc_ex_i_28_port, 
      dp_npc_ex_i_29_port, dp_npc_ex_i_30_port, dp_npc_ex_i_31_port, 
      dp_imm_ex_i_0_port, dp_imm_ex_i_1_port, dp_imm_ex_i_2_port, 
      dp_imm_ex_i_3_port, dp_imm_ex_i_4_port, dp_imm_ex_i_5_port, 
      dp_imm_ex_i_6_port, dp_imm_ex_i_7_port, dp_imm_ex_i_8_port, 
      dp_imm_ex_i_9_port, dp_imm_ex_i_10_port, dp_imm_ex_i_11_port, 
      dp_imm_ex_i_12_port, dp_imm_ex_i_13_port, dp_imm_ex_i_14_port, 
      dp_imm_ex_i_15_port, dp_imm_ex_i_16_port, dp_imm_ex_i_17_port, 
      dp_imm_ex_i_18_port, dp_imm_ex_i_19_port, dp_imm_ex_i_20_port, 
      dp_imm_ex_i_21_port, dp_imm_ex_i_22_port, dp_imm_ex_i_23_port, 
      dp_imm_ex_i_24_port, dp_imm_ex_i_25_port, dp_imm_ex_i_26_port, 
      dp_imm_ex_i_27_port, dp_imm_ex_i_28_port, dp_imm_ex_i_29_port, 
      dp_imm_ex_i_30_port, dp_imm_ex_i_31_port, dp_rf_out1_ex_i_0_port, 
      dp_rf_out1_ex_i_1_port, dp_rf_out1_ex_i_2_port, dp_rf_out1_ex_i_3_port, 
      dp_rf_out1_ex_i_4_port, dp_rf_out1_ex_i_5_port, dp_rf_out1_ex_i_6_port, 
      dp_rf_out1_ex_i_7_port, dp_rf_out1_ex_i_8_port, dp_rf_out1_ex_i_9_port, 
      dp_rf_out1_ex_i_10_port, dp_rf_out1_ex_i_11_port, dp_rf_out1_ex_i_12_port
      , dp_rf_out1_ex_i_13_port, dp_rf_out1_ex_i_14_port, 
      dp_rf_out1_ex_i_15_port, dp_rf_out1_ex_i_16_port, dp_rf_out1_ex_i_17_port
      , dp_rf_out1_ex_i_18_port, dp_rf_out1_ex_i_19_port, 
      dp_rf_out1_ex_i_20_port, dp_rf_out1_ex_i_21_port, dp_rf_out1_ex_i_22_port
      , dp_rf_out1_ex_i_23_port, dp_rf_out1_ex_i_24_port, 
      dp_rf_out1_ex_i_25_port, dp_rf_out1_ex_i_26_port, dp_rf_out1_ex_i_27_port
      , dp_rf_out1_ex_i_28_port, dp_rf_out1_ex_i_29_port, 
      dp_rf_out1_ex_i_30_port, dp_rf_out1_ex_i_31_port, dp_rd_fwd_id_o_0_port, 
      dp_rd_fwd_id_o_1_port, dp_rd_fwd_id_o_2_port, dp_rd_fwd_id_o_3_port, 
      dp_rd_fwd_id_o_4_port, dp_npc_id_o_0_port, dp_npc_id_o_1_port, 
      dp_npc_id_o_2_port, dp_npc_id_o_3_port, dp_npc_id_o_4_port, 
      dp_npc_id_o_5_port, dp_npc_id_o_6_port, dp_npc_id_o_7_port, 
      dp_npc_id_o_8_port, dp_npc_id_o_9_port, dp_npc_id_o_10_port, 
      dp_npc_id_o_11_port, dp_npc_id_o_12_port, dp_npc_id_o_13_port, 
      dp_npc_id_o_14_port, dp_npc_id_o_15_port, dp_npc_id_o_16_port, 
      dp_npc_id_o_17_port, dp_npc_id_o_18_port, dp_npc_id_o_19_port, 
      dp_npc_id_o_20_port, dp_npc_id_o_21_port, dp_npc_id_o_22_port, 
      dp_npc_id_o_23_port, dp_npc_id_o_24_port, dp_npc_id_o_25_port, 
      dp_npc_id_o_26_port, dp_npc_id_o_27_port, dp_npc_id_o_28_port, 
      dp_npc_id_o_29_port, dp_npc_id_o_30_port, dp_npc_id_o_31_port, 
      dp_imm_id_o_0_port, dp_imm_id_o_1_port, dp_imm_id_o_2_port, 
      dp_imm_id_o_3_port, dp_imm_id_o_4_port, dp_imm_id_o_5_port, 
      dp_imm_id_o_6_port, dp_imm_id_o_7_port, dp_imm_id_o_8_port, 
      dp_imm_id_o_9_port, dp_imm_id_o_10_port, dp_imm_id_o_11_port, 
      dp_imm_id_o_12_port, dp_imm_id_o_13_port, dp_imm_id_o_14_port, 
      dp_imm_id_o_15_port, dp_imm_id_o_16_port, dp_imm_id_o_17_port, 
      dp_imm_id_o_18_port, dp_imm_id_o_19_port, dp_imm_id_o_20_port, 
      dp_imm_id_o_21_port, dp_imm_id_o_22_port, dp_imm_id_o_23_port, 
      dp_imm_id_o_24_port, dp_imm_id_o_31_port, dp_rf_out2_id_o_0_port, 
      dp_rf_out2_id_o_1_port, dp_rf_out2_id_o_2_port, dp_rf_out2_id_o_3_port, 
      dp_rf_out2_id_o_4_port, dp_rf_out2_id_o_5_port, dp_rf_out2_id_o_6_port, 
      dp_rf_out2_id_o_7_port, dp_rf_out2_id_o_8_port, dp_rf_out2_id_o_9_port, 
      dp_rf_out2_id_o_10_port, dp_rf_out2_id_o_11_port, dp_rf_out2_id_o_12_port
      , dp_rf_out2_id_o_13_port, dp_rf_out2_id_o_14_port, 
      dp_rf_out2_id_o_15_port, dp_rf_out2_id_o_16_port, dp_rf_out2_id_o_17_port
      , dp_rf_out2_id_o_18_port, dp_rf_out2_id_o_19_port, 
      dp_rf_out2_id_o_20_port, dp_rf_out2_id_o_21_port, dp_rf_out2_id_o_22_port
      , dp_rf_out2_id_o_23_port, dp_rf_out2_id_o_24_port, 
      dp_rf_out2_id_o_25_port, dp_rf_out2_id_o_26_port, dp_rf_out2_id_o_27_port
      , dp_rf_out2_id_o_28_port, dp_rf_out2_id_o_29_port, 
      dp_rf_out2_id_o_30_port, dp_rf_out2_id_o_31_port, dp_rf_out1_id_o_0_port,
      dp_rf_out1_id_o_1_port, dp_rf_out1_id_o_2_port, dp_rf_out1_id_o_3_port, 
      dp_rf_out1_id_o_4_port, dp_rf_out1_id_o_5_port, dp_rf_out1_id_o_6_port, 
      dp_rf_out1_id_o_7_port, dp_rf_out1_id_o_8_port, dp_rf_out1_id_o_9_port, 
      dp_rf_out1_id_o_10_port, dp_rf_out1_id_o_11_port, dp_rf_out1_id_o_12_port
      , dp_rf_out1_id_o_13_port, dp_rf_out1_id_o_14_port, 
      dp_rf_out1_id_o_15_port, dp_rf_out1_id_o_16_port, dp_rf_out1_id_o_17_port
      , dp_rf_out1_id_o_18_port, dp_rf_out1_id_o_19_port, 
      dp_rf_out1_id_o_20_port, dp_rf_out1_id_o_21_port, dp_rf_out1_id_o_22_port
      , dp_rf_out1_id_o_23_port, dp_rf_out1_id_o_24_port, 
      dp_rf_out1_id_o_25_port, dp_rf_out1_id_o_26_port, dp_rf_out1_id_o_27_port
      , dp_rf_out1_id_o_28_port, dp_rf_out1_id_o_29_port, 
      dp_rf_out1_id_o_30_port, dp_rf_out1_id_o_31_port, dp_wr_data_id_i_0_port,
      dp_wr_data_id_i_1_port, dp_wr_data_id_i_2_port, dp_wr_data_id_i_3_port, 
      dp_wr_data_id_i_4_port, dp_wr_data_id_i_5_port, dp_wr_data_id_i_6_port, 
      dp_wr_data_id_i_7_port, dp_wr_data_id_i_8_port, dp_wr_data_id_i_9_port, 
      dp_wr_data_id_i_10_port, dp_wr_data_id_i_11_port, dp_wr_data_id_i_12_port
      , dp_wr_data_id_i_13_port, dp_wr_data_id_i_14_port, 
      dp_wr_data_id_i_15_port, dp_wr_data_id_i_16_port, dp_wr_data_id_i_17_port
      , dp_wr_data_id_i_18_port, dp_wr_data_id_i_19_port, 
      dp_wr_data_id_i_20_port, dp_wr_data_id_i_21_port, dp_wr_data_id_i_22_port
      , dp_wr_data_id_i_23_port, dp_wr_data_id_i_24_port, 
      dp_wr_data_id_i_25_port, dp_wr_data_id_i_26_port, dp_wr_data_id_i_27_port
      , dp_wr_data_id_i_28_port, dp_wr_data_id_i_29_port, 
      dp_wr_data_id_i_30_port, dp_wr_data_id_i_31_port, dp_rd_fwd_wb_i_0_port, 
      dp_rd_fwd_wb_i_1_port, dp_rd_fwd_wb_i_2_port, dp_rd_fwd_wb_i_3_port, 
      dp_rd_fwd_wb_i_4_port, dp_ir_0_port, dp_ir_1_port, dp_ir_2_port, 
      dp_ir_3_port, dp_ir_4_port, dp_ir_5_port, dp_ir_6_port, dp_ir_7_port, 
      dp_ir_8_port, dp_ir_9_port, dp_ir_10_port, dp_ir_11_port, dp_ir_12_port, 
      dp_ir_13_port, dp_ir_14_port, dp_ir_15_port, dp_ir_16_port, dp_ir_17_port
      , dp_ir_18_port, dp_ir_19_port, dp_ir_20_port, dp_ir_21_port, 
      dp_ir_22_port, dp_ir_23_port, dp_ir_24_port, dp_ir_25_port, 
      dp_npc_if_o_0_port, dp_npc_if_o_1_port, dp_npc_if_o_2_port, 
      dp_npc_if_o_3_port, dp_npc_if_o_4_port, dp_npc_if_o_5_port, 
      dp_npc_if_o_6_port, dp_npc_if_o_7_port, dp_npc_if_o_8_port, 
      dp_npc_if_o_9_port, dp_npc_if_o_10_port, dp_npc_if_o_11_port, 
      dp_npc_if_o_12_port, dp_npc_if_o_13_port, dp_npc_if_o_14_port, 
      dp_npc_if_o_15_port, dp_npc_if_o_16_port, dp_npc_if_o_17_port, 
      dp_npc_if_o_18_port, dp_npc_if_o_19_port, dp_npc_if_o_20_port, 
      dp_npc_if_o_21_port, dp_npc_if_o_22_port, dp_npc_if_o_23_port, 
      dp_npc_if_o_24_port, dp_npc_if_o_25_port, dp_npc_if_o_26_port, 
      dp_npc_if_o_27_port, dp_npc_if_o_28_port, dp_npc_if_o_29_port, 
      dp_npc_if_o_30_port, dp_npc_if_o_31_port, dp_if_stage_n41, 
      dp_if_stage_n40, dp_if_stage_n39, dp_if_stage_n38, dp_if_stage_n37, 
      dp_if_stage_n36, dp_if_stage_n35, dp_if_stage_n34, dp_if_stage_n33, 
      dp_if_stage_n16, dp_if_stage_n15, dp_if_stage_n14, dp_if_stage_n13, 
      dp_if_stage_n12, dp_if_stage_n11, dp_if_stage_n10, dp_if_stage_n9, 
      dp_if_stage_n8, dp_if_stage_n7, dp_if_stage_n6, dp_if_stage_n5, 
      dp_if_stage_n4, dp_if_stage_n3, dp_if_stage_n2, dp_if_stage_n1, 
      dp_if_stage_n98, dp_if_stage_n97, dp_if_stage_n95, dp_if_stage_n94, 
      dp_if_stage_n93, dp_if_stage_n92, dp_if_stage_n91, dp_if_stage_n90, 
      dp_if_stage_n89, dp_if_stage_n88, dp_if_stage_n87, dp_if_stage_n86, 
      dp_if_stage_n85, dp_if_stage_n84, dp_if_stage_n83, dp_if_stage_n82, 
      dp_if_stage_n81, dp_if_stage_n64, dp_if_stage_n63, dp_if_stage_n62, 
      dp_if_stage_n61, dp_if_stage_n60, dp_if_stage_n59, dp_if_stage_n58, 
      dp_if_stage_n57, dp_if_stage_n56, dp_if_stage_n55, dp_if_stage_n54, 
      dp_if_stage_n53, dp_if_stage_n52, dp_if_stage_n51, dp_if_stage_n50, 
      dp_if_stage_n49, dp_if_stage_n32, dp_if_stage_n31, dp_if_stage_n30, 
      dp_if_stage_n29, dp_if_stage_n28, dp_if_stage_n27, dp_if_stage_n26, 
      dp_if_stage_n25, dp_if_stage_n24, dp_if_stage_n23, dp_if_stage_n22, 
      dp_if_stage_n21, dp_if_stage_n20, dp_if_stage_n19, dp_if_stage_n18, 
      dp_if_stage_n17, dp_if_stage_NPC_4_i_0_port, dp_if_stage_NPC_4_i_1_port, 
      dp_if_stage_NPC_4_i_2_port, dp_if_stage_NPC_4_i_3_port, 
      dp_if_stage_NPC_4_i_4_port, dp_if_stage_NPC_4_i_5_port, 
      dp_if_stage_NPC_4_i_6_port, dp_if_stage_NPC_4_i_7_port, 
      dp_if_stage_NPC_4_i_8_port, dp_if_stage_NPC_4_i_9_port, 
      dp_if_stage_NPC_4_i_10_port, dp_if_stage_NPC_4_i_11_port, 
      dp_if_stage_NPC_4_i_12_port, dp_if_stage_NPC_4_i_13_port, 
      dp_if_stage_NPC_4_i_14_port, dp_if_stage_NPC_4_i_15_port, 
      dp_if_stage_NPC_4_i_16_port, dp_if_stage_NPC_4_i_17_port, 
      dp_if_stage_NPC_4_i_18_port, dp_if_stage_NPC_4_i_19_port, 
      dp_if_stage_NPC_4_i_20_port, dp_if_stage_NPC_4_i_21_port, 
      dp_if_stage_NPC_4_i_22_port, dp_if_stage_NPC_4_i_23_port, 
      dp_if_stage_NPC_4_i_24_port, dp_if_stage_NPC_4_i_25_port, 
      dp_if_stage_NPC_4_i_26_port, dp_if_stage_NPC_4_i_27_port, 
      dp_if_stage_NPC_4_i_28_port, dp_if_stage_NPC_4_i_29_port, 
      dp_if_stage_NPC_4_i_30_port, dp_if_stage_NPC_4_i_31_port, 
      dp_if_stage_Logic0_port, dp_if_stage_Logic1_port, dp_if_stage_mux_n7, 
      dp_if_stage_mux_n6, dp_if_stage_mux_n5, dp_if_stage_mux_n4, 
      dp_if_stage_mux_n3, dp_if_stage_mux_n2, dp_if_stage_mux_n1, 
      dp_if_stage_mux_n65, dp_if_stage_mux_n64, dp_if_stage_mux_n63, 
      dp_if_stage_mux_n62, dp_if_stage_mux_n61, dp_if_stage_mux_n60, 
      dp_if_stage_mux_n59, dp_if_stage_mux_n54, dp_if_stage_mux_n43, 
      dp_if_stage_mux_n40, dp_if_stage_mux_n39, dp_if_stage_mux_n38, 
      dp_if_stage_mux_n37, dp_if_stage_mux_n36, dp_if_stage_mux_n35, 
      dp_if_stage_mux_n34, dp_if_stage_add_77_n61, dp_if_stage_add_77_n60, 
      dp_if_stage_add_77_n59, dp_if_stage_add_77_n58, dp_if_stage_add_77_n57, 
      dp_if_stage_add_77_n56, dp_if_stage_add_77_n55, dp_if_stage_add_77_n54, 
      dp_if_stage_add_77_n53, dp_if_stage_add_77_n52, dp_if_stage_add_77_n51, 
      dp_if_stage_add_77_n50, dp_if_stage_add_77_n49, dp_if_stage_add_77_n48, 
      dp_if_stage_add_77_n47, dp_if_stage_add_77_n46, dp_if_stage_add_77_n45, 
      dp_if_stage_add_77_n44, dp_if_stage_add_77_n43, dp_if_stage_add_77_n42, 
      dp_if_stage_add_77_n41, dp_if_stage_add_77_n40, dp_if_stage_add_77_n39, 
      dp_if_stage_add_77_n38, dp_if_stage_add_77_n37, dp_if_stage_add_77_n36, 
      dp_if_stage_add_77_n35, dp_if_stage_add_77_n34, dp_if_stage_add_77_n33, 
      dp_if_stage_add_77_n32, dp_if_stage_add_77_n31, dp_if_stage_add_77_n30, 
      dp_if_stage_add_77_n29, dp_if_stage_add_77_n28, dp_if_stage_add_77_n27, 
      dp_if_stage_add_77_n26, dp_if_stage_add_77_n25, dp_if_stage_add_77_n24, 
      dp_if_stage_add_77_n23, dp_if_stage_add_77_n22, dp_if_stage_add_77_n21, 
      dp_if_stage_add_77_n20, dp_if_stage_add_77_n19, dp_if_stage_add_77_n18, 
      dp_if_stage_add_77_n16, dp_if_stage_add_77_n15, dp_if_stage_add_77_n14, 
      dp_if_stage_add_77_n13, dp_if_stage_add_77_n12, dp_if_stage_add_77_n11, 
      dp_if_stage_add_77_n10, dp_if_stage_add_77_n9, dp_if_stage_add_77_n8, 
      dp_if_stage_add_77_n7, dp_if_stage_add_77_n6, dp_if_stage_add_77_n5, 
      dp_if_stage_add_77_n4, dp_if_stage_add_77_n3, dp_if_stage_add_77_n2, 
      dp_if_stage_add_77_n1, dp_id_stage_n40, dp_id_stage_n39, dp_id_stage_n38,
      dp_id_stage_n37, dp_id_stage_n36, dp_id_stage_n35, dp_id_stage_n34, 
      dp_id_stage_n33, dp_id_stage_n32, dp_id_stage_n31, dp_id_stage_n30, 
      dp_id_stage_n29, dp_id_stage_n28, dp_id_stage_n27, dp_id_stage_n26, 
      dp_id_stage_n25, dp_id_stage_n24, dp_id_stage_n16, dp_id_stage_n15, 
      dp_id_stage_n14, dp_id_stage_n13, dp_id_stage_n12, dp_id_stage_n11, 
      dp_id_stage_n10, dp_id_stage_n9, dp_id_stage_n8, dp_id_stage_n7, 
      dp_id_stage_n6, dp_id_stage_n5, dp_id_stage_n4, dp_id_stage_n3, 
      dp_id_stage_n2, dp_id_stage_n1, dp_id_stage_n23, dp_id_stage_n22, 
      dp_id_stage_n21, dp_id_stage_n20, dp_id_stage_n19, dp_id_stage_n18, 
      dp_id_stage_n17, dp_id_stage_out2_i_0_port, dp_id_stage_out2_i_1_port, 
      dp_id_stage_out2_i_2_port, dp_id_stage_out2_i_3_port, 
      dp_id_stage_out2_i_4_port, dp_id_stage_out2_i_5_port, 
      dp_id_stage_out2_i_6_port, dp_id_stage_out2_i_7_port, 
      dp_id_stage_out2_i_8_port, dp_id_stage_out2_i_9_port, 
      dp_id_stage_out2_i_10_port, dp_id_stage_out2_i_11_port, 
      dp_id_stage_out2_i_12_port, dp_id_stage_out2_i_13_port, 
      dp_id_stage_out2_i_14_port, dp_id_stage_out2_i_15_port, 
      dp_id_stage_out2_i_16_port, dp_id_stage_out2_i_17_port, 
      dp_id_stage_out2_i_18_port, dp_id_stage_out2_i_19_port, 
      dp_id_stage_out2_i_20_port, dp_id_stage_out2_i_21_port, 
      dp_id_stage_out2_i_22_port, dp_id_stage_out2_i_23_port, 
      dp_id_stage_out2_i_24_port, dp_id_stage_out2_i_25_port, 
      dp_id_stage_out2_i_26_port, dp_id_stage_out2_i_27_port, 
      dp_id_stage_out2_i_28_port, dp_id_stage_out2_i_29_port, 
      dp_id_stage_out2_i_30_port, dp_id_stage_out2_i_31_port, 
      dp_id_stage_out1_i_0_port, dp_id_stage_out1_i_1_port, 
      dp_id_stage_out1_i_2_port, dp_id_stage_out1_i_3_port, 
      dp_id_stage_out1_i_4_port, dp_id_stage_out1_i_5_port, 
      dp_id_stage_out1_i_6_port, dp_id_stage_out1_i_7_port, 
      dp_id_stage_out1_i_8_port, dp_id_stage_out1_i_9_port, 
      dp_id_stage_out1_i_10_port, dp_id_stage_out1_i_11_port, 
      dp_id_stage_out1_i_12_port, dp_id_stage_out1_i_13_port, 
      dp_id_stage_out1_i_14_port, dp_id_stage_out1_i_15_port, 
      dp_id_stage_out1_i_16_port, dp_id_stage_out1_i_17_port, 
      dp_id_stage_out1_i_18_port, dp_id_stage_out1_i_19_port, 
      dp_id_stage_out1_i_20_port, dp_id_stage_out1_i_21_port, 
      dp_id_stage_out1_i_22_port, dp_id_stage_out1_i_23_port, 
      dp_id_stage_out1_i_24_port, dp_id_stage_out1_i_25_port, 
      dp_id_stage_out1_i_26_port, dp_id_stage_out1_i_27_port, 
      dp_id_stage_out1_i_28_port, dp_id_stage_out1_i_29_port, 
      dp_id_stage_out1_i_30_port, dp_id_stage_out1_i_31_port, 
      dp_id_stage_p_addr_wRD_0_port, dp_id_stage_p_addr_wRD_1_port, 
      dp_id_stage_p_addr_wRD_2_port, dp_id_stage_p_addr_wRD_3_port, 
      dp_id_stage_p_addr_wRD_4_port, dp_id_stage_p_addr_wRS2_0_port, 
      dp_id_stage_p_addr_wRS2_1_port, dp_id_stage_p_addr_wRS2_2_port, 
      dp_id_stage_p_addr_wRS2_3_port, dp_id_stage_p_addr_wRS2_4_port, 
      dp_id_stage_p_addr_wRS1_0_port, dp_id_stage_p_addr_wRS1_1_port, 
      dp_id_stage_p_addr_wRS1_2_port, dp_id_stage_p_addr_wRS1_3_port, 
      dp_id_stage_p_addr_wRS1_4_port, dp_id_stage_regfile_cpu_work, 
      dp_id_stage_regfile_sel_wp, dp_id_stage_regfile_end_sf, 
      dp_id_stage_regfile_canrestore, dp_id_stage_regfile_cansave, 
      dp_id_stage_regfile_up_dwn_rest, dp_id_stage_regfile_up_dwn_save, 
      dp_id_stage_regfile_up_dwn_cwp, dp_id_stage_regfile_up_dwn_swp, 
      dp_id_stage_regfile_rst_spill_fill, dp_id_stage_regfile_rst_swp, 
      dp_id_stage_regfile_cnt_save, dp_id_stage_regfile_cnt_cwp, 
      dp_id_stage_regfile_cnt_swp, dp_id_stage_regfile_rst_rf, 
      dp_id_stage_regfile_rf_enable, dp_id_stage_regfile_wr_cu, 
      dp_id_stage_regfile_rd_cu, dp_id_stage_regfile_ControlUnit_n41, 
      dp_id_stage_regfile_ControlUnit_n15, dp_id_stage_regfile_ControlUnit_n10,
      dp_id_stage_regfile_ControlUnit_n9, dp_id_stage_regfile_ControlUnit_n6, 
      dp_id_stage_regfile_ControlUnit_n5, dp_id_stage_regfile_ControlUnit_n4, 
      dp_id_stage_regfile_ControlUnit_n3, dp_id_stage_regfile_ControlUnit_n1, 
      dp_id_stage_regfile_ControlUnit_n40, dp_id_stage_regfile_ControlUnit_n39,
      dp_id_stage_regfile_ControlUnit_n38, dp_id_stage_regfile_ControlUnit_n37,
      dp_id_stage_regfile_ControlUnit_n36, dp_id_stage_regfile_ControlUnit_n35,
      dp_id_stage_regfile_ControlUnit_n34, dp_id_stage_regfile_ControlUnit_n33,
      dp_id_stage_regfile_ControlUnit_n32, dp_id_stage_regfile_ControlUnit_n31,
      dp_id_stage_regfile_ControlUnit_n30, dp_id_stage_regfile_ControlUnit_n29,
      dp_id_stage_regfile_ControlUnit_n28, dp_id_stage_regfile_ControlUnit_n27,
      dp_id_stage_regfile_ControlUnit_n26, dp_id_stage_regfile_ControlUnit_n25,
      dp_id_stage_regfile_ControlUnit_n24, dp_id_stage_regfile_ControlUnit_n23,
      dp_id_stage_regfile_ControlUnit_n22, dp_id_stage_regfile_ControlUnit_n21,
      dp_id_stage_regfile_ControlUnit_n20, dp_id_stage_regfile_ControlUnit_n19,
      dp_id_stage_regfile_ControlUnit_n18, dp_id_stage_regfile_ControlUnit_n17,
      dp_id_stage_regfile_ControlUnit_n16, dp_id_stage_regfile_ControlUnit_n14,
      dp_id_stage_regfile_ControlUnit_n13, dp_id_stage_regfile_ControlUnit_n12,
      dp_id_stage_regfile_ControlUnit_current_state_0_port, 
      dp_id_stage_regfile_ControlUnit_current_state_2_port, 
      dp_id_stage_regfile_ControlUnit_current_state_3_port, 
      dp_id_stage_regfile_ControlUnit_next_state_0_port, 
      dp_id_stage_regfile_ControlUnit_next_state_1_port, 
      dp_id_stage_regfile_ControlUnit_next_state_2_port, 
      dp_id_stage_regfile_ControlUnit_next_state_3_port, 
      dp_id_stage_regfile_DataPath_mux_en_control_out, 
      dp_id_stage_regfile_DataPath_mux_wr_control_out, 
      dp_id_stage_regfile_DataPath_mux_rd2_control_out, 
      dp_id_stage_regfile_DataPath_mux_rd1_control_out, 
      dp_id_stage_regfile_DataPath_mux_wr_out_0_port, 
      dp_id_stage_regfile_DataPath_mux_wr_out_1_port, 
      dp_id_stage_regfile_DataPath_mux_wr_out_2_port, 
      dp_id_stage_regfile_DataPath_mux_wr_out_3_port, 
      dp_id_stage_regfile_DataPath_mux_wr_out_4_port, 
      dp_id_stage_regfile_DataPath_mux_wr_out_5_port, 
      dp_id_stage_regfile_DataPath_mux_rd_out_0_port, 
      dp_id_stage_regfile_DataPath_mux_rd_out_1_port, 
      dp_id_stage_regfile_DataPath_mux_rd_out_2_port, 
      dp_id_stage_regfile_DataPath_mux_rd_out_3_port, 
      dp_id_stage_regfile_DataPath_mux_rd_out_4_port, 
      dp_id_stage_regfile_DataPath_mux_rd_out_5_port, 
      dp_id_stage_regfile_DataPath_cwp_1_0_port, 
      dp_id_stage_regfile_DataPath_spill_fill_addr_0_port, 
      dp_id_stage_regfile_DataPath_spill_fill_addr_1_port, 
      dp_id_stage_regfile_DataPath_spill_fill_addr_2_port, 
      dp_id_stage_regfile_DataPath_spill_fill_addr_3_port, 
      dp_id_stage_regfile_DataPath_spill_fill_addr_4_port, 
      dp_id_stage_regfile_DataPath_spill_fill_addr_5_port, 
      dp_id_stage_regfile_DataPath_sf_wp_0_port, 
      dp_id_stage_regfile_DataPath_addr_sf_in_0_port, 
      dp_id_stage_regfile_DataPath_addr_sf_in_1_port, 
      dp_id_stage_regfile_DataPath_addr_sf_in_2_port, 
      dp_id_stage_regfile_DataPath_addr_w_p_0_port, 
      dp_id_stage_regfile_DataPath_addr_w_p_1_port, 
      dp_id_stage_regfile_DataPath_addr_w_p_2_port, 
      dp_id_stage_regfile_DataPath_addr_w_p_3_port, 
      dp_id_stage_regfile_DataPath_addr_w_p_4_port, 
      dp_id_stage_regfile_DataPath_addr_w_p_5_port, 
      dp_id_stage_regfile_DataPath_addr_rd2_p_0_port, 
      dp_id_stage_regfile_DataPath_addr_rd2_p_1_port, 
      dp_id_stage_regfile_DataPath_addr_rd2_p_2_port, 
      dp_id_stage_regfile_DataPath_addr_rd2_p_3_port, 
      dp_id_stage_regfile_DataPath_addr_rd2_p_4_port, 
      dp_id_stage_regfile_DataPath_addr_rd2_p_5_port, 
      dp_id_stage_regfile_DataPath_addr_rd1_p_0_port, 
      dp_id_stage_regfile_DataPath_addr_rd1_p_1_port, 
      dp_id_stage_regfile_DataPath_addr_rd1_p_2_port, 
      dp_id_stage_regfile_DataPath_addr_rd1_p_3_port, 
      dp_id_stage_regfile_DataPath_addr_rd1_p_4_port, 
      dp_id_stage_regfile_DataPath_addr_rd1_p_5_port, 
      dp_id_stage_regfile_DataPath_CWP_0_port, 
      dp_id_stage_regfile_DataPath_Logic0_port, 
      dp_id_stage_regfile_DataPath_Logic1_port, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n8, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n4, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n3, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n2, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n1, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n22, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n21, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n20, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n19, 
      dp_id_stage_regfile_DataPath_Conv_RD1_n18, 
      dp_id_stage_regfile_DataPath_Conv_RD1_N5, 
      dp_id_stage_regfile_DataPath_Conv_RD1_N1_port, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n13, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n12, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n11, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n10, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n9, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n8, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n4, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n3, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n2, 
      dp_id_stage_regfile_DataPath_Conv_RD2_n1, 
      dp_id_stage_regfile_DataPath_Conv_RD2_N5, 
      dp_id_stage_regfile_DataPath_Conv_RD2_N1_port, 
      dp_id_stage_regfile_DataPath_Conv_W_n13, 
      dp_id_stage_regfile_DataPath_Conv_W_n12, 
      dp_id_stage_regfile_DataPath_Conv_W_n11, 
      dp_id_stage_regfile_DataPath_Conv_W_n10, 
      dp_id_stage_regfile_DataPath_Conv_W_n9, 
      dp_id_stage_regfile_DataPath_Conv_W_n8, 
      dp_id_stage_regfile_DataPath_Conv_W_n4, 
      dp_id_stage_regfile_DataPath_Conv_W_n3, 
      dp_id_stage_regfile_DataPath_Conv_W_n2, 
      dp_id_stage_regfile_DataPath_Conv_W_n1, 
      dp_id_stage_regfile_DataPath_Conv_W_N5, 
      dp_id_stage_regfile_DataPath_Conv_W_N1_port, 
      dp_id_stage_regfile_DataPath_SF_converter_n10, 
      dp_id_stage_regfile_DataPath_SF_converter_n9, 
      dp_id_stage_regfile_DataPath_SF_converter_n8, 
      dp_id_stage_regfile_DataPath_SF_converter_n7, 
      dp_id_stage_regfile_DataPath_SF_converter_n6, 
      dp_id_stage_regfile_DataPath_SF_converter_n5, 
      dp_id_stage_regfile_DataPath_SF_converter_n4, 
      dp_id_stage_regfile_DataPath_SF_converter_n3, 
      dp_id_stage_regfile_DataPath_SF_converter_n2, 
      dp_id_stage_regfile_DataPath_SF_converter_n1, 
      dp_id_stage_regfile_DataPath_SF_converter_N5_port, 
      dp_id_stage_regfile_DataPath_SF_converter_N1_port, 
      dp_id_stage_regfile_DataPath_Cwp_counter_n4, 
      dp_id_stage_regfile_DataPath_Cwp_counter_n2, 
      dp_id_stage_regfile_DataPath_Cwp_counter_n5, 
      dp_id_stage_regfile_DataPath_Cwp_counter_n3, 
      dp_id_stage_regfile_DataPath_Cwp_counter_n1, 
      dp_id_stage_regfile_DataPath_Swp_counter_n8, 
      dp_id_stage_regfile_DataPath_Swp_counter_n7, 
      dp_id_stage_regfile_DataPath_Swp_counter_n6, 
      dp_id_stage_regfile_DataPath_Swp_counter_n4, 
      dp_id_stage_regfile_DataPath_Swp_counter_n2, 
      dp_id_stage_regfile_DataPath_Swp_counter_Q_0_port, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n16, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n12, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n4, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n3, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n2, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n1, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n21, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n20, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n19, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n18, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n17, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n15, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n14, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n13, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n11, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n10, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n9, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n8, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n7, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n6, 
      dp_id_stage_regfile_DataPath_Spill_fill_counter_n5, 
      dp_id_stage_regfile_DataPath_CANSAVE_counter_n8, 
      dp_id_stage_regfile_DataPath_CANSAVE_counter_n7, 
      dp_id_stage_regfile_DataPath_CANSAVE_counter_n6, 
      dp_id_stage_regfile_DataPath_CANSAVE_counter_n4, 
      dp_id_stage_regfile_DataPath_CANSAVE_counter_n2, 
      dp_id_stage_regfile_DataPath_CANRESTORE_counter_n8, 
      dp_id_stage_regfile_DataPath_CANRESTORE_counter_n7, 
      dp_id_stage_regfile_DataPath_CANRESTORE_counter_n6, 
      dp_id_stage_regfile_DataPath_CANRESTORE_counter_n4, 
      dp_id_stage_regfile_DataPath_CANRESTORE_counter_n2, 
      dp_id_stage_regfile_DataPath_Mux_rd_n1, 
      dp_id_stage_regfile_DataPath_Mux_rd_n13, 
      dp_id_stage_regfile_DataPath_Mux_rd_n12, 
      dp_id_stage_regfile_DataPath_Mux_rd_n11, 
      dp_id_stage_regfile_DataPath_Mux_rd_n10, 
      dp_id_stage_regfile_DataPath_Mux_rd_n9, 
      dp_id_stage_regfile_DataPath_Mux_rd_n8, 
      dp_id_stage_regfile_DataPath_Mux_wr_n7, 
      dp_id_stage_regfile_DataPath_Mux_wr_n6, 
      dp_id_stage_regfile_DataPath_Mux_wr_n5, 
      dp_id_stage_regfile_DataPath_Mux_wr_n4, 
      dp_id_stage_regfile_DataPath_Mux_wr_n3, 
      dp_id_stage_regfile_DataPath_Mux_wr_n2, 
      dp_id_stage_regfile_DataPath_Mux_wr_n1, 
      dp_id_stage_regfile_DataPath_Mux_sf_n1, 
      dp_id_stage_regfile_DataPath_Mux_sf_n3, 
      dp_id_stage_regfile_DataPath_Mux_rd1_control_n2, 
      dp_id_stage_regfile_DataPath_Mux_rd1_control_n3, 
      dp_id_stage_regfile_DataPath_Mux_rd2_control_n4, 
      dp_id_stage_regfile_DataPath_Mux_rd2_control_n2, 
      dp_id_stage_regfile_DataPath_Mux_wr_control_n4, 
      dp_id_stage_regfile_DataPath_Mux_wr_control_n2, 
      dp_id_stage_regfile_DataPath_Mux_en_control_n4, 
      dp_id_stage_regfile_DataPath_Mux_en_control_n2, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4270, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4269, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4268, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4267, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4266, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4265, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4264, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4263, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4262, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4261, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4260, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4259, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4258, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4257, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4256, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4255, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4254, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4253, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4252, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4251, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4250, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4249, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4248, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4247, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4246, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4245, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4244, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4243, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4242, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4241, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4240, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4239, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4238, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4237, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4236, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4235, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4234, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4233, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4232, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4231, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4230, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4229, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4228, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4227, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4226, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4225, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4224, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4223, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4222, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4221, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4220, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4219, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4218, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4217, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4216, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4215, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4214, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4213, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4212, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4211, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4210, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4209, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4208, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4207, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4206, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4205, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4204, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4203, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4202, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4201, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4200, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4199, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4198, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4197, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4196, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4195, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4194, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4193, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4192, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4191, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4190, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4189, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4186, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4185, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4184, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4183, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4182, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4181, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4180, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4179, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4178, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4175, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4174, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4173, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4172, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4171, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4170, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4169, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4168, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4167, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4164, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4163, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4162, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4161, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4160, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4159, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4158, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4157, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4156, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4153, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4152, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4151, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4150, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4149, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4148, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4147, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4146, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4145, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4144, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4143, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4142, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4141, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4140, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4139, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4138, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4137, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4136, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4135, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4134, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4133, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4132, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4131, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4130, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4129, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4128, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4127, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4126, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4125, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4124, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4123, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4122, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4121, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4120, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4119, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4118, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4117, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4116, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4115, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4114, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4113, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4112, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4111, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4110, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4109, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4108, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4107, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4106, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4105, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4104, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4103, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4102, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4101, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4100, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4099, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4098, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4097, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4096, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4093, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4092, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4091, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4090, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4089, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4088, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4087, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4086, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4085, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4082, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4081, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4080, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4079, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4078, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4077, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4076, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4075, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4074, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4073, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4072, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4071, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4070, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4069, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4068, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4067, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4066, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4065, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4064, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4063, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4062, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4061, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4060, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4059, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4058, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4057, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4056, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4053, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4052, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4051, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4050, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4049, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4048, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4047, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4046, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4045, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4042, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4041, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4040, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4039, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4038, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4037, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4036, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4035, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4034, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4033, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4032, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4031, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4030, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4029, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4028, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4027, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4026, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4025, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4024, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4023, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4022, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4021, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4020, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4019, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4018, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4017, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4016, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4015, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4014, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4013, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4012, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4011, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4010, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4009, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4008, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4007, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4006, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4005, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4002, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4001, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4000, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3999, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3998, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3997, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3996, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3995, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3994, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3991, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3990, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3989, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3988, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3987, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3986, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3985, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3984, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3983, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3982, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3981, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3980, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3979, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3978, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3977, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3976, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3975, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3974, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3973, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3972, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3971, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3970, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3969, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3968, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3967, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3966, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3965, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3964, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3961, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3960, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3959, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3958, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3957, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3956, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3955, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3954, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3953, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3950, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3949, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3948, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3947, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3946, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3945, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3944, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3943, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3942, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3941, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3940, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3939, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3938, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3937, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3936, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3935, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3934, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3933, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3932, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3931, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3930, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3929, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3928, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3927, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3926, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3925, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3924, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3923, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3922, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3921, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3920, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3919, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3918, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3917, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3916, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3915, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3914, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3911, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3910, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3909, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3908, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3907, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3906, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3905, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3904, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3903, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3900, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3899, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3898, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3897, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3896, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3895, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3894, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3893, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3892, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3891, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3890, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3889, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3888, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3887, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3886, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3885, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3884, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3883, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3882, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3881, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3880, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3879, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3878, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3877, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3876, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3875, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3874, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3873, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3872, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3869, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3868, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3867, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3866, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3865, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3864, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3863, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3862, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3861, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3858, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3857, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3856, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3855, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3854, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3853, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3852, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3851, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3850, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3849, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3848, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3847, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3846, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3845, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3844, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3843, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3842, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3841, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3840, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3839, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3838, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3837, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3836, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3835, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3834, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3833, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3832, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3831, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3830, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3829, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3828, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3827, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3826, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3825, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3824, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3823, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3822, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3821, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3820, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3816, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3815, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3814, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3813, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3812, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3811, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3810, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3809, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3808, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3807, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3806, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3805, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3804, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3803, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3802, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3801, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3800, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3799, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3798, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3797, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3796, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3795, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3794, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3793, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3792, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3791, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3790, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3789, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3788, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3787, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3786, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3785, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3784, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3783, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3782, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3781, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3780, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3779, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3778, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3777, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3776, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3775, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3774, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3773, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3772, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3771, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3770, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3769, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3768, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3767, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3766, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3765, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3764, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3763, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3762, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3761, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3760, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3759, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3758, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3757, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3756, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3755, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3754, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3753, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3752, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3751, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3750, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3749, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3748, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3747, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3746, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3745, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3744, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3743, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3742, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3741, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3740, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3739, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3738, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3737, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3736, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3735, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3734, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3733, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3732, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3731, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3730, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3729, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3728, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3727, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3726, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3725, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3724, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3723, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3722, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3721, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3720, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3719, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3718, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3717, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3716, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3715, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3714, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3713, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3712, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3708, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3707, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3706, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3705, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3704, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3703, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3702, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3701, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3700, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3699, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3698, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3697, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3696, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3695, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3694, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3693, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1926, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1925, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1858, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1857, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1756, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1755, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1688, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1687, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1586, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1585, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1518, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1516, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1348, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1346, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1343, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1340, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1236, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1235, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1234, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1233, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1232, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1231, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1230, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1229, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1228, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1227, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1226, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1225, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1224, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1223, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1222, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1221, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1220, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1219, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1218, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1217, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1216, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1215, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1214, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1213, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1212, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1211, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1210, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1209, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1208, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1207, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1206, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1205, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1204, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1203, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1202, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1200, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1189, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1188, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1187, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1186, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1185, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1184, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1183, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1182, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1181, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1180, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1179, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1178, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1177, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1176, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1175, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1174, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1173, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1172, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1171, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1170, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1169, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1168, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1167, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1166, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1165, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1164, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1163, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1162, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1161, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1160, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1159, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1158, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1157, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1156, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1155, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1154, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3692, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3691, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3690, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3689, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3688, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3687, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3686, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3685, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3684, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3683, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3682, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3681, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3680, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3679, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3678, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3677, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3676, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3675, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3674, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3673, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3672, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3671, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3670, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3669, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3668, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3667, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3666, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3665, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3664, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3663, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3662, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3661, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3660, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3659, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3658, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3657, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3656, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3655, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3654, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3653, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3652, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3651, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3650, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3649, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3648, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3647, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3646, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3645, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3644, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3643, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3642, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3641, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3640, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3639, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3638, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3637, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3636, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3635, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3634, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3633, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3632, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3631, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3630, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3629, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3628, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3627, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3626, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3625, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3624, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3623, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3622, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3621, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3620, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3619, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3618, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3617, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3616, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3615, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3614, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3613, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3612, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3611, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3610, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3609, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3608, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3607, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3606, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3605, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3604, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3603, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3602, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3601, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3600, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3599, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3598, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3597, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3596, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3595, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3594, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3593, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3592, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3591, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3590, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3589, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3588, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3587, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3586, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3585, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3584, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3583, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3582, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3581, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3580, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3579, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3578, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3577, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3576, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3575, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3574, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3573, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3572, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3571, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3570, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3569, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3568, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3567, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3566, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3565, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3564, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3563, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3562, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3561, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3560, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3559, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3558, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3557, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3556, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3555, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3554, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3553, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3552, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3551, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3550, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3549, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3548, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3547, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3546, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3545, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3544, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3543, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3542, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3541, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3540, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3539, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3538, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3537, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3536, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3535, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3534, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3533, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3532, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3531, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3530, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3529, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3528, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3527, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3526, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3525, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3524, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3523, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3522, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3521, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3520, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3519, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3518, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3517, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3516, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3515, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3514, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3513, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3512, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3511, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3510, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3509, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3508, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3507, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3506, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3505, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3504, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3503, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3502, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3501, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3500, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3499, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3498, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3497, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3496, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3495, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3494, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3493, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3492, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3491, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3490, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3489, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3488, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3487, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3486, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3485, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3484, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3483, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3482, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3481, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3480, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3479, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3478, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3477, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3476, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3475, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3474, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3473, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3472, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3471, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3470, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3469, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3468, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3467, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3466, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3465, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3464, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3463, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3462, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3461, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3460, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3459, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3458, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3457, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3456, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3455, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3454, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3453, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3452, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3451, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3450, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3449, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3448, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3447, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3446, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3445, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3444, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3443, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3442, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3441, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3440, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3439, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3438, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3437, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3436, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3435, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3434, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3433, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3432, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3431, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3430, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3429, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3428, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3427, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3426, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3425, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3424, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3423, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3422, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3421, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3420, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3419, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3418, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3417, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3416, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3415, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3414, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3413, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3412, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3411, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3410, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3409, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3408, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3407, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3406, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3405, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3404, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3403, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3402, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3401, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3400, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3399, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3398, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3397, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3396, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3395, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3394, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3393, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3392, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3391, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3390, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3389, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3388, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3387, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3386, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3385, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3384, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3383, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3382, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3381, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3380, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3379, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3378, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3377, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3376, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3375, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3374, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3373, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3372, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3371, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3370, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3369, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3368, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3367, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3366, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3365, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3364, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3363, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3362, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3361, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3360, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3359, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3358, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3357, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3356, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3355, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3354, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3353, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3352, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3351, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3350, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3349, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3348, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3347, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3346, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3345, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3344, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3343, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3342, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3341, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3340, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3339, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3338, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3337, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3336, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3335, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3334, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3333, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3332, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3331, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3330, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3329, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3328, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3327, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3326, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3325, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3324, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3323, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3322, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3321, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3320, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3319, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3318, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3317, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3316, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3315, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3314, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3313, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3312, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3311, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3310, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3309, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3308, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3307, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3306, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3305, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3304, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3303, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3302, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3301, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3300, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3299, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3298, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3297, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3296, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3295, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3294, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3293, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3292, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3291, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3290, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3289, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3288, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3287, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3286, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3285, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3284, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3283, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3282, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3281, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3280, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3279, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3278, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3277, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3276, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3275, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3274, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3273, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3272, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3271, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3270, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3269, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3268, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3267, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3266, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3265, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3264, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3263, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3262, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3261, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3260, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3259, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3258, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3257, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3256, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3255, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3254, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3253, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3252, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3251, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3250, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3249, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3248, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3247, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3246, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3245, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3244, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3243, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3242, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3241, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3240, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3239, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3238, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3237, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3236, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3235, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3234, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3233, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3232, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3231, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3230, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3229, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3228, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3227, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3226, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3225, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3224, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3223, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3222, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3221, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3220, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3219, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3218, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3217, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3216, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3215, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3214, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3213, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3212, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3211, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3210, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3209, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3208, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3207, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3206, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3205, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3204, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3203, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3202, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3201, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3200, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3199, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3198, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3197, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3196, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3195, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3194, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3193, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3192, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3191, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3190, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3189, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3188, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3187, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3186, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3185, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3184, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3183, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3182, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3181, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3180, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3179, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3178, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3177, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3176, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3175, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3174, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3173, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3172, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3171, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3170, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3169, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3168, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3167, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3166, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3165, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3164, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3163, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3162, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3161, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3158, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3155, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3154, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3153, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3152, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3151, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3150, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3149, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3148, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3147, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3146, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3145, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3144, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3143, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3142, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3141, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3140, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3139, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3138, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3137, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3136, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3135, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3134, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3133, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3132, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3131, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3130, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3129, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3128, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3127, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3126, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3125, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3124, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3123, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3122, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3121, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3120, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3119, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3118, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3117, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3116, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3115, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3114, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3113, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3112, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3111, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3110, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3109, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3108, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3107, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3106, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3105, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3104, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3103, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3102, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3101, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3100, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3099, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3098, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3097, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3096, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3095, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3094, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3093, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3092, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3091, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3090, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3089, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3088, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3087, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3086, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3085, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3084, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3083, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3082, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3081, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3080, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3079, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3078, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3077, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3076, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3075, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3074, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3073, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3072, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3071, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3070, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3069, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3068, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3067, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3066, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3065, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3064, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3063, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3062, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3061, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3060, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3059, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3058, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3057, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3056, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3055, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3054, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3053, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3052, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3051, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3050, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3049, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3048, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3047, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3046, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3045, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3044, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3043, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3042, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3041, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3040, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3039, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3038, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3037, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3036, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3035, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3034, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3033, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3032, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3031, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3030, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3029, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3028, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3027, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3026, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3025, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3024, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3023, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3022, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3021, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3020, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3019, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3018, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3017, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3016, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3015, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3014, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3013, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3012, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3011, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3010, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3009, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3008, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3007, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3006, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3005, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3004, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3003, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3002, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3001, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3000, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2999, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2998, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2997, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2996, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2995, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2994, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2993, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2992, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2991, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2990, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2989, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2988, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2987, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2986, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2985, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2984, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2983, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2982, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2981, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2980, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2979, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2978, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2977, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2976, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2975, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2974, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2973, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2972, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2971, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2970, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2969, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2968, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2967, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2966, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2965, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2964, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2963, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2962, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2961, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2960, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2959, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2958, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2957, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2956, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2955, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2954, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2953, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2952, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2951, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2950, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2949, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2948, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2947, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2946, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2945, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2944, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2943, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2942, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2941, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2940, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2939, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2938, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2937, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2936, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2935, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2934, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2933, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2932, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2931, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2930, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2929, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2928, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2927, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2926, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2925, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2924, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2923, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2922, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2921, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2920, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2919, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2918, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2917, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2916, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2915, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2914, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2913, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2912, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2911, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2910, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2909, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2908, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2907, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2906, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2905, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2904, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2903, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2902, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2901, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2900, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2899, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2898, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2897, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2896, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2895, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2894, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2893, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2892, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2891, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2890, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2889, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2888, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2887, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2886, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2885, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2884, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2883, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2882, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2881, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2880, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2879, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2878, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2877, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2876, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2875, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2874, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2873, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2872, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2871, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2870, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2869, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2868, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2867, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2866, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2865, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2864, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2863, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2862, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2861, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2860, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2859, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2858, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2857, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2856, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2855, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2854, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2853, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2852, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2851, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2850, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2849, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2848, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2847, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2846, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2845, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2844, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2843, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2842, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2841, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2840, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2839, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2838, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2837, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2836, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2835, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2834, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2833, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2832, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2831, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2830, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2829, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2828, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2827, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2826, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2825, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2824, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2823, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2822, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2821, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2820, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2819, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2818, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2817, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2816, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2815, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2814, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2813, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2812, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2811, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2810, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2809, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2808, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2807, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2806, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2805, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2804, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2803, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2802, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2801, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2800, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2799, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2798, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2797, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2796, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2795, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2794, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2793, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2792, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2791, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2790, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2789, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2788, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2787, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2786, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2785, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2784, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2783, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2782, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2781, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2780, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2779, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2778, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2777, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2776, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2775, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2774, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2773, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2772, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2771, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2770, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2769, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2768, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2767, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2766, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2765, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2764, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2763, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2762, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2761, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2760, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2759, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2758, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2757, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2756, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2755, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2754, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2753, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2752, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2751, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2750, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2749, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2748, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2747, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2746, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2745, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2744, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2743, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2742, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2741, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2740, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2739, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2738, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2737, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2736, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2735, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2734, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2733, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2732, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2731, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2730, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2729, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2728, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2727, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2726, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2725, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2724, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2723, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2722, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2721, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2720, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2719, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2718, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2717, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2716, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2715, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2714, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2713, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2712, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2711, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2710, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2709, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2708, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2707, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2706, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2705, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2704, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2703, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2702, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2701, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2700, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2699, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2698, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2697, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2696, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2695, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2694, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2693, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2692, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2691, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2690, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2689, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2688, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2687, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2686, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2685, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2684, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2683, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2682, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2681, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2680, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2679, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2678, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2677, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2676, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2675, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2674, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2673, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2672, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2671, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2670, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2669, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2668, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2667, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2666, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2665, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2664, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2663, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2662, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2661, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2660, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2659, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2658, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2657, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2656, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2655, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2654, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2653, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2652, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2651, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2650, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2649, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2648, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2647, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2646, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2645, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2644, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2643, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2642, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2641, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2640, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2639, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2638, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2637, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2636, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2635, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2634, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2633, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2632, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2631, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2630, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2629, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2628, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2627, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2626, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2625, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2624, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2623, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2622, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2621, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2620, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2619, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2618, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2617, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2616, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2615, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2614, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2613, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2612, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2611, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2610, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2609, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2608, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2607, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2606, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2605, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2604, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2603, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2602, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2601, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2600, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2599, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2598, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2597, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2596, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2595, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2594, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2593, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2592, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2591, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2590, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2589, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2588, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2587, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2586, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2585, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2584, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2583, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2582, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2581, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2580, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2579, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2578, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2577, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2576, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2575, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2574, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2573, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2572, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2571, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2570, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2569, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2568, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2567, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2566, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2565, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2564, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2563, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2562, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2561, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2560, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2559, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2558, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2557, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2556, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2555, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2554, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2553, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2552, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2551, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2550, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2549, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2548, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2547, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2546, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2545, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2544, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2543, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2542, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2541, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2540, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2539, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2538, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2537, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2536, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2535, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2534, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2531, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2528, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2527, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2526, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2525, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2524, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2523, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2522, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2521, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2520, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2519, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2518, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2517, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2516, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2515, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2514, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2513, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2512, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2511, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2510, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2509, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2508, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2507, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2506, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2505, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2504, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2503, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2502, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2501, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2500, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2499, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2498, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2497, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2496, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2495, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2494, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2493, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2492, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2491, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2490, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2489, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2488, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2487, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2486, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2485, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2484, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2483, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2482, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2481, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2480, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2479, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2478, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2477, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2476, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2475, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2474, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2473, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2472, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2471, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2470, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2469, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2468, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2467, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2466, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2465, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2464, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2463, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2462, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2461, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2460, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2459, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2458, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2457, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2456, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2455, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2454, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2453, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2452, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2451, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2450, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2449, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2448, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2447, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2446, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2445, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2444, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2443, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2442, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2441, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2440, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2439, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2438, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2437, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2436, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2435, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2434, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2433, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2432, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2431, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2430, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2429, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2428, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2427, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2426, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2425, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2424, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2423, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2422, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2421, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2420, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2419, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2418, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2417, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2416, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2415, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2414, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2413, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2412, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2411, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2410, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2409, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2408, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2407, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2406, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2405, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2404, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2403, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2402, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2401, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2400, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2399, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2398, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2397, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2396, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2395, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2394, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2393, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2392, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2391, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2390, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2389, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2388, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2387, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2386, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2385, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2384, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2383, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2382, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2381, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2380, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2379, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2378, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2377, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2376, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2375, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2374, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2373, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2372, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2371, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2370, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2369, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2368, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2367, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2366, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2365, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2364, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2363, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2362, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2361, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2360, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2359, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2358, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2357, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2356, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2355, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2354, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2353, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2352, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2351, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2350, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2349, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2348, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2347, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2346, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2345, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2344, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2343, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2342, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2341, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2340, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2339, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2338, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2337, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2336, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2335, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2334, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2333, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2332, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2331, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2330, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2329, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2328, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2327, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2326, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2325, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2324, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2323, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2322, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2321, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2320, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2319, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2318, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2317, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2316, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2315, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2314, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2313, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2312, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2311, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2310, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2309, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2308, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2307, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2306, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2305, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2304, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2303, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2302, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2301, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2300, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2299, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2298, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2297, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2296, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2295, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2294, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2293, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2292, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2291, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2290, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2289, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2288, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2287, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2286, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2285, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2284, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2283, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2282, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2281, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2280, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2279, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2278, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2277, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2276, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2275, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2274, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2273, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2272, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2271, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2270, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2269, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2268, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2267, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2266, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2265, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2264, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2263, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2262, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2261, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2260, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2259, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2258, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2257, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2256, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2255, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2254, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2253, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2252, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2251, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2250, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2249, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2248, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2247, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2246, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2245, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2244, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2243, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2242, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2241, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2240, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2239, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2238, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2237, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2236, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2235, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2234, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2233, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2232, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2231, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2230, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2229, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2228, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2227, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2226, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2225, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2224, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2223, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2222, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2221, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2220, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2219, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2218, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2217, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2216, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2215, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2214, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2213, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2212, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2211, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2210, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2209, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2208, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2207, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2206, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2205, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2204, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2203, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2202, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2201, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2200, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2199, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2198, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2197, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2196, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2195, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2194, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2193, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2192, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2191, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2190, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2189, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2188, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2187, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2186, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2185, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2184, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2183, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2182, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2181, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2180, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2179, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2178, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2177, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2176, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2175, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2174, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2173, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2172, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2171, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2170, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2169, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2168, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2167, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2166, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2165, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2164, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2163, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2162, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2161, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2160, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2159, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2158, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2157, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2156, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2155, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2154, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2153, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2152, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2151, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2150, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2149, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2148, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2147, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2146, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2145, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2144, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2143, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2142, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2141, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2140, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2139, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2138, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2137, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2136, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2135, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2134, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2133, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2132, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2131, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2130, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2129, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2128, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2127, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2126, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2125, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2124, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2123, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2122, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2121, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2120, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2119, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2118, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2117, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2116, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2115, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2114, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2113, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2112, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2111, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2110, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2109, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2108, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2107, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2106, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2105, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2104, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2103, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2102, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2101, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2100, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2099, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2098, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2097, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2096, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2095, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2094, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2093, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2092, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2091, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2090, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2089, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2088, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2087, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2086, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2085, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2084, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2083, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2082, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2081, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2080, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2079, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2078, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2077, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2076, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2075, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2074, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2073, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2072, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2071, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2070, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2069, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2068, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2067, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2066, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2065, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2064, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2063, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2062, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2061, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2060, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2059, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2058, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2057, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2056, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2055, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2054, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2053, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2052, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2051, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2050, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2049, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2048, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2047, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2046, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2045, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2044, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2043, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2042, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2041, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2040, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2039, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2038, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2037, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2036, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2035, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2034, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2033, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2032, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2031, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2030, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2029, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2028, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2027, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2026, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2025, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2024, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2023, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2022, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2021, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2020, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2019, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2018, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2017, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2016, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2015, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2014, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2013, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2012, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2011, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2010, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2009, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2008, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2007, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2006, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2005, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2004, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2003, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2002, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2001, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2000, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1999, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1998, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1997, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1996, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1995, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1994, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1993, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1992, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1991, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1990, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1989, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1988, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1987, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1986, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1985, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1984, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1983, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1982, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1981, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1980, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1979, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1978, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1977, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1976, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1975, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1974, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1973, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1972, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1971, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1970, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1969, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1968, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1967, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1966, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1965, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1964, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1963, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1962, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1961, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1960, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1959, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1958, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1957, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1956, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1955, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1954, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1953, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1952, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1951, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1950, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1949, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1948, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1947, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1946, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1945, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1944, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1943, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1942, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1941, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1940, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1939, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1938, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1937, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1936, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1935, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1934, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1933, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1932, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1931, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1930, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1929, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1928, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1927, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1924, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1923, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1922, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1921, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1920, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1919, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1918, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1917, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1916, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1915, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1914, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1913, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1912, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1911, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1910, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1909, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1908, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1907, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1906, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1905, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1904, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1903, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1902, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1901, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1900, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1899, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1898, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1897, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1896, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1895, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1894, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1893, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1892, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1891, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1890, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1889, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1888, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1887, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1886, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1885, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1884, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1883, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1882, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1881, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1880, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1879, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1878, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1877, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1876, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1875, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1874, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1873, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1872, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1871, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1870, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1869, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1868, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1867, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1866, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1865, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1864, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1863, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1862, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1861, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1860, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1859, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1856, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1855, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1854, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1853, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1852, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1851, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1850, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1849, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1848, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1847, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1846, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1845, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1844, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1843, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1842, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1841, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1840, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1839, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1838, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1837, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1836, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1835, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1834, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1833, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1832, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1831, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1830, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1829, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1828, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1827, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1826, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1825, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1824, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1823, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1822, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1821, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1820, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1819, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1818, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1817, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1816, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1815, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1814, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1813, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1812, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1811, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1810, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1809, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1808, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1807, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1806, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1805, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1804, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1803, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1802, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1801, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1800, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1799, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1798, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1797, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1796, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1795, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1794, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1793, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1792, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1791, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1790, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1789, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1788, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1787, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1786, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1785, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1784, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1783, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1782, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1781, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1780, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1779, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1778, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1777, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1776, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1775, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1774, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1773, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1772, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1771, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1770, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1769, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1768, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1767, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1766, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1765, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1764, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1763, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1762, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1761, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1760, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1759, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1758, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1757, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1754, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1753, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1752, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1751, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1750, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1749, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1748, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1747, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1746, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1745, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1744, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1743, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1742, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1741, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1740, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1739, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1738, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1737, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1736, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1735, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1734, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1733, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1732, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1731, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1730, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1729, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1728, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1727, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1726, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1725, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1724, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1723, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1722, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1721, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1720, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1719, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1718, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1717, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1716, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1715, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1714, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1713, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1712, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1711, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1710, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1709, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1708, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1707, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1706, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1705, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1704, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1703, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1702, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1701, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1700, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1699, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1698, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1697, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1696, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1695, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1694, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1693, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1692, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1691, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1690, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1689, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1686, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1685, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1684, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1683, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1682, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1681, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1680, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1679, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1678, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1677, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1676, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1675, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1674, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1673, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1672, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1671, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1670, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1669, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1668, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1667, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1666, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1665, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1664, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1663, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1662, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1661, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1660, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1659, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1658, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1657, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1656, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1655, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1654, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1653, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1652, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1651, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1650, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1649, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1648, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1647, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1646, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1645, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1644, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1643, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1642, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1641, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1640, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1639, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1638, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1637, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1636, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1635, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1634, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1633, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1632, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1631, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1630, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1629, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1628, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1627, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1626, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1625, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1624, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1623, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1622, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1621, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1620, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1619, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1618, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1617, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1616, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1615, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1614, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1613, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1612, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1611, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1610, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1609, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1608, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1607, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1606, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1605, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1604, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1603, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1602, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1601, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1600, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1599, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1598, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1597, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1596, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1595, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1594, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1593, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1592, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1591, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1590, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1589, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1588, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1587, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1584, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1583, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1582, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1581, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1580, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1579, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1578, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1577, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1576, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1575, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1574, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1573, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1572, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1571, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1570, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1569, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1568, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1567, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1566, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1565, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1564, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1563, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1562, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1561, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1560, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1559, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1558, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1557, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1556, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1555, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1554, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1553, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1552, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1551, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1550, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1549, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1548, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1547, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1546, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1545, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1544, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1543, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1542, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1541, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1540, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1539, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1538, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1537, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1536, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1535, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1534, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1533, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1532, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1531, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1530, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1529, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1528, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1527, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1526, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1525, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1524, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1523, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1522, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1521, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1520, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1519, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1517, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1515, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1514, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1513, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1512, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1511, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1510, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1509, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1508, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1507, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1506, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1505, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1504, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1503, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1502, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1501, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1500, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1499, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1498, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1497, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1496, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1495, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1494, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1493, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1492, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1491, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1490, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1489, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1488, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1487, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1486, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1485, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1484, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1483, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1482, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1481, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1480, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1479, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1478, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1477, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1476, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1475, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1474, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1473, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1472, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1471, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1470, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1469, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1468, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1467, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1466, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1465, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1464, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1463, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1462, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1461, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1460, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1459, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1458, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1457, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1456, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1455, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1454, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1453, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1452, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1451, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1450, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1449, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1448, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1447, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1446, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1445, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1444, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1443, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1442, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1441, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1440, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1439, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1438, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1437, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1436, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1435, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1434, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1433, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1432, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1431, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1430, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1429, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1428, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1427, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1426, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1425, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1424, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1423, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1422, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1421, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1420, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1419, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1418, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1417, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1416, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1415, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1414, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1413, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1412, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1411, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1410, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1409, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1408, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1407, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1406, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1405, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1404, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1403, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1402, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1401, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1400, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1399, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1398, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1397, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1396, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1395, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1394, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1393, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1392, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1391, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1390, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1389, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1388, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1387, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1386, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1385, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1384, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1383, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1382, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1381, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1380, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1379, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1378, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1377, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1376, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1375, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1374, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1373, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1372, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1371, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1370, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1369, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1368, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1367, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1366, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1365, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1364, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1363, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1362, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1361, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1360, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1359, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1358, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1357, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1356, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1355, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1354, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1353, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1352, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1351, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1350, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1349, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1347, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1345, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1344, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1342, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1341, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1339, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1338, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1337, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1336, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1335, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1334, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1333, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1332, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1331, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1330, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1329, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1328, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1327, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1326, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1325, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1324, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1323, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1322, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1321, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1320, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1319, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1318, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1317, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1316, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1315, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1314, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1313, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1312, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1311, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1310, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1309, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1308, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1307, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1306, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1305, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1304, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1303, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1302, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1301, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1300, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1299, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1298, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1297, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1296, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1295, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1294, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1293, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1292, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1291, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1290, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1289, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1288, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1287, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1286, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1285, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1284, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1283, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1282, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1281, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1280, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1279, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1278, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1277, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1276, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1275, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1274, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1273, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1272, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1271, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1270, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1269, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1268, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1267, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1266, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1265, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1264, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1263, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1262, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1261, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1260, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1259, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1258, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1257, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1256, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1255, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1254, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1253, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1252, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1251, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1250, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1249, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1248, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1247, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1246, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1245, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1244, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1243, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1242, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1241, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1240, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1239, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1238, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1237, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1201, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1199, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1198, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1197, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1196, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1195, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1194, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1193, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1192, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1191, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1190, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1153, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1152, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1151, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1150, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1149, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1148, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1147, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1146, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1145, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1144, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1143, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1142, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1141, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1140, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1139, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1138, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1137, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1136, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1135, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1134, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1133, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1132, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1131, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1130, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1129, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1128, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1127, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1126, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1125, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1124, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1123, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1122, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1121, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1120, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1119, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1118, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1117, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1116, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1115, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1114, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1113, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1112, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1111, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1110, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1109, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1108, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1107, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1106, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1105, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1104, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1103, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1102, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1101, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1100, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1099, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1098, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1097, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1096, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1095, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1094, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1093, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1092, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1091, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1090, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1089, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1088, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1087, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1086, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1085, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1084, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1083, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1082, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1081, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1080, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1079, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1078, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1077, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1076, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1075, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1074, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1073, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1072, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1071, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1070, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1069, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1068, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1067, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1066, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1065, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1064, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1063, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1062, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1061, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1060, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1059, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1058, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1057, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1056, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1055, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1054, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1053, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1052, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1051, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1050, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1049, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1048, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1047, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1046, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1045, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1044, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1043, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1042, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1041, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1040, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1039, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1038, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1037, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1036, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1035, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1034, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1033, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1032, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1031, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1030, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1029, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1028, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1027, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1026, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1025, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1024, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1023, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1022, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1021, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1020, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1019, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1018, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1017, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1016, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1015, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1014, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1013, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1012, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1011, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1010, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1009, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1008, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1007, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1006, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1005, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1004, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1003, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1002, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1001, 
      dp_id_stage_regfile_DataPath_Physical_RF_n1000, 
      dp_id_stage_regfile_DataPath_Physical_RF_n999, 
      dp_id_stage_regfile_DataPath_Physical_RF_n998, 
      dp_id_stage_regfile_DataPath_Physical_RF_n997, 
      dp_id_stage_regfile_DataPath_Physical_RF_n996, 
      dp_id_stage_regfile_DataPath_Physical_RF_n995, 
      dp_id_stage_regfile_DataPath_Physical_RF_n994, 
      dp_id_stage_regfile_DataPath_Physical_RF_n993, 
      dp_id_stage_regfile_DataPath_Physical_RF_n992, 
      dp_id_stage_regfile_DataPath_Physical_RF_n991, 
      dp_id_stage_regfile_DataPath_Physical_RF_n990, 
      dp_id_stage_regfile_DataPath_Physical_RF_n989, 
      dp_id_stage_regfile_DataPath_Physical_RF_n988, 
      dp_id_stage_regfile_DataPath_Physical_RF_n987, 
      dp_id_stage_regfile_DataPath_Physical_RF_n986, 
      dp_id_stage_regfile_DataPath_Physical_RF_n985, 
      dp_id_stage_regfile_DataPath_Physical_RF_n984, 
      dp_id_stage_regfile_DataPath_Physical_RF_n983, 
      dp_id_stage_regfile_DataPath_Physical_RF_n982, 
      dp_id_stage_regfile_DataPath_Physical_RF_n981, 
      dp_id_stage_regfile_DataPath_Physical_RF_n980, 
      dp_id_stage_regfile_DataPath_Physical_RF_n979, 
      dp_id_stage_regfile_DataPath_Physical_RF_n978, 
      dp_id_stage_regfile_DataPath_Physical_RF_n977, 
      dp_id_stage_regfile_DataPath_Physical_RF_n976, 
      dp_id_stage_regfile_DataPath_Physical_RF_n975, 
      dp_id_stage_regfile_DataPath_Physical_RF_n974, 
      dp_id_stage_regfile_DataPath_Physical_RF_n973, 
      dp_id_stage_regfile_DataPath_Physical_RF_n972, 
      dp_id_stage_regfile_DataPath_Physical_RF_n971, 
      dp_id_stage_regfile_DataPath_Physical_RF_n970, 
      dp_id_stage_regfile_DataPath_Physical_RF_n969, 
      dp_id_stage_regfile_DataPath_Physical_RF_n968, 
      dp_id_stage_regfile_DataPath_Physical_RF_n967, 
      dp_id_stage_regfile_DataPath_Physical_RF_n966, 
      dp_id_stage_regfile_DataPath_Physical_RF_n965, 
      dp_id_stage_regfile_DataPath_Physical_RF_n964, 
      dp_id_stage_regfile_DataPath_Physical_RF_n963, 
      dp_id_stage_regfile_DataPath_Physical_RF_n962, 
      dp_id_stage_regfile_DataPath_Physical_RF_n961, 
      dp_id_stage_regfile_DataPath_Physical_RF_n960, 
      dp_id_stage_regfile_DataPath_Physical_RF_n959, 
      dp_id_stage_regfile_DataPath_Physical_RF_n958, 
      dp_id_stage_regfile_DataPath_Physical_RF_n957, 
      dp_id_stage_regfile_DataPath_Physical_RF_n956, 
      dp_id_stage_regfile_DataPath_Physical_RF_n955, 
      dp_id_stage_regfile_DataPath_Physical_RF_n954, 
      dp_id_stage_regfile_DataPath_Physical_RF_n953, 
      dp_id_stage_regfile_DataPath_Physical_RF_n952, 
      dp_id_stage_regfile_DataPath_Physical_RF_n951, 
      dp_id_stage_regfile_DataPath_Physical_RF_n950, 
      dp_id_stage_regfile_DataPath_Physical_RF_n949, 
      dp_id_stage_regfile_DataPath_Physical_RF_n948, 
      dp_id_stage_regfile_DataPath_Physical_RF_n947, 
      dp_id_stage_regfile_DataPath_Physical_RF_n946, 
      dp_id_stage_regfile_DataPath_Physical_RF_n945, 
      dp_id_stage_regfile_DataPath_Physical_RF_n944, 
      dp_id_stage_regfile_DataPath_Physical_RF_n943, 
      dp_id_stage_regfile_DataPath_Physical_RF_n942, 
      dp_id_stage_regfile_DataPath_Physical_RF_n941, 
      dp_id_stage_regfile_DataPath_Physical_RF_n940, 
      dp_id_stage_regfile_DataPath_Physical_RF_n939, 
      dp_id_stage_regfile_DataPath_Physical_RF_n938, 
      dp_id_stage_regfile_DataPath_Physical_RF_n937, 
      dp_id_stage_regfile_DataPath_Physical_RF_n936, 
      dp_id_stage_regfile_DataPath_Physical_RF_n935, 
      dp_id_stage_regfile_DataPath_Physical_RF_n934, 
      dp_id_stage_regfile_DataPath_Physical_RF_n933, 
      dp_id_stage_regfile_DataPath_Physical_RF_n932, 
      dp_id_stage_regfile_DataPath_Physical_RF_n931, 
      dp_id_stage_regfile_DataPath_Physical_RF_n930, 
      dp_id_stage_regfile_DataPath_Physical_RF_n929, 
      dp_id_stage_regfile_DataPath_Physical_RF_n928, 
      dp_id_stage_regfile_DataPath_Physical_RF_n927, 
      dp_id_stage_regfile_DataPath_Physical_RF_n926, 
      dp_id_stage_regfile_DataPath_Physical_RF_n925, 
      dp_id_stage_regfile_DataPath_Physical_RF_n924, 
      dp_id_stage_regfile_DataPath_Physical_RF_n923, 
      dp_id_stage_regfile_DataPath_Physical_RF_n922, 
      dp_id_stage_regfile_DataPath_Physical_RF_n921, 
      dp_id_stage_regfile_DataPath_Physical_RF_n920, 
      dp_id_stage_regfile_DataPath_Physical_RF_n919, 
      dp_id_stage_regfile_DataPath_Physical_RF_n918, 
      dp_id_stage_regfile_DataPath_Physical_RF_n917, 
      dp_id_stage_regfile_DataPath_Physical_RF_n916, 
      dp_id_stage_regfile_DataPath_Physical_RF_n915, 
      dp_id_stage_regfile_DataPath_Physical_RF_n914, 
      dp_id_stage_regfile_DataPath_Physical_RF_n913, 
      dp_id_stage_regfile_DataPath_Physical_RF_n912, 
      dp_id_stage_regfile_DataPath_Physical_RF_n911, 
      dp_id_stage_regfile_DataPath_Physical_RF_n910, 
      dp_id_stage_regfile_DataPath_Physical_RF_n909, 
      dp_id_stage_regfile_DataPath_Physical_RF_n908, 
      dp_id_stage_regfile_DataPath_Physical_RF_n907, 
      dp_id_stage_regfile_DataPath_Physical_RF_n906, 
      dp_id_stage_regfile_DataPath_Physical_RF_n905, 
      dp_id_stage_regfile_DataPath_Physical_RF_n904, 
      dp_id_stage_regfile_DataPath_Physical_RF_n903, 
      dp_id_stage_regfile_DataPath_Physical_RF_n902, 
      dp_id_stage_regfile_DataPath_Physical_RF_n901, 
      dp_id_stage_regfile_DataPath_Physical_RF_n900, 
      dp_id_stage_regfile_DataPath_Physical_RF_n899, 
      dp_id_stage_regfile_DataPath_Physical_RF_n898, 
      dp_id_stage_regfile_DataPath_Physical_RF_n897, 
      dp_id_stage_regfile_DataPath_Physical_RF_n896, 
      dp_id_stage_regfile_DataPath_Physical_RF_n895, 
      dp_id_stage_regfile_DataPath_Physical_RF_n894, 
      dp_id_stage_regfile_DataPath_Physical_RF_n893, 
      dp_id_stage_regfile_DataPath_Physical_RF_n892, 
      dp_id_stage_regfile_DataPath_Physical_RF_n891, 
      dp_id_stage_regfile_DataPath_Physical_RF_n890, 
      dp_id_stage_regfile_DataPath_Physical_RF_n889, 
      dp_id_stage_regfile_DataPath_Physical_RF_n888, 
      dp_id_stage_regfile_DataPath_Physical_RF_n887, 
      dp_id_stage_regfile_DataPath_Physical_RF_n886, 
      dp_id_stage_regfile_DataPath_Physical_RF_n885, 
      dp_id_stage_regfile_DataPath_Physical_RF_n884, 
      dp_id_stage_regfile_DataPath_Physical_RF_n883, 
      dp_id_stage_regfile_DataPath_Physical_RF_n882, 
      dp_id_stage_regfile_DataPath_Physical_RF_n881, 
      dp_id_stage_regfile_DataPath_Physical_RF_n880, 
      dp_id_stage_regfile_DataPath_Physical_RF_n879, 
      dp_id_stage_regfile_DataPath_Physical_RF_n878, 
      dp_id_stage_regfile_DataPath_Physical_RF_n877, 
      dp_id_stage_regfile_DataPath_Physical_RF_n876, 
      dp_id_stage_regfile_DataPath_Physical_RF_n875, 
      dp_id_stage_regfile_DataPath_Physical_RF_n874, 
      dp_id_stage_regfile_DataPath_Physical_RF_n873, 
      dp_id_stage_regfile_DataPath_Physical_RF_n872, 
      dp_id_stage_regfile_DataPath_Physical_RF_n871, 
      dp_id_stage_regfile_DataPath_Physical_RF_n870, 
      dp_id_stage_regfile_DataPath_Physical_RF_n869, 
      dp_id_stage_regfile_DataPath_Physical_RF_n868, 
      dp_id_stage_regfile_DataPath_Physical_RF_n867, 
      dp_id_stage_regfile_DataPath_Physical_RF_n866, 
      dp_id_stage_regfile_DataPath_Physical_RF_n865, 
      dp_id_stage_regfile_DataPath_Physical_RF_n864, 
      dp_id_stage_regfile_DataPath_Physical_RF_n863, 
      dp_id_stage_regfile_DataPath_Physical_RF_n862, 
      dp_id_stage_regfile_DataPath_Physical_RF_n861, 
      dp_id_stage_regfile_DataPath_Physical_RF_n860, 
      dp_id_stage_regfile_DataPath_Physical_RF_n859, 
      dp_id_stage_regfile_DataPath_Physical_RF_n858, 
      dp_id_stage_regfile_DataPath_Physical_RF_n857, 
      dp_id_stage_regfile_DataPath_Physical_RF_n856, 
      dp_id_stage_regfile_DataPath_Physical_RF_n855, 
      dp_id_stage_regfile_DataPath_Physical_RF_n854, 
      dp_id_stage_regfile_DataPath_Physical_RF_n853, 
      dp_id_stage_regfile_DataPath_Physical_RF_n852, 
      dp_id_stage_regfile_DataPath_Physical_RF_n851, 
      dp_id_stage_regfile_DataPath_Physical_RF_n850, 
      dp_id_stage_regfile_DataPath_Physical_RF_n849, 
      dp_id_stage_regfile_DataPath_Physical_RF_n848, 
      dp_id_stage_regfile_DataPath_Physical_RF_n847, 
      dp_id_stage_regfile_DataPath_Physical_RF_n846, 
      dp_id_stage_regfile_DataPath_Physical_RF_n845, 
      dp_id_stage_regfile_DataPath_Physical_RF_n844, 
      dp_id_stage_regfile_DataPath_Physical_RF_n843, 
      dp_id_stage_regfile_DataPath_Physical_RF_n842, 
      dp_id_stage_regfile_DataPath_Physical_RF_n841, 
      dp_id_stage_regfile_DataPath_Physical_RF_n840, 
      dp_id_stage_regfile_DataPath_Physical_RF_n839, 
      dp_id_stage_regfile_DataPath_Physical_RF_n838, 
      dp_id_stage_regfile_DataPath_Physical_RF_n837, 
      dp_id_stage_regfile_DataPath_Physical_RF_n836, 
      dp_id_stage_regfile_DataPath_Physical_RF_n835, 
      dp_id_stage_regfile_DataPath_Physical_RF_n834, 
      dp_id_stage_regfile_DataPath_Physical_RF_n833, 
      dp_id_stage_regfile_DataPath_Physical_RF_n832, 
      dp_id_stage_regfile_DataPath_Physical_RF_n831, 
      dp_id_stage_regfile_DataPath_Physical_RF_n830, 
      dp_id_stage_regfile_DataPath_Physical_RF_n829, 
      dp_id_stage_regfile_DataPath_Physical_RF_n828, 
      dp_id_stage_regfile_DataPath_Physical_RF_n827, 
      dp_id_stage_regfile_DataPath_Physical_RF_n826, 
      dp_id_stage_regfile_DataPath_Physical_RF_n825, 
      dp_id_stage_regfile_DataPath_Physical_RF_n824, 
      dp_id_stage_regfile_DataPath_Physical_RF_n823, 
      dp_id_stage_regfile_DataPath_Physical_RF_n822, 
      dp_id_stage_regfile_DataPath_Physical_RF_n821, 
      dp_id_stage_regfile_DataPath_Physical_RF_n820, 
      dp_id_stage_regfile_DataPath_Physical_RF_n819, 
      dp_id_stage_regfile_DataPath_Physical_RF_n818, 
      dp_id_stage_regfile_DataPath_Physical_RF_n817, 
      dp_id_stage_regfile_DataPath_Physical_RF_n816, 
      dp_id_stage_regfile_DataPath_Physical_RF_n815, 
      dp_id_stage_regfile_DataPath_Physical_RF_n814, 
      dp_id_stage_regfile_DataPath_Physical_RF_n813, 
      dp_id_stage_regfile_DataPath_Physical_RF_n812, 
      dp_id_stage_regfile_DataPath_Physical_RF_n811, 
      dp_id_stage_regfile_DataPath_Physical_RF_n810, 
      dp_id_stage_regfile_DataPath_Physical_RF_n809, 
      dp_id_stage_regfile_DataPath_Physical_RF_n808, 
      dp_id_stage_regfile_DataPath_Physical_RF_n807, 
      dp_id_stage_regfile_DataPath_Physical_RF_n806, 
      dp_id_stage_regfile_DataPath_Physical_RF_n805, 
      dp_id_stage_regfile_DataPath_Physical_RF_n804, 
      dp_id_stage_regfile_DataPath_Physical_RF_n803, 
      dp_id_stage_regfile_DataPath_Physical_RF_n802, 
      dp_id_stage_regfile_DataPath_Physical_RF_n801, 
      dp_id_stage_regfile_DataPath_Physical_RF_n800, 
      dp_id_stage_regfile_DataPath_Physical_RF_n799, 
      dp_id_stage_regfile_DataPath_Physical_RF_n798, 
      dp_id_stage_regfile_DataPath_Physical_RF_n797, 
      dp_id_stage_regfile_DataPath_Physical_RF_n796, 
      dp_id_stage_regfile_DataPath_Physical_RF_n795, 
      dp_id_stage_regfile_DataPath_Physical_RF_n794, 
      dp_id_stage_regfile_DataPath_Physical_RF_n793, 
      dp_id_stage_regfile_DataPath_Physical_RF_n792, 
      dp_id_stage_regfile_DataPath_Physical_RF_n791, 
      dp_id_stage_regfile_DataPath_Physical_RF_n790, 
      dp_id_stage_regfile_DataPath_Physical_RF_n789, 
      dp_id_stage_regfile_DataPath_Physical_RF_n788, 
      dp_id_stage_regfile_DataPath_Physical_RF_n787, 
      dp_id_stage_regfile_DataPath_Physical_RF_n786, 
      dp_id_stage_regfile_DataPath_Physical_RF_n785, 
      dp_id_stage_regfile_DataPath_Physical_RF_n784, 
      dp_id_stage_regfile_DataPath_Physical_RF_n783, 
      dp_id_stage_regfile_DataPath_Physical_RF_n782, 
      dp_id_stage_regfile_DataPath_Physical_RF_n781, 
      dp_id_stage_regfile_DataPath_Physical_RF_n780, 
      dp_id_stage_regfile_DataPath_Physical_RF_n779, 
      dp_id_stage_regfile_DataPath_Physical_RF_n778, 
      dp_id_stage_regfile_DataPath_Physical_RF_n777, 
      dp_id_stage_regfile_DataPath_Physical_RF_n776, 
      dp_id_stage_regfile_DataPath_Physical_RF_n775, 
      dp_id_stage_regfile_DataPath_Physical_RF_n774, 
      dp_id_stage_regfile_DataPath_Physical_RF_n773, 
      dp_id_stage_regfile_DataPath_Physical_RF_n772, 
      dp_id_stage_regfile_DataPath_Physical_RF_n771, 
      dp_id_stage_regfile_DataPath_Physical_RF_n770, 
      dp_id_stage_regfile_DataPath_Physical_RF_n769, 
      dp_id_stage_regfile_DataPath_Physical_RF_n768, 
      dp_id_stage_regfile_DataPath_Physical_RF_n767, 
      dp_id_stage_regfile_DataPath_Physical_RF_n766, 
      dp_id_stage_regfile_DataPath_Physical_RF_n765, 
      dp_id_stage_regfile_DataPath_Physical_RF_n764, 
      dp_id_stage_regfile_DataPath_Physical_RF_n763, 
      dp_id_stage_regfile_DataPath_Physical_RF_n762, 
      dp_id_stage_regfile_DataPath_Physical_RF_n761, 
      dp_id_stage_regfile_DataPath_Physical_RF_n760, 
      dp_id_stage_regfile_DataPath_Physical_RF_n759, 
      dp_id_stage_regfile_DataPath_Physical_RF_n758, 
      dp_id_stage_regfile_DataPath_Physical_RF_n757, 
      dp_id_stage_regfile_DataPath_Physical_RF_n756, 
      dp_id_stage_regfile_DataPath_Physical_RF_n755, 
      dp_id_stage_regfile_DataPath_Physical_RF_n754, 
      dp_id_stage_regfile_DataPath_Physical_RF_n753, 
      dp_id_stage_regfile_DataPath_Physical_RF_n752, 
      dp_id_stage_regfile_DataPath_Physical_RF_n751, 
      dp_id_stage_regfile_DataPath_Physical_RF_n750, 
      dp_id_stage_regfile_DataPath_Physical_RF_n749, 
      dp_id_stage_regfile_DataPath_Physical_RF_n748, 
      dp_id_stage_regfile_DataPath_Physical_RF_n747, 
      dp_id_stage_regfile_DataPath_Physical_RF_n746, 
      dp_id_stage_regfile_DataPath_Physical_RF_n745, 
      dp_id_stage_regfile_DataPath_Physical_RF_n744, 
      dp_id_stage_regfile_DataPath_Physical_RF_n743, 
      dp_id_stage_regfile_DataPath_Physical_RF_n742, 
      dp_id_stage_regfile_DataPath_Physical_RF_n741, 
      dp_id_stage_regfile_DataPath_Physical_RF_n740, 
      dp_id_stage_regfile_DataPath_Physical_RF_n739, 
      dp_id_stage_regfile_DataPath_Physical_RF_n738, 
      dp_id_stage_regfile_DataPath_Physical_RF_n737, 
      dp_id_stage_regfile_DataPath_Physical_RF_n736, 
      dp_id_stage_regfile_DataPath_Physical_RF_n735, 
      dp_id_stage_regfile_DataPath_Physical_RF_n734, 
      dp_id_stage_regfile_DataPath_Physical_RF_n733, 
      dp_id_stage_regfile_DataPath_Physical_RF_n732, 
      dp_id_stage_regfile_DataPath_Physical_RF_n731, 
      dp_id_stage_regfile_DataPath_Physical_RF_n730, 
      dp_id_stage_regfile_DataPath_Physical_RF_n729, 
      dp_id_stage_regfile_DataPath_Physical_RF_n728, 
      dp_id_stage_regfile_DataPath_Physical_RF_n727, 
      dp_id_stage_regfile_DataPath_Physical_RF_n726, 
      dp_id_stage_regfile_DataPath_Physical_RF_n725, 
      dp_id_stage_regfile_DataPath_Physical_RF_n724, 
      dp_id_stage_regfile_DataPath_Physical_RF_n723, 
      dp_id_stage_regfile_DataPath_Physical_RF_n722, 
      dp_id_stage_regfile_DataPath_Physical_RF_n721, 
      dp_id_stage_regfile_DataPath_Physical_RF_n720, 
      dp_id_stage_regfile_DataPath_Physical_RF_n719, 
      dp_id_stage_regfile_DataPath_Physical_RF_n718, 
      dp_id_stage_regfile_DataPath_Physical_RF_n717, 
      dp_id_stage_regfile_DataPath_Physical_RF_n716, 
      dp_id_stage_regfile_DataPath_Physical_RF_n715, 
      dp_id_stage_regfile_DataPath_Physical_RF_n714, 
      dp_id_stage_regfile_DataPath_Physical_RF_n713, 
      dp_id_stage_regfile_DataPath_Physical_RF_n712, 
      dp_id_stage_regfile_DataPath_Physical_RF_n711, 
      dp_id_stage_regfile_DataPath_Physical_RF_n710, 
      dp_id_stage_regfile_DataPath_Physical_RF_n709, 
      dp_id_stage_regfile_DataPath_Physical_RF_n708, 
      dp_id_stage_regfile_DataPath_Physical_RF_n707, 
      dp_id_stage_regfile_DataPath_Physical_RF_n706, 
      dp_id_stage_regfile_DataPath_Physical_RF_n705, 
      dp_id_stage_regfile_DataPath_Physical_RF_n704, 
      dp_id_stage_regfile_DataPath_Physical_RF_n703, 
      dp_id_stage_regfile_DataPath_Physical_RF_n702, 
      dp_id_stage_regfile_DataPath_Physical_RF_n701, 
      dp_id_stage_regfile_DataPath_Physical_RF_n700, 
      dp_id_stage_regfile_DataPath_Physical_RF_n699, 
      dp_id_stage_regfile_DataPath_Physical_RF_n698, 
      dp_id_stage_regfile_DataPath_Physical_RF_n697, 
      dp_id_stage_regfile_DataPath_Physical_RF_n696, 
      dp_id_stage_regfile_DataPath_Physical_RF_n695, 
      dp_id_stage_regfile_DataPath_Physical_RF_n694, 
      dp_id_stage_regfile_DataPath_Physical_RF_n693, 
      dp_id_stage_regfile_DataPath_Physical_RF_n692, 
      dp_id_stage_regfile_DataPath_Physical_RF_n691, 
      dp_id_stage_regfile_DataPath_Physical_RF_n690, 
      dp_id_stage_regfile_DataPath_Physical_RF_n689, 
      dp_id_stage_regfile_DataPath_Physical_RF_n688, 
      dp_id_stage_regfile_DataPath_Physical_RF_n687, 
      dp_id_stage_regfile_DataPath_Physical_RF_n686, 
      dp_id_stage_regfile_DataPath_Physical_RF_n685, 
      dp_id_stage_regfile_DataPath_Physical_RF_n684, 
      dp_id_stage_regfile_DataPath_Physical_RF_n683, 
      dp_id_stage_regfile_DataPath_Physical_RF_n682, 
      dp_id_stage_regfile_DataPath_Physical_RF_n681, 
      dp_id_stage_regfile_DataPath_Physical_RF_n680, 
      dp_id_stage_regfile_DataPath_Physical_RF_n679, 
      dp_id_stage_regfile_DataPath_Physical_RF_n678, 
      dp_id_stage_regfile_DataPath_Physical_RF_n677, 
      dp_id_stage_regfile_DataPath_Physical_RF_n676, 
      dp_id_stage_regfile_DataPath_Physical_RF_n675, 
      dp_id_stage_regfile_DataPath_Physical_RF_n674, 
      dp_id_stage_regfile_DataPath_Physical_RF_n673, 
      dp_id_stage_regfile_DataPath_Physical_RF_n672, 
      dp_id_stage_regfile_DataPath_Physical_RF_n671, 
      dp_id_stage_regfile_DataPath_Physical_RF_n670, 
      dp_id_stage_regfile_DataPath_Physical_RF_n669, 
      dp_id_stage_regfile_DataPath_Physical_RF_n668, 
      dp_id_stage_regfile_DataPath_Physical_RF_n667, 
      dp_id_stage_regfile_DataPath_Physical_RF_n666, 
      dp_id_stage_regfile_DataPath_Physical_RF_n665, 
      dp_id_stage_regfile_DataPath_Physical_RF_n664, 
      dp_id_stage_regfile_DataPath_Physical_RF_n663, 
      dp_id_stage_regfile_DataPath_Physical_RF_n662, 
      dp_id_stage_regfile_DataPath_Physical_RF_n661, 
      dp_id_stage_regfile_DataPath_Physical_RF_n660, 
      dp_id_stage_regfile_DataPath_Physical_RF_n659, 
      dp_id_stage_regfile_DataPath_Physical_RF_n658, 
      dp_id_stage_regfile_DataPath_Physical_RF_n657, 
      dp_id_stage_regfile_DataPath_Physical_RF_n656, 
      dp_id_stage_regfile_DataPath_Physical_RF_n655, 
      dp_id_stage_regfile_DataPath_Physical_RF_n654, 
      dp_id_stage_regfile_DataPath_Physical_RF_n653, 
      dp_id_stage_regfile_DataPath_Physical_RF_n652, 
      dp_id_stage_regfile_DataPath_Physical_RF_n651, 
      dp_id_stage_regfile_DataPath_Physical_RF_n650, 
      dp_id_stage_regfile_DataPath_Physical_RF_n649, 
      dp_id_stage_regfile_DataPath_Physical_RF_n648, 
      dp_id_stage_regfile_DataPath_Physical_RF_n647, 
      dp_id_stage_regfile_DataPath_Physical_RF_n646, 
      dp_id_stage_regfile_DataPath_Physical_RF_n645, 
      dp_id_stage_regfile_DataPath_Physical_RF_n644, 
      dp_id_stage_regfile_DataPath_Physical_RF_n643, 
      dp_id_stage_regfile_DataPath_Physical_RF_n642, 
      dp_id_stage_regfile_DataPath_Physical_RF_n641, 
      dp_id_stage_regfile_DataPath_Physical_RF_n640, 
      dp_id_stage_regfile_DataPath_Physical_RF_n639, 
      dp_id_stage_regfile_DataPath_Physical_RF_n638, 
      dp_id_stage_regfile_DataPath_Physical_RF_n637, 
      dp_id_stage_regfile_DataPath_Physical_RF_n636, 
      dp_id_stage_regfile_DataPath_Physical_RF_n635, 
      dp_id_stage_regfile_DataPath_Physical_RF_n634, 
      dp_id_stage_regfile_DataPath_Physical_RF_n633, 
      dp_id_stage_regfile_DataPath_Physical_RF_n632, 
      dp_id_stage_regfile_DataPath_Physical_RF_n631, 
      dp_id_stage_regfile_DataPath_Physical_RF_n630, 
      dp_id_stage_regfile_DataPath_Physical_RF_n629, 
      dp_id_stage_regfile_DataPath_Physical_RF_n628, 
      dp_id_stage_regfile_DataPath_Physical_RF_n627, 
      dp_id_stage_regfile_DataPath_Physical_RF_n626, 
      dp_id_stage_regfile_DataPath_Physical_RF_n625, 
      dp_id_stage_regfile_DataPath_Physical_RF_n624, 
      dp_id_stage_regfile_DataPath_Physical_RF_n623, 
      dp_id_stage_regfile_DataPath_Physical_RF_n622, 
      dp_id_stage_regfile_DataPath_Physical_RF_n621, 
      dp_id_stage_regfile_DataPath_Physical_RF_n620, 
      dp_id_stage_regfile_DataPath_Physical_RF_n619, 
      dp_id_stage_regfile_DataPath_Physical_RF_n618, 
      dp_id_stage_regfile_DataPath_Physical_RF_n617, 
      dp_id_stage_regfile_DataPath_Physical_RF_n616, 
      dp_id_stage_regfile_DataPath_Physical_RF_n615, 
      dp_id_stage_regfile_DataPath_Physical_RF_n614, 
      dp_id_stage_regfile_DataPath_Physical_RF_n613, 
      dp_id_stage_regfile_DataPath_Physical_RF_n612, 
      dp_id_stage_regfile_DataPath_Physical_RF_n611, 
      dp_id_stage_regfile_DataPath_Physical_RF_n610, 
      dp_id_stage_regfile_DataPath_Physical_RF_n609, 
      dp_id_stage_regfile_DataPath_Physical_RF_n608, 
      dp_id_stage_regfile_DataPath_Physical_RF_n607, 
      dp_id_stage_regfile_DataPath_Physical_RF_n606, 
      dp_id_stage_regfile_DataPath_Physical_RF_n605, 
      dp_id_stage_regfile_DataPath_Physical_RF_n604, 
      dp_id_stage_regfile_DataPath_Physical_RF_n603, 
      dp_id_stage_regfile_DataPath_Physical_RF_n602, 
      dp_id_stage_regfile_DataPath_Physical_RF_n601, 
      dp_id_stage_regfile_DataPath_Physical_RF_n600, 
      dp_id_stage_regfile_DataPath_Physical_RF_n599, 
      dp_id_stage_regfile_DataPath_Physical_RF_n598, 
      dp_id_stage_regfile_DataPath_Physical_RF_n597, 
      dp_id_stage_regfile_DataPath_Physical_RF_n596, 
      dp_id_stage_regfile_DataPath_Physical_RF_n595, 
      dp_id_stage_regfile_DataPath_Physical_RF_n594, 
      dp_id_stage_regfile_DataPath_Physical_RF_n593, 
      dp_id_stage_regfile_DataPath_Physical_RF_n592, 
      dp_id_stage_regfile_DataPath_Physical_RF_n591, 
      dp_id_stage_regfile_DataPath_Physical_RF_n590, 
      dp_id_stage_regfile_DataPath_Physical_RF_n589, 
      dp_id_stage_regfile_DataPath_Physical_RF_n588, 
      dp_id_stage_regfile_DataPath_Physical_RF_n587, 
      dp_id_stage_regfile_DataPath_Physical_RF_n586, 
      dp_id_stage_regfile_DataPath_Physical_RF_n585, 
      dp_id_stage_regfile_DataPath_Physical_RF_n584, 
      dp_id_stage_regfile_DataPath_Physical_RF_n583, 
      dp_id_stage_regfile_DataPath_Physical_RF_n582, 
      dp_id_stage_regfile_DataPath_Physical_RF_n581, 
      dp_id_stage_regfile_DataPath_Physical_RF_n580, 
      dp_id_stage_regfile_DataPath_Physical_RF_n579, 
      dp_id_stage_regfile_DataPath_Physical_RF_n578, 
      dp_id_stage_regfile_DataPath_Physical_RF_n577, 
      dp_id_stage_regfile_DataPath_Physical_RF_n576, 
      dp_id_stage_regfile_DataPath_Physical_RF_n575, 
      dp_id_stage_regfile_DataPath_Physical_RF_n574, 
      dp_id_stage_regfile_DataPath_Physical_RF_n573, 
      dp_id_stage_regfile_DataPath_Physical_RF_n572, 
      dp_id_stage_regfile_DataPath_Physical_RF_n571, 
      dp_id_stage_regfile_DataPath_Physical_RF_n570, 
      dp_id_stage_regfile_DataPath_Physical_RF_n569, 
      dp_id_stage_regfile_DataPath_Physical_RF_n568, 
      dp_id_stage_regfile_DataPath_Physical_RF_n567, 
      dp_id_stage_regfile_DataPath_Physical_RF_n566, 
      dp_id_stage_regfile_DataPath_Physical_RF_n565, 
      dp_id_stage_regfile_DataPath_Physical_RF_n564, 
      dp_id_stage_regfile_DataPath_Physical_RF_n563, 
      dp_id_stage_regfile_DataPath_Physical_RF_n562, 
      dp_id_stage_regfile_DataPath_Physical_RF_n561, 
      dp_id_stage_regfile_DataPath_Physical_RF_n560, 
      dp_id_stage_regfile_DataPath_Physical_RF_n559, 
      dp_id_stage_regfile_DataPath_Physical_RF_n558, 
      dp_id_stage_regfile_DataPath_Physical_RF_n557, 
      dp_id_stage_regfile_DataPath_Physical_RF_n556, 
      dp_id_stage_regfile_DataPath_Physical_RF_n555, 
      dp_id_stage_regfile_DataPath_Physical_RF_n554, 
      dp_id_stage_regfile_DataPath_Physical_RF_n553, 
      dp_id_stage_regfile_DataPath_Physical_RF_n552, 
      dp_id_stage_regfile_DataPath_Physical_RF_n551, 
      dp_id_stage_regfile_DataPath_Physical_RF_n550, 
      dp_id_stage_regfile_DataPath_Physical_RF_n549, 
      dp_id_stage_regfile_DataPath_Physical_RF_n548, 
      dp_id_stage_regfile_DataPath_Physical_RF_n547, 
      dp_id_stage_regfile_DataPath_Physical_RF_n546, 
      dp_id_stage_regfile_DataPath_Physical_RF_n545, 
      dp_id_stage_regfile_DataPath_Physical_RF_n544, 
      dp_id_stage_regfile_DataPath_Physical_RF_n543, 
      dp_id_stage_regfile_DataPath_Physical_RF_n542, 
      dp_id_stage_regfile_DataPath_Physical_RF_n541, 
      dp_id_stage_regfile_DataPath_Physical_RF_n540, 
      dp_id_stage_regfile_DataPath_Physical_RF_n539, 
      dp_id_stage_regfile_DataPath_Physical_RF_n538, 
      dp_id_stage_regfile_DataPath_Physical_RF_n537, 
      dp_id_stage_regfile_DataPath_Physical_RF_n536, 
      dp_id_stage_regfile_DataPath_Physical_RF_n535, 
      dp_id_stage_regfile_DataPath_Physical_RF_n534, 
      dp_id_stage_regfile_DataPath_Physical_RF_n533, 
      dp_id_stage_regfile_DataPath_Physical_RF_n532, 
      dp_id_stage_regfile_DataPath_Physical_RF_n531, 
      dp_id_stage_regfile_DataPath_Physical_RF_n530, 
      dp_id_stage_regfile_DataPath_Physical_RF_n529, 
      dp_id_stage_regfile_DataPath_Physical_RF_n528, 
      dp_id_stage_regfile_DataPath_Physical_RF_n527, 
      dp_id_stage_regfile_DataPath_Physical_RF_n526, 
      dp_id_stage_regfile_DataPath_Physical_RF_n525, 
      dp_id_stage_regfile_DataPath_Physical_RF_n524, 
      dp_id_stage_regfile_DataPath_Physical_RF_n523, 
      dp_id_stage_regfile_DataPath_Physical_RF_n522, 
      dp_id_stage_regfile_DataPath_Physical_RF_n521, 
      dp_id_stage_regfile_DataPath_Physical_RF_n520, 
      dp_id_stage_regfile_DataPath_Physical_RF_n519, 
      dp_id_stage_regfile_DataPath_Physical_RF_n518, 
      dp_id_stage_regfile_DataPath_Physical_RF_n517, 
      dp_id_stage_regfile_DataPath_Physical_RF_n516, 
      dp_id_stage_regfile_DataPath_Physical_RF_n515, 
      dp_id_stage_regfile_DataPath_Physical_RF_n514, 
      dp_id_stage_regfile_DataPath_Physical_RF_n513, 
      dp_id_stage_regfile_DataPath_Physical_RF_n512, 
      dp_id_stage_regfile_DataPath_Physical_RF_n511, 
      dp_id_stage_regfile_DataPath_Physical_RF_n510, 
      dp_id_stage_regfile_DataPath_Physical_RF_n509, 
      dp_id_stage_regfile_DataPath_Physical_RF_n508, 
      dp_id_stage_regfile_DataPath_Physical_RF_n507, 
      dp_id_stage_regfile_DataPath_Physical_RF_n506, 
      dp_id_stage_regfile_DataPath_Physical_RF_n505, 
      dp_id_stage_regfile_DataPath_Physical_RF_n504, 
      dp_id_stage_regfile_DataPath_Physical_RF_n503, 
      dp_id_stage_regfile_DataPath_Physical_RF_n502, 
      dp_id_stage_regfile_DataPath_Physical_RF_n501, 
      dp_id_stage_regfile_DataPath_Physical_RF_n500, 
      dp_id_stage_regfile_DataPath_Physical_RF_n499, 
      dp_id_stage_regfile_DataPath_Physical_RF_n498, 
      dp_id_stage_regfile_DataPath_Physical_RF_n497, 
      dp_id_stage_regfile_DataPath_Physical_RF_n496, 
      dp_id_stage_regfile_DataPath_Physical_RF_n495, 
      dp_id_stage_regfile_DataPath_Physical_RF_n494, 
      dp_id_stage_regfile_DataPath_Physical_RF_n493, 
      dp_id_stage_regfile_DataPath_Physical_RF_n492, 
      dp_id_stage_regfile_DataPath_Physical_RF_n491, 
      dp_id_stage_regfile_DataPath_Physical_RF_n490, 
      dp_id_stage_regfile_DataPath_Physical_RF_n489, 
      dp_id_stage_regfile_DataPath_Physical_RF_n488, 
      dp_id_stage_regfile_DataPath_Physical_RF_n487, 
      dp_id_stage_regfile_DataPath_Physical_RF_n486, 
      dp_id_stage_regfile_DataPath_Physical_RF_n485, 
      dp_id_stage_regfile_DataPath_Physical_RF_n484, 
      dp_id_stage_regfile_DataPath_Physical_RF_n483, 
      dp_id_stage_regfile_DataPath_Physical_RF_n482, 
      dp_id_stage_regfile_DataPath_Physical_RF_n481, 
      dp_id_stage_regfile_DataPath_Physical_RF_n480, 
      dp_id_stage_regfile_DataPath_Physical_RF_n479, 
      dp_id_stage_regfile_DataPath_Physical_RF_n478, 
      dp_id_stage_regfile_DataPath_Physical_RF_n477, 
      dp_id_stage_regfile_DataPath_Physical_RF_n476, 
      dp_id_stage_regfile_DataPath_Physical_RF_n475, 
      dp_id_stage_regfile_DataPath_Physical_RF_n474, 
      dp_id_stage_regfile_DataPath_Physical_RF_n473, 
      dp_id_stage_regfile_DataPath_Physical_RF_n472, 
      dp_id_stage_regfile_DataPath_Physical_RF_n471, 
      dp_id_stage_regfile_DataPath_Physical_RF_n470, 
      dp_id_stage_regfile_DataPath_Physical_RF_n469, 
      dp_id_stage_regfile_DataPath_Physical_RF_n468, 
      dp_id_stage_regfile_DataPath_Physical_RF_n467, 
      dp_id_stage_regfile_DataPath_Physical_RF_n466, 
      dp_id_stage_regfile_DataPath_Physical_RF_n465, 
      dp_id_stage_regfile_DataPath_Physical_RF_n464, 
      dp_id_stage_regfile_DataPath_Physical_RF_n463, 
      dp_id_stage_regfile_DataPath_Physical_RF_n462, 
      dp_id_stage_regfile_DataPath_Physical_RF_n461, 
      dp_id_stage_regfile_DataPath_Physical_RF_n460, 
      dp_id_stage_regfile_DataPath_Physical_RF_n459, 
      dp_id_stage_regfile_DataPath_Physical_RF_n458, 
      dp_id_stage_regfile_DataPath_Physical_RF_n457, 
      dp_id_stage_regfile_DataPath_Physical_RF_n456, 
      dp_id_stage_regfile_DataPath_Physical_RF_n455, 
      dp_id_stage_regfile_DataPath_Physical_RF_n454, 
      dp_id_stage_regfile_DataPath_Physical_RF_n453, 
      dp_id_stage_regfile_DataPath_Physical_RF_n452, 
      dp_id_stage_regfile_DataPath_Physical_RF_n451, 
      dp_id_stage_regfile_DataPath_Physical_RF_n450, 
      dp_id_stage_regfile_DataPath_Physical_RF_n449, 
      dp_id_stage_regfile_DataPath_Physical_RF_n448, 
      dp_id_stage_regfile_DataPath_Physical_RF_n447, 
      dp_id_stage_regfile_DataPath_Physical_RF_n446, 
      dp_id_stage_regfile_DataPath_Physical_RF_n445, 
      dp_id_stage_regfile_DataPath_Physical_RF_n444, 
      dp_id_stage_regfile_DataPath_Physical_RF_n443, 
      dp_id_stage_regfile_DataPath_Physical_RF_n442, 
      dp_id_stage_regfile_DataPath_Physical_RF_n441, 
      dp_id_stage_regfile_DataPath_Physical_RF_n440, 
      dp_id_stage_regfile_DataPath_Physical_RF_n439, 
      dp_id_stage_regfile_DataPath_Physical_RF_n438, 
      dp_id_stage_regfile_DataPath_Physical_RF_n437, 
      dp_id_stage_regfile_DataPath_Physical_RF_n436, 
      dp_id_stage_regfile_DataPath_Physical_RF_n435, 
      dp_id_stage_regfile_DataPath_Physical_RF_n434, 
      dp_id_stage_regfile_DataPath_Physical_RF_n433, 
      dp_id_stage_regfile_DataPath_Physical_RF_n432, 
      dp_id_stage_regfile_DataPath_Physical_RF_n431, 
      dp_id_stage_regfile_DataPath_Physical_RF_n430, 
      dp_id_stage_regfile_DataPath_Physical_RF_n429, 
      dp_id_stage_regfile_DataPath_Physical_RF_n428, 
      dp_id_stage_regfile_DataPath_Physical_RF_n427, 
      dp_id_stage_regfile_DataPath_Physical_RF_n426, 
      dp_id_stage_regfile_DataPath_Physical_RF_n425, 
      dp_id_stage_regfile_DataPath_Physical_RF_n424, 
      dp_id_stage_regfile_DataPath_Physical_RF_n423, 
      dp_id_stage_regfile_DataPath_Physical_RF_n422, 
      dp_id_stage_regfile_DataPath_Physical_RF_n421, 
      dp_id_stage_regfile_DataPath_Physical_RF_n420, 
      dp_id_stage_regfile_DataPath_Physical_RF_n419, 
      dp_id_stage_regfile_DataPath_Physical_RF_n418, 
      dp_id_stage_regfile_DataPath_Physical_RF_n417, 
      dp_id_stage_regfile_DataPath_Physical_RF_n416, 
      dp_id_stage_regfile_DataPath_Physical_RF_n415, 
      dp_id_stage_regfile_DataPath_Physical_RF_n414, 
      dp_id_stage_regfile_DataPath_Physical_RF_n413, 
      dp_id_stage_regfile_DataPath_Physical_RF_n412, 
      dp_id_stage_regfile_DataPath_Physical_RF_n411, 
      dp_id_stage_regfile_DataPath_Physical_RF_n410, 
      dp_id_stage_regfile_DataPath_Physical_RF_n409, 
      dp_id_stage_regfile_DataPath_Physical_RF_n408, 
      dp_id_stage_regfile_DataPath_Physical_RF_n407, 
      dp_id_stage_regfile_DataPath_Physical_RF_n406, 
      dp_id_stage_regfile_DataPath_Physical_RF_n405, 
      dp_id_stage_regfile_DataPath_Physical_RF_n404, 
      dp_id_stage_regfile_DataPath_Physical_RF_n403, 
      dp_id_stage_regfile_DataPath_Physical_RF_n402, 
      dp_id_stage_regfile_DataPath_Physical_RF_n401, 
      dp_id_stage_regfile_DataPath_Physical_RF_n400, 
      dp_id_stage_regfile_DataPath_Physical_RF_n399, 
      dp_id_stage_regfile_DataPath_Physical_RF_n398, 
      dp_id_stage_regfile_DataPath_Physical_RF_n397, 
      dp_id_stage_regfile_DataPath_Physical_RF_n396, 
      dp_id_stage_regfile_DataPath_Physical_RF_n395, 
      dp_id_stage_regfile_DataPath_Physical_RF_n394, 
      dp_id_stage_regfile_DataPath_Physical_RF_n393, 
      dp_id_stage_regfile_DataPath_Physical_RF_n392, 
      dp_id_stage_regfile_DataPath_Physical_RF_n391, 
      dp_id_stage_regfile_DataPath_Physical_RF_n390, 
      dp_id_stage_regfile_DataPath_Physical_RF_n389, 
      dp_id_stage_regfile_DataPath_Physical_RF_n388, 
      dp_id_stage_regfile_DataPath_Physical_RF_n387, 
      dp_id_stage_regfile_DataPath_Physical_RF_n386, 
      dp_id_stage_regfile_DataPath_Physical_RF_n385, 
      dp_id_stage_regfile_DataPath_Physical_RF_n384, 
      dp_id_stage_regfile_DataPath_Physical_RF_n383, 
      dp_id_stage_regfile_DataPath_Physical_RF_n382, 
      dp_id_stage_regfile_DataPath_Physical_RF_n381, 
      dp_id_stage_regfile_DataPath_Physical_RF_n380, 
      dp_id_stage_regfile_DataPath_Physical_RF_n379, 
      dp_id_stage_regfile_DataPath_Physical_RF_n378, 
      dp_id_stage_regfile_DataPath_Physical_RF_n377, 
      dp_id_stage_regfile_DataPath_Physical_RF_n376, 
      dp_id_stage_regfile_DataPath_Physical_RF_n375, 
      dp_id_stage_regfile_DataPath_Physical_RF_n374, 
      dp_id_stage_regfile_DataPath_Physical_RF_n373, 
      dp_id_stage_regfile_DataPath_Physical_RF_n372, 
      dp_id_stage_regfile_DataPath_Physical_RF_n371, 
      dp_id_stage_regfile_DataPath_Physical_RF_n370, 
      dp_id_stage_regfile_DataPath_Physical_RF_n369, 
      dp_id_stage_regfile_DataPath_Physical_RF_n368, 
      dp_id_stage_regfile_DataPath_Physical_RF_n367, 
      dp_id_stage_regfile_DataPath_Physical_RF_n366, 
      dp_id_stage_regfile_DataPath_Physical_RF_n365, 
      dp_id_stage_regfile_DataPath_Physical_RF_n364, 
      dp_id_stage_regfile_DataPath_Physical_RF_n363, 
      dp_id_stage_regfile_DataPath_Physical_RF_n362, 
      dp_id_stage_regfile_DataPath_Physical_RF_n361, 
      dp_id_stage_regfile_DataPath_Physical_RF_n360, 
      dp_id_stage_regfile_DataPath_Physical_RF_n359, 
      dp_id_stage_regfile_DataPath_Physical_RF_n358, 
      dp_id_stage_regfile_DataPath_Physical_RF_n357, 
      dp_id_stage_regfile_DataPath_Physical_RF_n356, 
      dp_id_stage_regfile_DataPath_Physical_RF_n355, 
      dp_id_stage_regfile_DataPath_Physical_RF_n354, 
      dp_id_stage_regfile_DataPath_Physical_RF_n353, 
      dp_id_stage_regfile_DataPath_Physical_RF_n352, 
      dp_id_stage_regfile_DataPath_Physical_RF_n351, 
      dp_id_stage_regfile_DataPath_Physical_RF_n350, 
      dp_id_stage_regfile_DataPath_Physical_RF_n349, 
      dp_id_stage_regfile_DataPath_Physical_RF_n348, 
      dp_id_stage_regfile_DataPath_Physical_RF_n347, 
      dp_id_stage_regfile_DataPath_Physical_RF_n346, 
      dp_id_stage_regfile_DataPath_Physical_RF_n345, 
      dp_id_stage_regfile_DataPath_Physical_RF_n344, 
      dp_id_stage_regfile_DataPath_Physical_RF_n343, 
      dp_id_stage_regfile_DataPath_Physical_RF_n342, 
      dp_id_stage_regfile_DataPath_Physical_RF_n341, 
      dp_id_stage_regfile_DataPath_Physical_RF_n340, 
      dp_id_stage_regfile_DataPath_Physical_RF_n339, 
      dp_id_stage_regfile_DataPath_Physical_RF_n338, 
      dp_id_stage_regfile_DataPath_Physical_RF_n337, 
      dp_id_stage_regfile_DataPath_Physical_RF_n336, 
      dp_id_stage_regfile_DataPath_Physical_RF_n335, 
      dp_id_stage_regfile_DataPath_Physical_RF_n334, 
      dp_id_stage_regfile_DataPath_Physical_RF_n333, 
      dp_id_stage_regfile_DataPath_Physical_RF_n332, 
      dp_id_stage_regfile_DataPath_Physical_RF_n331, 
      dp_id_stage_regfile_DataPath_Physical_RF_n330, 
      dp_id_stage_regfile_DataPath_Physical_RF_n329, 
      dp_id_stage_regfile_DataPath_Physical_RF_n328, 
      dp_id_stage_regfile_DataPath_Physical_RF_n327, 
      dp_id_stage_regfile_DataPath_Physical_RF_n326, 
      dp_id_stage_regfile_DataPath_Physical_RF_n325, 
      dp_id_stage_regfile_DataPath_Physical_RF_n324, 
      dp_id_stage_regfile_DataPath_Physical_RF_n323, 
      dp_id_stage_regfile_DataPath_Physical_RF_n322, 
      dp_id_stage_regfile_DataPath_Physical_RF_n321, 
      dp_id_stage_regfile_DataPath_Physical_RF_n320, 
      dp_id_stage_regfile_DataPath_Physical_RF_n319, 
      dp_id_stage_regfile_DataPath_Physical_RF_n318, 
      dp_id_stage_regfile_DataPath_Physical_RF_n317, 
      dp_id_stage_regfile_DataPath_Physical_RF_n316, 
      dp_id_stage_regfile_DataPath_Physical_RF_n315, 
      dp_id_stage_regfile_DataPath_Physical_RF_n314, 
      dp_id_stage_regfile_DataPath_Physical_RF_n313, 
      dp_id_stage_regfile_DataPath_Physical_RF_n312, 
      dp_id_stage_regfile_DataPath_Physical_RF_n311, 
      dp_id_stage_regfile_DataPath_Physical_RF_n310, 
      dp_id_stage_regfile_DataPath_Physical_RF_n309, 
      dp_id_stage_regfile_DataPath_Physical_RF_n308, 
      dp_id_stage_regfile_DataPath_Physical_RF_n307, 
      dp_id_stage_regfile_DataPath_Physical_RF_n306, 
      dp_id_stage_regfile_DataPath_Physical_RF_n305, 
      dp_id_stage_regfile_DataPath_Physical_RF_n304, 
      dp_id_stage_regfile_DataPath_Physical_RF_n303, 
      dp_id_stage_regfile_DataPath_Physical_RF_n302, 
      dp_id_stage_regfile_DataPath_Physical_RF_n301, 
      dp_id_stage_regfile_DataPath_Physical_RF_n300, 
      dp_id_stage_regfile_DataPath_Physical_RF_n299, 
      dp_id_stage_regfile_DataPath_Physical_RF_n298, 
      dp_id_stage_regfile_DataPath_Physical_RF_n297, 
      dp_id_stage_regfile_DataPath_Physical_RF_n296, 
      dp_id_stage_regfile_DataPath_Physical_RF_n295, 
      dp_id_stage_regfile_DataPath_Physical_RF_n294, 
      dp_id_stage_regfile_DataPath_Physical_RF_n293, 
      dp_id_stage_regfile_DataPath_Physical_RF_n292, 
      dp_id_stage_regfile_DataPath_Physical_RF_n291, 
      dp_id_stage_regfile_DataPath_Physical_RF_n290, 
      dp_id_stage_regfile_DataPath_Physical_RF_n289, 
      dp_id_stage_regfile_DataPath_Physical_RF_n288, 
      dp_id_stage_regfile_DataPath_Physical_RF_n287, 
      dp_id_stage_regfile_DataPath_Physical_RF_n286, 
      dp_id_stage_regfile_DataPath_Physical_RF_n285, 
      dp_id_stage_regfile_DataPath_Physical_RF_n284, 
      dp_id_stage_regfile_DataPath_Physical_RF_n283, 
      dp_id_stage_regfile_DataPath_Physical_RF_n282, 
      dp_id_stage_regfile_DataPath_Physical_RF_n281, 
      dp_id_stage_regfile_DataPath_Physical_RF_n280, 
      dp_id_stage_regfile_DataPath_Physical_RF_n279, 
      dp_id_stage_regfile_DataPath_Physical_RF_n278, 
      dp_id_stage_regfile_DataPath_Physical_RF_n277, 
      dp_id_stage_regfile_DataPath_Physical_RF_n276, 
      dp_id_stage_regfile_DataPath_Physical_RF_n275, 
      dp_id_stage_regfile_DataPath_Physical_RF_n274, 
      dp_id_stage_regfile_DataPath_Physical_RF_n273, 
      dp_id_stage_regfile_DataPath_Physical_RF_n272, 
      dp_id_stage_regfile_DataPath_Physical_RF_n271, 
      dp_id_stage_regfile_DataPath_Physical_RF_n270, 
      dp_id_stage_regfile_DataPath_Physical_RF_n269, 
      dp_id_stage_regfile_DataPath_Physical_RF_n268, 
      dp_id_stage_regfile_DataPath_Physical_RF_n267, 
      dp_id_stage_regfile_DataPath_Physical_RF_n266, 
      dp_id_stage_regfile_DataPath_Physical_RF_n265, 
      dp_id_stage_regfile_DataPath_Physical_RF_n264, 
      dp_id_stage_regfile_DataPath_Physical_RF_n263, 
      dp_id_stage_regfile_DataPath_Physical_RF_n262, 
      dp_id_stage_regfile_DataPath_Physical_RF_n261, 
      dp_id_stage_regfile_DataPath_Physical_RF_n260, 
      dp_id_stage_regfile_DataPath_Physical_RF_n259, 
      dp_id_stage_regfile_DataPath_Physical_RF_n258, 
      dp_id_stage_regfile_DataPath_Physical_RF_n257, 
      dp_id_stage_regfile_DataPath_Physical_RF_n256, 
      dp_id_stage_regfile_DataPath_Physical_RF_n255, 
      dp_id_stage_regfile_DataPath_Physical_RF_n254, 
      dp_id_stage_regfile_DataPath_Physical_RF_n253, 
      dp_id_stage_regfile_DataPath_Physical_RF_n252, 
      dp_id_stage_regfile_DataPath_Physical_RF_n251, 
      dp_id_stage_regfile_DataPath_Physical_RF_n250, 
      dp_id_stage_regfile_DataPath_Physical_RF_n249, 
      dp_id_stage_regfile_DataPath_Physical_RF_n248, 
      dp_id_stage_regfile_DataPath_Physical_RF_n247, 
      dp_id_stage_regfile_DataPath_Physical_RF_n246, 
      dp_id_stage_regfile_DataPath_Physical_RF_n245, 
      dp_id_stage_regfile_DataPath_Physical_RF_n244, 
      dp_id_stage_regfile_DataPath_Physical_RF_n243, 
      dp_id_stage_regfile_DataPath_Physical_RF_n242, 
      dp_id_stage_regfile_DataPath_Physical_RF_n241, 
      dp_id_stage_regfile_DataPath_Physical_RF_n240, 
      dp_id_stage_regfile_DataPath_Physical_RF_n239, 
      dp_id_stage_regfile_DataPath_Physical_RF_n238, 
      dp_id_stage_regfile_DataPath_Physical_RF_n237, 
      dp_id_stage_regfile_DataPath_Physical_RF_n236, 
      dp_id_stage_regfile_DataPath_Physical_RF_n235, 
      dp_id_stage_regfile_DataPath_Physical_RF_n234, 
      dp_id_stage_regfile_DataPath_Physical_RF_n233, 
      dp_id_stage_regfile_DataPath_Physical_RF_n232, 
      dp_id_stage_regfile_DataPath_Physical_RF_n231, 
      dp_id_stage_regfile_DataPath_Physical_RF_n230, 
      dp_id_stage_regfile_DataPath_Physical_RF_n229, 
      dp_id_stage_regfile_DataPath_Physical_RF_n228, 
      dp_id_stage_regfile_DataPath_Physical_RF_n227, 
      dp_id_stage_regfile_DataPath_Physical_RF_n226, 
      dp_id_stage_regfile_DataPath_Physical_RF_n225, 
      dp_id_stage_regfile_DataPath_Physical_RF_n224, 
      dp_id_stage_regfile_DataPath_Physical_RF_n223, 
      dp_id_stage_regfile_DataPath_Physical_RF_n222, 
      dp_id_stage_regfile_DataPath_Physical_RF_n221, 
      dp_id_stage_regfile_DataPath_Physical_RF_n220, 
      dp_id_stage_regfile_DataPath_Physical_RF_n219, 
      dp_id_stage_regfile_DataPath_Physical_RF_n218, 
      dp_id_stage_regfile_DataPath_Physical_RF_n217, 
      dp_id_stage_regfile_DataPath_Physical_RF_n216, 
      dp_id_stage_regfile_DataPath_Physical_RF_n215, 
      dp_id_stage_regfile_DataPath_Physical_RF_n214, 
      dp_id_stage_regfile_DataPath_Physical_RF_n213, 
      dp_id_stage_regfile_DataPath_Physical_RF_n212, 
      dp_id_stage_regfile_DataPath_Physical_RF_n211, 
      dp_id_stage_regfile_DataPath_Physical_RF_n210, 
      dp_id_stage_regfile_DataPath_Physical_RF_n209, 
      dp_id_stage_regfile_DataPath_Physical_RF_n208, 
      dp_id_stage_regfile_DataPath_Physical_RF_n207, 
      dp_id_stage_regfile_DataPath_Physical_RF_n206, 
      dp_id_stage_regfile_DataPath_Physical_RF_n205, 
      dp_id_stage_regfile_DataPath_Physical_RF_n204, 
      dp_id_stage_regfile_DataPath_Physical_RF_n203, 
      dp_id_stage_regfile_DataPath_Physical_RF_n202, 
      dp_id_stage_regfile_DataPath_Physical_RF_n201, 
      dp_id_stage_regfile_DataPath_Physical_RF_n200, 
      dp_id_stage_regfile_DataPath_Physical_RF_n199, 
      dp_id_stage_regfile_DataPath_Physical_RF_n198, 
      dp_id_stage_regfile_DataPath_Physical_RF_n197, 
      dp_id_stage_regfile_DataPath_Physical_RF_n196, 
      dp_id_stage_regfile_DataPath_Physical_RF_n195, 
      dp_id_stage_regfile_DataPath_Physical_RF_n194, 
      dp_id_stage_regfile_DataPath_Physical_RF_n193, 
      dp_id_stage_regfile_DataPath_Physical_RF_n192, 
      dp_id_stage_regfile_DataPath_Physical_RF_n191, 
      dp_id_stage_regfile_DataPath_Physical_RF_n190, 
      dp_id_stage_regfile_DataPath_Physical_RF_n189, 
      dp_id_stage_regfile_DataPath_Physical_RF_n188, 
      dp_id_stage_regfile_DataPath_Physical_RF_n187, 
      dp_id_stage_regfile_DataPath_Physical_RF_n186, 
      dp_id_stage_regfile_DataPath_Physical_RF_n185, 
      dp_id_stage_regfile_DataPath_Physical_RF_n184, 
      dp_id_stage_regfile_DataPath_Physical_RF_n183, 
      dp_id_stage_regfile_DataPath_Physical_RF_n182, 
      dp_id_stage_regfile_DataPath_Physical_RF_n181, 
      dp_id_stage_regfile_DataPath_Physical_RF_n180, 
      dp_id_stage_regfile_DataPath_Physical_RF_n179, 
      dp_id_stage_regfile_DataPath_Physical_RF_n178, 
      dp_id_stage_regfile_DataPath_Physical_RF_n177, 
      dp_id_stage_regfile_DataPath_Physical_RF_n176, 
      dp_id_stage_regfile_DataPath_Physical_RF_n175, 
      dp_id_stage_regfile_DataPath_Physical_RF_n174, 
      dp_id_stage_regfile_DataPath_Physical_RF_n173, 
      dp_id_stage_regfile_DataPath_Physical_RF_n172, 
      dp_id_stage_regfile_DataPath_Physical_RF_n171, 
      dp_id_stage_regfile_DataPath_Physical_RF_n170, 
      dp_id_stage_regfile_DataPath_Physical_RF_n169, 
      dp_id_stage_regfile_DataPath_Physical_RF_n168, 
      dp_id_stage_regfile_DataPath_Physical_RF_n167, 
      dp_id_stage_regfile_DataPath_Physical_RF_n166, 
      dp_id_stage_regfile_DataPath_Physical_RF_n165, 
      dp_id_stage_regfile_DataPath_Physical_RF_n164, 
      dp_id_stage_regfile_DataPath_Physical_RF_n163, 
      dp_id_stage_regfile_DataPath_Physical_RF_n162, 
      dp_id_stage_regfile_DataPath_Physical_RF_n161, 
      dp_id_stage_regfile_DataPath_Physical_RF_n160, 
      dp_id_stage_regfile_DataPath_Physical_RF_n159, 
      dp_id_stage_regfile_DataPath_Physical_RF_n158, 
      dp_id_stage_regfile_DataPath_Physical_RF_n157, 
      dp_id_stage_regfile_DataPath_Physical_RF_n156, 
      dp_id_stage_regfile_DataPath_Physical_RF_n155, 
      dp_id_stage_regfile_DataPath_Physical_RF_n154, 
      dp_id_stage_regfile_DataPath_Physical_RF_n153, 
      dp_id_stage_regfile_DataPath_Physical_RF_n152, 
      dp_id_stage_regfile_DataPath_Physical_RF_n151, 
      dp_id_stage_regfile_DataPath_Physical_RF_n150, 
      dp_id_stage_regfile_DataPath_Physical_RF_n149, 
      dp_id_stage_regfile_DataPath_Physical_RF_n148, 
      dp_id_stage_regfile_DataPath_Physical_RF_n147, 
      dp_id_stage_regfile_DataPath_Physical_RF_n146, 
      dp_id_stage_regfile_DataPath_Physical_RF_n145, 
      dp_id_stage_regfile_DataPath_Physical_RF_n144, 
      dp_id_stage_regfile_DataPath_Physical_RF_n143, 
      dp_id_stage_regfile_DataPath_Physical_RF_n142, 
      dp_id_stage_regfile_DataPath_Physical_RF_n141, 
      dp_id_stage_regfile_DataPath_Physical_RF_n140, 
      dp_id_stage_regfile_DataPath_Physical_RF_n139, 
      dp_id_stage_regfile_DataPath_Physical_RF_n138, 
      dp_id_stage_regfile_DataPath_Physical_RF_n137, 
      dp_id_stage_regfile_DataPath_Physical_RF_n136, 
      dp_id_stage_regfile_DataPath_Physical_RF_n135, 
      dp_id_stage_regfile_DataPath_Physical_RF_n134, 
      dp_id_stage_regfile_DataPath_Physical_RF_n133, 
      dp_id_stage_regfile_DataPath_Physical_RF_n132, 
      dp_id_stage_regfile_DataPath_Physical_RF_n131, 
      dp_id_stage_regfile_DataPath_Physical_RF_n130, 
      dp_id_stage_regfile_DataPath_Physical_RF_n129, 
      dp_id_stage_regfile_DataPath_Physical_RF_n128, 
      dp_id_stage_regfile_DataPath_Physical_RF_n127, 
      dp_id_stage_regfile_DataPath_Physical_RF_n126, 
      dp_id_stage_regfile_DataPath_Physical_RF_n125, 
      dp_id_stage_regfile_DataPath_Physical_RF_n124, 
      dp_id_stage_regfile_DataPath_Physical_RF_n123, 
      dp_id_stage_regfile_DataPath_Physical_RF_n122, 
      dp_id_stage_regfile_DataPath_Physical_RF_n121, 
      dp_id_stage_regfile_DataPath_Physical_RF_n120, 
      dp_id_stage_regfile_DataPath_Physical_RF_n119, 
      dp_id_stage_regfile_DataPath_Physical_RF_n118, 
      dp_id_stage_regfile_DataPath_Physical_RF_n117, 
      dp_id_stage_regfile_DataPath_Physical_RF_n116, 
      dp_id_stage_regfile_DataPath_Physical_RF_n115, 
      dp_id_stage_regfile_DataPath_Physical_RF_n114, 
      dp_id_stage_regfile_DataPath_Physical_RF_n113, 
      dp_id_stage_regfile_DataPath_Physical_RF_n112, 
      dp_id_stage_regfile_DataPath_Physical_RF_n111, 
      dp_id_stage_regfile_DataPath_Physical_RF_n110, 
      dp_id_stage_regfile_DataPath_Physical_RF_n109, 
      dp_id_stage_regfile_DataPath_Physical_RF_n108, 
      dp_id_stage_regfile_DataPath_Physical_RF_n107, 
      dp_id_stage_regfile_DataPath_Physical_RF_n106, 
      dp_id_stage_regfile_DataPath_Physical_RF_n105, 
      dp_id_stage_regfile_DataPath_Physical_RF_n104, 
      dp_id_stage_regfile_DataPath_Physical_RF_n103, 
      dp_id_stage_regfile_DataPath_Physical_RF_n102, 
      dp_id_stage_regfile_DataPath_Physical_RF_n101, 
      dp_id_stage_regfile_DataPath_Physical_RF_n100, 
      dp_id_stage_regfile_DataPath_Physical_RF_n99, 
      dp_id_stage_regfile_DataPath_Physical_RF_n98, 
      dp_id_stage_regfile_DataPath_Physical_RF_n97, 
      dp_id_stage_regfile_DataPath_Physical_RF_n96, 
      dp_id_stage_regfile_DataPath_Physical_RF_n95, 
      dp_id_stage_regfile_DataPath_Physical_RF_n94, 
      dp_id_stage_regfile_DataPath_Physical_RF_n93, 
      dp_id_stage_regfile_DataPath_Physical_RF_n92, 
      dp_id_stage_regfile_DataPath_Physical_RF_n91, 
      dp_id_stage_regfile_DataPath_Physical_RF_n90, 
      dp_id_stage_regfile_DataPath_Physical_RF_n89, 
      dp_id_stage_regfile_DataPath_Physical_RF_n88, 
      dp_id_stage_regfile_DataPath_Physical_RF_n87, 
      dp_id_stage_regfile_DataPath_Physical_RF_n86, 
      dp_id_stage_regfile_DataPath_Physical_RF_n85, 
      dp_id_stage_regfile_DataPath_Physical_RF_n84, 
      dp_id_stage_regfile_DataPath_Physical_RF_n83, 
      dp_id_stage_regfile_DataPath_Physical_RF_n82, 
      dp_id_stage_regfile_DataPath_Physical_RF_n81, 
      dp_id_stage_regfile_DataPath_Physical_RF_n80, 
      dp_id_stage_regfile_DataPath_Physical_RF_n79, 
      dp_id_stage_regfile_DataPath_Physical_RF_n78, 
      dp_id_stage_regfile_DataPath_Physical_RF_n77, 
      dp_id_stage_regfile_DataPath_Physical_RF_n76, 
      dp_id_stage_regfile_DataPath_Physical_RF_n75, 
      dp_id_stage_regfile_DataPath_Physical_RF_n74, 
      dp_id_stage_regfile_DataPath_Physical_RF_n73, 
      dp_id_stage_regfile_DataPath_Physical_RF_n72, 
      dp_id_stage_regfile_DataPath_Physical_RF_n71, 
      dp_id_stage_regfile_DataPath_Physical_RF_n70, 
      dp_id_stage_regfile_DataPath_Physical_RF_n69, 
      dp_id_stage_regfile_DataPath_Physical_RF_n68, 
      dp_id_stage_regfile_DataPath_Physical_RF_n67, 
      dp_id_stage_regfile_DataPath_Physical_RF_n66, 
      dp_id_stage_regfile_DataPath_Physical_RF_n65, 
      dp_id_stage_regfile_DataPath_Physical_RF_n64, 
      dp_id_stage_regfile_DataPath_Physical_RF_n63, 
      dp_id_stage_regfile_DataPath_Physical_RF_n62, 
      dp_id_stage_regfile_DataPath_Physical_RF_n61, 
      dp_id_stage_regfile_DataPath_Physical_RF_n60, 
      dp_id_stage_regfile_DataPath_Physical_RF_n59, 
      dp_id_stage_regfile_DataPath_Physical_RF_n58, 
      dp_id_stage_regfile_DataPath_Physical_RF_n57, 
      dp_id_stage_regfile_DataPath_Physical_RF_n56, 
      dp_id_stage_regfile_DataPath_Physical_RF_n55, 
      dp_id_stage_regfile_DataPath_Physical_RF_n54, 
      dp_id_stage_regfile_DataPath_Physical_RF_n53, 
      dp_id_stage_regfile_DataPath_Physical_RF_n52, 
      dp_id_stage_regfile_DataPath_Physical_RF_n51, 
      dp_id_stage_regfile_DataPath_Physical_RF_n50, 
      dp_id_stage_regfile_DataPath_Physical_RF_n49, 
      dp_id_stage_regfile_DataPath_Physical_RF_n48, 
      dp_id_stage_regfile_DataPath_Physical_RF_n47, 
      dp_id_stage_regfile_DataPath_Physical_RF_n46, 
      dp_id_stage_regfile_DataPath_Physical_RF_n45, 
      dp_id_stage_regfile_DataPath_Physical_RF_n44, 
      dp_id_stage_regfile_DataPath_Physical_RF_n43, 
      dp_id_stage_regfile_DataPath_Physical_RF_n42, 
      dp_id_stage_regfile_DataPath_Physical_RF_n41, 
      dp_id_stage_regfile_DataPath_Physical_RF_n40, 
      dp_id_stage_regfile_DataPath_Physical_RF_n39, 
      dp_id_stage_regfile_DataPath_Physical_RF_n38, 
      dp_id_stage_regfile_DataPath_Physical_RF_n37, 
      dp_id_stage_regfile_DataPath_Physical_RF_n36, 
      dp_id_stage_regfile_DataPath_Physical_RF_n35, 
      dp_id_stage_regfile_DataPath_Physical_RF_n34, 
      dp_id_stage_regfile_DataPath_Physical_RF_n33, 
      dp_id_stage_regfile_DataPath_Physical_RF_n32, 
      dp_id_stage_regfile_DataPath_Physical_RF_n31, 
      dp_id_stage_regfile_DataPath_Physical_RF_n30, 
      dp_id_stage_regfile_DataPath_Physical_RF_n29, 
      dp_id_stage_regfile_DataPath_Physical_RF_n28, 
      dp_id_stage_regfile_DataPath_Physical_RF_n27, 
      dp_id_stage_regfile_DataPath_Physical_RF_n26, 
      dp_id_stage_regfile_DataPath_Physical_RF_n25, 
      dp_id_stage_regfile_DataPath_Physical_RF_n24, 
      dp_id_stage_regfile_DataPath_Physical_RF_n23, 
      dp_id_stage_regfile_DataPath_Physical_RF_n22, 
      dp_id_stage_regfile_DataPath_Physical_RF_n21, 
      dp_id_stage_regfile_DataPath_Physical_RF_n20, 
      dp_id_stage_regfile_DataPath_Physical_RF_n19, 
      dp_id_stage_regfile_DataPath_Physical_RF_n18, 
      dp_id_stage_regfile_DataPath_Physical_RF_n17, 
      dp_id_stage_regfile_DataPath_Physical_RF_n16, 
      dp_id_stage_regfile_DataPath_Physical_RF_n15, 
      dp_id_stage_regfile_DataPath_Physical_RF_n14, 
      dp_id_stage_regfile_DataPath_Physical_RF_n13, 
      dp_id_stage_regfile_DataPath_Physical_RF_n12, 
      dp_id_stage_regfile_DataPath_Physical_RF_n11, 
      dp_id_stage_regfile_DataPath_Physical_RF_n10, 
      dp_id_stage_regfile_DataPath_Physical_RF_n9, 
      dp_id_stage_regfile_DataPath_Physical_RF_n8, 
      dp_id_stage_regfile_DataPath_Physical_RF_n7, 
      dp_id_stage_regfile_DataPath_Physical_RF_n6, 
      dp_id_stage_regfile_DataPath_Physical_RF_n5, 
      dp_id_stage_regfile_DataPath_Physical_RF_n4, 
      dp_id_stage_regfile_DataPath_Physical_RF_n3, 
      dp_id_stage_regfile_DataPath_Physical_RF_n2, 
      dp_id_stage_regfile_DataPath_Physical_RF_N429_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N428_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N427_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N426_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N425_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N424_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N423_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N422_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N421_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N420_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N419_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N418_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N417_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N416_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N415_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N414_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N413_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N412_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N411_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N410_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N409_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N408_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N407_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N406_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N405_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N404_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N403_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N402_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N401_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N400_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N399_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N398_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N397_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N396_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N359_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N358_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N357_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N356_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N355_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N354_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N353_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N352_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N351_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N350_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N349_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N348_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N347_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N346_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N345_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N344_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N343_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N342_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N341_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N340_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N339_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N338_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N337_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N336_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N335_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N334_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N333_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N332_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N331_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N330_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N329_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_N328_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_31_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_0_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_1_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_2_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_3_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_4_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_5_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_6_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_7_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_8_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_9_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_10_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_11_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_12_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_13_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_14_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_15_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_16_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_17_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_18_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_19_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_20_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_21_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_22_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_23_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_24_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_25_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_26_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_27_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_28_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_29_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_30_port, 
      dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_31_port, 
      dp_ex_stage_n10, dp_ex_stage_n9, dp_ex_stage_n8, dp_ex_stage_n7, 
      dp_ex_stage_n6, dp_ex_stage_n5, dp_ex_stage_n4, dp_ex_stage_n3, 
      dp_ex_stage_n2, dp_ex_stage_n1, dp_ex_stage_muxB_out_0_port, 
      dp_ex_stage_muxB_out_1_port, dp_ex_stage_muxB_out_2_port, 
      dp_ex_stage_muxB_out_3_port, dp_ex_stage_muxB_out_4_port, 
      dp_ex_stage_muxB_out_5_port, dp_ex_stage_muxB_out_6_port, 
      dp_ex_stage_muxB_out_7_port, dp_ex_stage_muxB_out_8_port, 
      dp_ex_stage_muxB_out_9_port, dp_ex_stage_muxB_out_10_port, 
      dp_ex_stage_muxB_out_11_port, dp_ex_stage_muxB_out_12_port, 
      dp_ex_stage_muxB_out_13_port, dp_ex_stage_muxB_out_14_port, 
      dp_ex_stage_muxB_out_15_port, dp_ex_stage_muxB_out_16_port, 
      dp_ex_stage_muxB_out_17_port, dp_ex_stage_muxB_out_18_port, 
      dp_ex_stage_muxB_out_19_port, dp_ex_stage_muxB_out_20_port, 
      dp_ex_stage_muxB_out_21_port, dp_ex_stage_muxB_out_22_port, 
      dp_ex_stage_muxB_out_23_port, dp_ex_stage_muxB_out_24_port, 
      dp_ex_stage_muxB_out_25_port, dp_ex_stage_muxB_out_26_port, 
      dp_ex_stage_muxB_out_27_port, dp_ex_stage_muxB_out_28_port, 
      dp_ex_stage_muxB_out_29_port, dp_ex_stage_muxB_out_30_port, 
      dp_ex_stage_muxB_out_31_port, dp_ex_stage_muxA_out_0_port, 
      dp_ex_stage_muxA_out_1_port, dp_ex_stage_muxA_out_2_port, 
      dp_ex_stage_muxA_out_3_port, dp_ex_stage_muxA_out_4_port, 
      dp_ex_stage_muxA_out_5_port, dp_ex_stage_muxA_out_6_port, 
      dp_ex_stage_muxA_out_7_port, dp_ex_stage_muxA_out_8_port, 
      dp_ex_stage_muxA_out_9_port, dp_ex_stage_muxA_out_10_port, 
      dp_ex_stage_muxA_out_11_port, dp_ex_stage_muxA_out_12_port, 
      dp_ex_stage_muxA_out_13_port, dp_ex_stage_muxA_out_14_port, 
      dp_ex_stage_muxA_out_15_port, dp_ex_stage_muxA_out_16_port, 
      dp_ex_stage_muxA_out_17_port, dp_ex_stage_muxA_out_18_port, 
      dp_ex_stage_muxA_out_19_port, dp_ex_stage_muxA_out_20_port, 
      dp_ex_stage_muxA_out_21_port, dp_ex_stage_muxA_out_22_port, 
      dp_ex_stage_muxA_out_23_port, dp_ex_stage_muxA_out_24_port, 
      dp_ex_stage_muxA_out_25_port, dp_ex_stage_muxA_out_26_port, 
      dp_ex_stage_muxA_out_27_port, dp_ex_stage_muxA_out_28_port, 
      dp_ex_stage_muxA_out_29_port, dp_ex_stage_muxA_out_30_port, 
      dp_ex_stage_muxA_out_31_port, dp_ex_stage_muxA_n27, dp_ex_stage_muxA_n8, 
      dp_ex_stage_muxA_n7, dp_ex_stage_muxA_n6, dp_ex_stage_muxA_n5, 
      dp_ex_stage_muxA_n4, dp_ex_stage_muxA_n3, dp_ex_stage_muxA_n2, 
      dp_ex_stage_muxB_n8, dp_ex_stage_muxB_n7, dp_ex_stage_muxB_n6, 
      dp_ex_stage_muxB_n5, dp_ex_stage_muxB_n4, dp_ex_stage_muxB_n3, 
      dp_ex_stage_muxB_n2, dp_ex_stage_muxB_n1, dp_ex_stage_alu_n311, 
      dp_ex_stage_alu_n310, dp_ex_stage_alu_n309, dp_ex_stage_alu_n308, 
      dp_ex_stage_alu_n307, dp_ex_stage_alu_n306, dp_ex_stage_alu_n305, 
      dp_ex_stage_alu_n304, dp_ex_stage_alu_n303, dp_ex_stage_alu_n302, 
      dp_ex_stage_alu_n301, dp_ex_stage_alu_n300, dp_ex_stage_alu_n299, 
      dp_ex_stage_alu_n298, dp_ex_stage_alu_n297, dp_ex_stage_alu_n296, 
      dp_ex_stage_alu_n295, dp_ex_stage_alu_n294, dp_ex_stage_alu_n293, 
      dp_ex_stage_alu_n292, dp_ex_stage_alu_n291, dp_ex_stage_alu_n290, 
      dp_ex_stage_alu_n289, dp_ex_stage_alu_n288, dp_ex_stage_alu_n287, 
      dp_ex_stage_alu_n286, dp_ex_stage_alu_n285, dp_ex_stage_alu_n284, 
      dp_ex_stage_alu_n283, dp_ex_stage_alu_n282, dp_ex_stage_alu_n281, 
      dp_ex_stage_alu_n280, dp_ex_stage_alu_n279, dp_ex_stage_alu_n278, 
      dp_ex_stage_alu_n277, dp_ex_stage_alu_n276, dp_ex_stage_alu_n275, 
      dp_ex_stage_alu_n274, dp_ex_stage_alu_n273, dp_ex_stage_alu_n272, 
      dp_ex_stage_alu_n271, dp_ex_stage_alu_n270, dp_ex_stage_alu_n269, 
      dp_ex_stage_alu_n268, dp_ex_stage_alu_n267, dp_ex_stage_alu_n266, 
      dp_ex_stage_alu_n265, dp_ex_stage_alu_n264, dp_ex_stage_alu_n263, 
      dp_ex_stage_alu_n262, dp_ex_stage_alu_n261, dp_ex_stage_alu_n260, 
      dp_ex_stage_alu_n259, dp_ex_stage_alu_n258, dp_ex_stage_alu_n257, 
      dp_ex_stage_alu_n256, dp_ex_stage_alu_n255, dp_ex_stage_alu_n254, 
      dp_ex_stage_alu_n253, dp_ex_stage_alu_n252, dp_ex_stage_alu_n251, 
      dp_ex_stage_alu_n250, dp_ex_stage_alu_n249, dp_ex_stage_alu_n248, 
      dp_ex_stage_alu_n247, dp_ex_stage_alu_n246, dp_ex_stage_alu_n245, 
      dp_ex_stage_alu_n244, dp_ex_stage_alu_n243, dp_ex_stage_alu_n242, 
      dp_ex_stage_alu_n241, dp_ex_stage_alu_n240, dp_ex_stage_alu_n239, 
      dp_ex_stage_alu_n238, dp_ex_stage_alu_n237, dp_ex_stage_alu_n236, 
      dp_ex_stage_alu_n235, dp_ex_stage_alu_n234, dp_ex_stage_alu_n233, 
      dp_ex_stage_alu_n232, dp_ex_stage_alu_n231, dp_ex_stage_alu_n230, 
      dp_ex_stage_alu_n229, dp_ex_stage_alu_n228, dp_ex_stage_alu_n227, 
      dp_ex_stage_alu_n226, dp_ex_stage_alu_n225, dp_ex_stage_alu_n224, 
      dp_ex_stage_alu_n223, dp_ex_stage_alu_n222, dp_ex_stage_alu_n221, 
      dp_ex_stage_alu_n220, dp_ex_stage_alu_n219, dp_ex_stage_alu_n218, 
      dp_ex_stage_alu_n217, dp_ex_stage_alu_n216, dp_ex_stage_alu_n215, 
      dp_ex_stage_alu_n214, dp_ex_stage_alu_n213, dp_ex_stage_alu_n212, 
      dp_ex_stage_alu_n211, dp_ex_stage_alu_n210, dp_ex_stage_alu_n209, 
      dp_ex_stage_alu_n207, dp_ex_stage_alu_n204, dp_ex_stage_alu_n203, 
      dp_ex_stage_alu_n202, dp_ex_stage_alu_n201, dp_ex_stage_alu_n200, 
      dp_ex_stage_alu_n199, dp_ex_stage_alu_n198, dp_ex_stage_alu_n197, 
      dp_ex_stage_alu_n196, dp_ex_stage_alu_n195, dp_ex_stage_alu_n194, 
      dp_ex_stage_alu_n193, dp_ex_stage_alu_n192, dp_ex_stage_alu_n191, 
      dp_ex_stage_alu_n93, dp_ex_stage_alu_n92, dp_ex_stage_alu_n89, 
      dp_ex_stage_alu_n88, dp_ex_stage_alu_n87, dp_ex_stage_alu_n86, 
      dp_ex_stage_alu_n85, dp_ex_stage_alu_n84, dp_ex_stage_alu_n83, 
      dp_ex_stage_alu_n82, dp_ex_stage_alu_n81, dp_ex_stage_alu_n80, 
      dp_ex_stage_alu_n79, dp_ex_stage_alu_n78, dp_ex_stage_alu_n77, 
      dp_ex_stage_alu_n76, dp_ex_stage_alu_n74, dp_ex_stage_alu_n73, 
      dp_ex_stage_alu_n72, dp_ex_stage_alu_n71, dp_ex_stage_alu_n70, 
      dp_ex_stage_alu_n69, dp_ex_stage_alu_n68, dp_ex_stage_alu_n67, 
      dp_ex_stage_alu_n66, dp_ex_stage_alu_n65, dp_ex_stage_alu_n64, 
      dp_ex_stage_alu_n63, dp_ex_stage_alu_n62, dp_ex_stage_alu_n61, 
      dp_ex_stage_alu_n60, dp_ex_stage_alu_n59, dp_ex_stage_alu_n58, 
      dp_ex_stage_alu_n57, dp_ex_stage_alu_n56, dp_ex_stage_alu_n55, 
      dp_ex_stage_alu_n54, dp_ex_stage_alu_n53, dp_ex_stage_alu_n52, 
      dp_ex_stage_alu_n51, dp_ex_stage_alu_n50, dp_ex_stage_alu_n49, 
      dp_ex_stage_alu_n48, dp_ex_stage_alu_n47, dp_ex_stage_alu_n46, 
      dp_ex_stage_alu_n45, dp_ex_stage_alu_n44, dp_ex_stage_alu_n43, 
      dp_ex_stage_alu_n42, dp_ex_stage_alu_n41, dp_ex_stage_alu_n40, 
      dp_ex_stage_alu_n39, dp_ex_stage_alu_n38, dp_ex_stage_alu_n37, 
      dp_ex_stage_alu_n36, dp_ex_stage_alu_n35, dp_ex_stage_alu_n34, 
      dp_ex_stage_alu_n33, dp_ex_stage_alu_n32, dp_ex_stage_alu_n31, 
      dp_ex_stage_alu_n30, dp_ex_stage_alu_n29, dp_ex_stage_alu_n28, 
      dp_ex_stage_alu_n27, dp_ex_stage_alu_n26, dp_ex_stage_alu_n25, 
      dp_ex_stage_alu_n24, dp_ex_stage_alu_n23, dp_ex_stage_alu_n22, 
      dp_ex_stage_alu_n21, dp_ex_stage_alu_n20, dp_ex_stage_alu_n19, 
      dp_ex_stage_alu_n18, dp_ex_stage_alu_n17, dp_ex_stage_alu_n16, 
      dp_ex_stage_alu_n15, dp_ex_stage_alu_n14, dp_ex_stage_alu_n11, 
      dp_ex_stage_alu_n10, dp_ex_stage_alu_n9, dp_ex_stage_alu_n8, 
      dp_ex_stage_alu_n7, dp_ex_stage_alu_n6, dp_ex_stage_alu_n5, 
      dp_ex_stage_alu_n4, dp_ex_stage_alu_n3, dp_ex_stage_alu_n2, 
      dp_ex_stage_alu_n1, dp_ex_stage_alu_n208, dp_ex_stage_alu_n206, 
      dp_ex_stage_alu_n205, dp_ex_stage_alu_n190, dp_ex_stage_alu_n189, 
      dp_ex_stage_alu_n188, dp_ex_stage_alu_n187, dp_ex_stage_alu_n186, 
      dp_ex_stage_alu_n185, dp_ex_stage_alu_n184, dp_ex_stage_alu_n183, 
      dp_ex_stage_alu_n182, dp_ex_stage_alu_n181, dp_ex_stage_alu_n180, 
      dp_ex_stage_alu_n179, dp_ex_stage_alu_n178, dp_ex_stage_alu_n177, 
      dp_ex_stage_alu_n176, dp_ex_stage_alu_n175, dp_ex_stage_alu_n174, 
      dp_ex_stage_alu_n173, dp_ex_stage_alu_n172, dp_ex_stage_alu_n171, 
      dp_ex_stage_alu_n170, dp_ex_stage_alu_n169, dp_ex_stage_alu_n168, 
      dp_ex_stage_alu_n167, dp_ex_stage_alu_n166, dp_ex_stage_alu_n165, 
      dp_ex_stage_alu_n164, dp_ex_stage_alu_n163, dp_ex_stage_alu_n162, 
      dp_ex_stage_alu_n161, dp_ex_stage_alu_n160, dp_ex_stage_alu_n159, 
      dp_ex_stage_alu_n158, dp_ex_stage_alu_n157, dp_ex_stage_alu_n156, 
      dp_ex_stage_alu_n155, dp_ex_stage_alu_n154, dp_ex_stage_alu_n153, 
      dp_ex_stage_alu_n152, dp_ex_stage_alu_n151, dp_ex_stage_alu_n150, 
      dp_ex_stage_alu_n149, dp_ex_stage_alu_n148, dp_ex_stage_alu_n147, 
      dp_ex_stage_alu_n146, dp_ex_stage_alu_n145, dp_ex_stage_alu_n144, 
      dp_ex_stage_alu_n143, dp_ex_stage_alu_n142, dp_ex_stage_alu_n141, 
      dp_ex_stage_alu_n140, dp_ex_stage_alu_n139, dp_ex_stage_alu_n138, 
      dp_ex_stage_alu_n137, dp_ex_stage_alu_n136, dp_ex_stage_alu_n135, 
      dp_ex_stage_alu_n134, dp_ex_stage_alu_n133, dp_ex_stage_alu_n132, 
      dp_ex_stage_alu_n131, dp_ex_stage_alu_n130, dp_ex_stage_alu_n129, 
      dp_ex_stage_alu_n128, dp_ex_stage_alu_n127, dp_ex_stage_alu_n126, 
      dp_ex_stage_alu_n125, dp_ex_stage_alu_n124, dp_ex_stage_alu_n123, 
      dp_ex_stage_alu_n122, dp_ex_stage_alu_n121, dp_ex_stage_alu_n120, 
      dp_ex_stage_alu_n119, dp_ex_stage_alu_n118, dp_ex_stage_alu_n117, 
      dp_ex_stage_alu_n116, dp_ex_stage_alu_n115, dp_ex_stage_alu_n114, 
      dp_ex_stage_alu_n113, dp_ex_stage_alu_n112, dp_ex_stage_alu_n111, 
      dp_ex_stage_alu_n110, dp_ex_stage_alu_n109, dp_ex_stage_alu_n108, 
      dp_ex_stage_alu_n107, dp_ex_stage_alu_n106, dp_ex_stage_alu_n105, 
      dp_ex_stage_alu_n104, dp_ex_stage_alu_n103, dp_ex_stage_alu_n102, 
      dp_ex_stage_alu_n101, dp_ex_stage_alu_n100, dp_ex_stage_alu_n99, 
      dp_ex_stage_alu_n98, dp_ex_stage_alu_n97, dp_ex_stage_alu_n96, 
      dp_ex_stage_alu_n95, dp_ex_stage_alu_n94, dp_ex_stage_alu_n91, 
      dp_ex_stage_alu_n90, dp_ex_stage_alu_n13, dp_ex_stage_alu_n12, 
      dp_ex_stage_alu_N23_port, dp_ex_stage_alu_shifter_out_0_port, 
      dp_ex_stage_alu_shifter_out_1_port, dp_ex_stage_alu_shifter_out_2_port, 
      dp_ex_stage_alu_shifter_out_3_port, dp_ex_stage_alu_shifter_out_4_port, 
      dp_ex_stage_alu_shifter_out_5_port, dp_ex_stage_alu_shifter_out_6_port, 
      dp_ex_stage_alu_shifter_out_7_port, dp_ex_stage_alu_shifter_out_8_port, 
      dp_ex_stage_alu_shifter_out_9_port, dp_ex_stage_alu_shifter_out_10_port, 
      dp_ex_stage_alu_shifter_out_11_port, dp_ex_stage_alu_shifter_out_12_port,
      dp_ex_stage_alu_shifter_out_13_port, dp_ex_stage_alu_shifter_out_14_port,
      dp_ex_stage_alu_shifter_out_15_port, dp_ex_stage_alu_shifter_out_16_port,
      dp_ex_stage_alu_shifter_out_17_port, dp_ex_stage_alu_shifter_out_18_port,
      dp_ex_stage_alu_shifter_out_19_port, dp_ex_stage_alu_shifter_out_20_port,
      dp_ex_stage_alu_shifter_out_21_port, dp_ex_stage_alu_shifter_out_22_port,
      dp_ex_stage_alu_shifter_out_23_port, dp_ex_stage_alu_shifter_out_24_port,
      dp_ex_stage_alu_shifter_out_25_port, dp_ex_stage_alu_shifter_out_26_port,
      dp_ex_stage_alu_shifter_out_27_port, dp_ex_stage_alu_shifter_out_28_port,
      dp_ex_stage_alu_shifter_out_29_port, dp_ex_stage_alu_shifter_out_30_port,
      dp_ex_stage_alu_shifter_out_31_port, dp_ex_stage_alu_shift_arith_i, 
      dp_ex_stage_alu_N22_port, dp_ex_stage_alu_N21_port, 
      dp_ex_stage_alu_N20_port, dp_ex_stage_alu_N19_port, 
      dp_ex_stage_alu_N18_port, dp_ex_stage_alu_N17_port, 
      dp_ex_stage_alu_N16_port, dp_ex_stage_alu_adder_out_0_port, 
      dp_ex_stage_alu_adder_out_1_port, dp_ex_stage_alu_adder_out_2_port, 
      dp_ex_stage_alu_adder_out_3_port, dp_ex_stage_alu_adder_out_4_port, 
      dp_ex_stage_alu_adder_out_5_port, dp_ex_stage_alu_adder_out_6_port, 
      dp_ex_stage_alu_adder_out_7_port, dp_ex_stage_alu_adder_out_8_port, 
      dp_ex_stage_alu_adder_out_9_port, dp_ex_stage_alu_adder_out_10_port, 
      dp_ex_stage_alu_adder_out_11_port, dp_ex_stage_alu_adder_out_12_port, 
      dp_ex_stage_alu_adder_out_13_port, dp_ex_stage_alu_adder_out_14_port, 
      dp_ex_stage_alu_adder_out_15_port, dp_ex_stage_alu_adder_out_16_port, 
      dp_ex_stage_alu_adder_out_17_port, dp_ex_stage_alu_adder_out_18_port, 
      dp_ex_stage_alu_adder_out_19_port, dp_ex_stage_alu_adder_out_20_port, 
      dp_ex_stage_alu_adder_out_21_port, dp_ex_stage_alu_adder_out_22_port, 
      dp_ex_stage_alu_adder_out_23_port, dp_ex_stage_alu_adder_out_24_port, 
      dp_ex_stage_alu_adder_out_25_port, dp_ex_stage_alu_adder_out_26_port, 
      dp_ex_stage_alu_adder_out_27_port, dp_ex_stage_alu_adder_out_28_port, 
      dp_ex_stage_alu_adder_out_29_port, dp_ex_stage_alu_adder_out_30_port, 
      dp_ex_stage_alu_adder_out_31_port, dp_ex_stage_alu_Logic1_port, 
      dp_ex_stage_alu_adder_n23, dp_ex_stage_alu_adder_n22, 
      dp_ex_stage_alu_adder_n21, dp_ex_stage_alu_adder_n20, 
      dp_ex_stage_alu_adder_n19, dp_ex_stage_alu_adder_n18, 
      dp_ex_stage_alu_adder_n17, dp_ex_stage_alu_adder_n16, 
      dp_ex_stage_alu_adder_n15, dp_ex_stage_alu_adder_n14, 
      dp_ex_stage_alu_adder_n13, dp_ex_stage_alu_adder_n12, 
      dp_ex_stage_alu_adder_n11, dp_ex_stage_alu_adder_n10, 
      dp_ex_stage_alu_adder_n9, dp_ex_stage_alu_adder_n8, 
      dp_ex_stage_alu_adder_n7, dp_ex_stage_alu_adder_n6, 
      dp_ex_stage_alu_adder_n5, dp_ex_stage_alu_adder_n4, 
      dp_ex_stage_alu_adder_n3, dp_ex_stage_alu_adder_n2, 
      dp_ex_stage_alu_adder_n1, dp_ex_stage_alu_adder_carries_0_port, 
      dp_ex_stage_alu_adder_carries_1_port, 
      dp_ex_stage_alu_adder_carries_2_port, 
      dp_ex_stage_alu_adder_carries_3_port, 
      dp_ex_stage_alu_adder_carries_4_port, 
      dp_ex_stage_alu_adder_carries_5_port, 
      dp_ex_stage_alu_adder_carries_6_port, 
      dp_ex_stage_alu_adder_carries_7_port, dp_ex_stage_alu_adder_B_xor_0_port,
      dp_ex_stage_alu_adder_B_xor_1_port, dp_ex_stage_alu_adder_B_xor_2_port, 
      dp_ex_stage_alu_adder_B_xor_3_port, dp_ex_stage_alu_adder_B_xor_4_port, 
      dp_ex_stage_alu_adder_B_xor_6_port, dp_ex_stage_alu_adder_B_xor_8_port, 
      dp_ex_stage_alu_adder_B_xor_9_port, dp_ex_stage_alu_adder_B_xor_10_port, 
      dp_ex_stage_alu_adder_B_xor_11_port, dp_ex_stage_alu_adder_B_xor_12_port,
      dp_ex_stage_alu_adder_B_xor_13_port, dp_ex_stage_alu_adder_B_xor_14_port,
      dp_ex_stage_alu_adder_B_xor_16_port, dp_ex_stage_alu_adder_B_xor_17_port,
      dp_ex_stage_alu_adder_B_xor_18_port, dp_ex_stage_alu_adder_B_xor_19_port,
      dp_ex_stage_alu_adder_B_xor_20_port, dp_ex_stage_alu_adder_B_xor_21_port,
      dp_ex_stage_alu_adder_B_xor_22_port, dp_ex_stage_alu_adder_B_xor_23_port,
      dp_ex_stage_alu_adder_B_xor_24_port, dp_ex_stage_alu_adder_B_xor_25_port,
      dp_ex_stage_alu_adder_B_xor_26_port, dp_ex_stage_alu_adder_B_xor_27_port,
      dp_ex_stage_alu_adder_B_xor_28_port, dp_ex_stage_alu_adder_B_xor_29_port,
      dp_ex_stage_alu_adder_B_xor_30_port, dp_ex_stage_alu_adder_B_xor_31_port,
      dp_ex_stage_alu_adder_Cout, dp_ex_stage_alu_adder_SparseTree_n4, 
      dp_ex_stage_alu_adder_SparseTree_n3, dp_ex_stage_alu_adder_SparseTree_n1,
      dp_ex_stage_alu_adder_SparseTree_prop_2_2_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_3_3_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_4_3_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_4_4_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_5_5_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_6_5_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_6_6_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_7_7_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_8_5_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_8_7_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_8_8_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_9_9_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_10_9_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_10_10_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_11_11_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_12_9_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_12_11_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_12_12_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_13_13_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_14_13_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_14_14_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_15_15_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_16_9_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_16_13_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_16_15_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_16_16_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_17_17_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_18_17_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_18_18_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_19_19_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_20_17_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_20_19_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_20_20_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_21_21_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_22_21_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_22_22_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_23_23_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_24_17_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_24_21_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_24_23_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_24_24_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_25_25_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_26_25_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_26_26_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_27_27_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_28_17_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_28_25_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_28_27_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_28_28_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_29_29_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_30_29_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_30_30_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_31_31_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_32_17_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_32_25_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_32_29_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_32_31_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_32_32_port, 
      dp_ex_stage_alu_adder_SparseTree_prop_1_1_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_2_0_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_2_2_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_3_3_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_4_3_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_4_4_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_5_5_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_6_5_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_6_6_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_7_7_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_8_5_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_8_7_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_8_8_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_9_9_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_10_9_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_10_10_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_11_11_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_12_9_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_12_11_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_12_12_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_13_13_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_14_13_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_14_14_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_15_15_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_16_9_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_16_13_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_16_15_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_16_16_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_17_17_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_18_17_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_18_18_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_19_19_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_20_17_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_20_19_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_20_20_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_21_21_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_22_21_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_22_22_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_23_23_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_24_17_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_24_21_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_24_23_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_24_24_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_25_25_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_26_25_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_26_26_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_27_27_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_28_17_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_28_25_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_28_27_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_28_28_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_29_29_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_30_29_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_30_30_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_31_31_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_32_17_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_32_25_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_32_29_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_32_31_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_32_32_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_1_0_port, 
      dp_ex_stage_alu_adder_SparseTree_gen_1_1_port, 
      dp_ex_stage_alu_adder_SparseTree_n9, dp_ex_stage_alu_adder_SparseTree_n8,
      dp_ex_stage_alu_adder_SparseTree_n7, 
      dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_n1, 
      dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_n1, 
      dp_ex_stage_alu_adder_SparseTree_G10_n2, 
      dp_ex_stage_alu_adder_SparseTree_G20_1_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_n2, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_n3, 
      dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_n3, 
      dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_n3, 
      dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_n3, 
      dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_n3, 
      dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_n3, 
      dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_n3, 
      dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_n3, 
      dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_n3, 
      dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_n3, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Logic0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Logic1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n9, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n8, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n7, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n6, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Logic0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Logic1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n13, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n12, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n11, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n10, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Logic0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Logic1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n13, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n12, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n11, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n10, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Logic0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Logic1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n13, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n12, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n11, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n10, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Logic0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Logic1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n13, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n12, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n11, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n10, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Logic0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Logic1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n14, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n13, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n12, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n11, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n10, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n1, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Logic0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Logic1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n4, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n3, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n2, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n1, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n14, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n13, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n12, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n11, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n10, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n1, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Logic0_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Logic1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_3_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_2_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_1_port, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_Co, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n14, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n13, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n12, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n11, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n10, 
      dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n1, dp_ex_stage_alu_shifter_n118
      , dp_ex_stage_alu_shifter_n117, dp_ex_stage_alu_shifter_n116, 
      dp_ex_stage_alu_shifter_n115, dp_ex_stage_alu_shifter_n114, 
      dp_ex_stage_alu_shifter_n113, dp_ex_stage_alu_shifter_n112, 
      dp_ex_stage_alu_shifter_n111, dp_ex_stage_alu_shifter_n110, 
      dp_ex_stage_alu_shifter_n109, dp_ex_stage_alu_shifter_n108, 
      dp_ex_stage_alu_shifter_n107, dp_ex_stage_alu_shifter_n106, 
      dp_ex_stage_alu_shifter_n105, dp_ex_stage_alu_shifter_n104, 
      dp_ex_stage_alu_shifter_n103, dp_ex_stage_alu_shifter_n102, 
      dp_ex_stage_alu_shifter_n101, dp_ex_stage_alu_shifter_n100, 
      dp_ex_stage_alu_shifter_n99, dp_ex_stage_alu_shifter_n98, 
      dp_ex_stage_alu_shifter_n97, dp_ex_stage_alu_shifter_n96, 
      dp_ex_stage_alu_shifter_n95, dp_ex_stage_alu_shifter_n94, 
      dp_ex_stage_alu_shifter_n93, dp_ex_stage_alu_shifter_n20, 
      dp_ex_stage_alu_shifter_n19, dp_ex_stage_alu_shifter_n12, 
      dp_ex_stage_alu_shifter_n11, dp_ex_stage_alu_shifter_n10, 
      dp_ex_stage_alu_shifter_n9, dp_ex_stage_alu_shifter_n8, 
      dp_ex_stage_alu_shifter_n7, dp_ex_stage_alu_shifter_n6, 
      dp_ex_stage_alu_shifter_n5, dp_ex_stage_alu_shifter_n4, 
      dp_ex_stage_alu_shifter_n3, dp_ex_stage_alu_shifter_n2, 
      dp_ex_stage_alu_shifter_n1, dp_ex_stage_alu_shifter_n92, 
      dp_ex_stage_alu_shifter_n91, dp_ex_stage_alu_shifter_n90, 
      dp_ex_stage_alu_shifter_n89, dp_ex_stage_alu_shifter_n88, 
      dp_ex_stage_alu_shifter_n87, dp_ex_stage_alu_shifter_n86, 
      dp_ex_stage_alu_shifter_n85, dp_ex_stage_alu_shifter_n84, 
      dp_ex_stage_alu_shifter_n83, dp_ex_stage_alu_shifter_n82, 
      dp_ex_stage_alu_shifter_n81, dp_ex_stage_alu_shifter_n80, 
      dp_ex_stage_alu_shifter_n79, dp_ex_stage_alu_shifter_n78, 
      dp_ex_stage_alu_shifter_n77, dp_ex_stage_alu_shifter_n76, 
      dp_ex_stage_alu_shifter_n75, dp_ex_stage_alu_shifter_n74, 
      dp_ex_stage_alu_shifter_n73, dp_ex_stage_alu_shifter_n72, 
      dp_ex_stage_alu_shifter_n71, dp_ex_stage_alu_shifter_n70, 
      dp_ex_stage_alu_shifter_n69, dp_ex_stage_alu_shifter_n68, 
      dp_ex_stage_alu_shifter_n67, dp_ex_stage_alu_shifter_n66, 
      dp_ex_stage_alu_shifter_n65, dp_ex_stage_alu_shifter_n64, 
      dp_ex_stage_alu_shifter_n63, dp_ex_stage_alu_shifter_n62, 
      dp_ex_stage_alu_shifter_n61, dp_ex_stage_alu_shifter_n60, 
      dp_ex_stage_alu_shifter_n59, dp_ex_stage_alu_shifter_n58, 
      dp_ex_stage_alu_shifter_n57, dp_ex_stage_alu_shifter_n56, 
      dp_ex_stage_alu_shifter_n55, dp_ex_stage_alu_shifter_n54, 
      dp_ex_stage_alu_shifter_n53, dp_ex_stage_alu_shifter_n52, 
      dp_ex_stage_alu_shifter_n51, dp_ex_stage_alu_shifter_n50, 
      dp_ex_stage_alu_shifter_n49, dp_ex_stage_alu_shifter_n48, 
      dp_ex_stage_alu_shifter_n47, dp_ex_stage_alu_shifter_n46, 
      dp_ex_stage_alu_shifter_n45, dp_ex_stage_alu_shifter_n44, 
      dp_ex_stage_alu_shifter_n43, dp_ex_stage_alu_shifter_n42, 
      dp_ex_stage_alu_shifter_n41, dp_ex_stage_alu_shifter_n40, 
      dp_ex_stage_alu_shifter_n39, dp_ex_stage_alu_shifter_n38, 
      dp_ex_stage_alu_shifter_n37, dp_ex_stage_alu_shifter_n36, 
      dp_ex_stage_alu_shifter_n35, dp_ex_stage_alu_shifter_n34, 
      dp_ex_stage_alu_shifter_n33, dp_ex_stage_alu_shifter_n32, 
      dp_ex_stage_alu_shifter_n31, dp_ex_stage_alu_shifter_n30, 
      dp_ex_stage_alu_shifter_n29, dp_ex_stage_alu_shifter_n28, 
      dp_ex_stage_alu_shifter_n27, dp_ex_stage_alu_shifter_n26, 
      dp_ex_stage_alu_shifter_n25, dp_ex_stage_alu_shifter_n24, 
      dp_ex_stage_alu_shifter_n23, dp_ex_stage_alu_shifter_n22, 
      dp_ex_stage_alu_shifter_n21, dp_ex_stage_alu_shifter_n18, 
      dp_ex_stage_alu_shifter_n17, dp_ex_stage_alu_shifter_n16, 
      dp_ex_stage_alu_shifter_n15, dp_ex_stage_alu_shifter_n14, 
      dp_ex_stage_alu_shifter_n13, dp_ex_stage_alu_shifter_N265, 
      dp_ex_stage_alu_shifter_N264, dp_ex_stage_alu_shifter_N263, 
      dp_ex_stage_alu_shifter_N262, dp_ex_stage_alu_shifter_N261, 
      dp_ex_stage_alu_shifter_N260, dp_ex_stage_alu_shifter_N259, 
      dp_ex_stage_alu_shifter_N258, dp_ex_stage_alu_shifter_N257, 
      dp_ex_stage_alu_shifter_N256, dp_ex_stage_alu_shifter_N255, 
      dp_ex_stage_alu_shifter_N254, dp_ex_stage_alu_shifter_N253, 
      dp_ex_stage_alu_shifter_N252, dp_ex_stage_alu_shifter_N251, 
      dp_ex_stage_alu_shifter_N250, dp_ex_stage_alu_shifter_N249, 
      dp_ex_stage_alu_shifter_N248, dp_ex_stage_alu_shifter_N247, 
      dp_ex_stage_alu_shifter_N246, dp_ex_stage_alu_shifter_N245, 
      dp_ex_stage_alu_shifter_N244, dp_ex_stage_alu_shifter_N243, 
      dp_ex_stage_alu_shifter_N242, dp_ex_stage_alu_shifter_N241, 
      dp_ex_stage_alu_shifter_N240, dp_ex_stage_alu_shifter_N239, 
      dp_ex_stage_alu_shifter_N238, dp_ex_stage_alu_shifter_N237, 
      dp_ex_stage_alu_shifter_N236, dp_ex_stage_alu_shifter_N235, 
      dp_ex_stage_alu_shifter_N234, dp_ex_stage_alu_shifter_N233, 
      dp_ex_stage_alu_shifter_N232, dp_ex_stage_alu_shifter_N231, 
      dp_ex_stage_alu_shifter_N230, dp_ex_stage_alu_shifter_N229, 
      dp_ex_stage_alu_shifter_N228, dp_ex_stage_alu_shifter_N227, 
      dp_ex_stage_alu_shifter_N226, dp_ex_stage_alu_shifter_N225, 
      dp_ex_stage_alu_shifter_N224, dp_ex_stage_alu_shifter_N223, 
      dp_ex_stage_alu_shifter_N222, dp_ex_stage_alu_shifter_N221, 
      dp_ex_stage_alu_shifter_N220, dp_ex_stage_alu_shifter_N219, 
      dp_ex_stage_alu_shifter_N218, dp_ex_stage_alu_shifter_N217, 
      dp_ex_stage_alu_shifter_N216, dp_ex_stage_alu_shifter_N215, 
      dp_ex_stage_alu_shifter_N214, dp_ex_stage_alu_shifter_N213, 
      dp_ex_stage_alu_shifter_N212, dp_ex_stage_alu_shifter_N211, 
      dp_ex_stage_alu_shifter_N210, dp_ex_stage_alu_shifter_N209, 
      dp_ex_stage_alu_shifter_N208, dp_ex_stage_alu_shifter_N207, 
      dp_ex_stage_alu_shifter_N206, dp_ex_stage_alu_shifter_N205, 
      dp_ex_stage_alu_shifter_N204, dp_ex_stage_alu_shifter_N203, 
      dp_ex_stage_alu_shifter_N202, dp_ex_stage_alu_shifter_N168, 
      dp_ex_stage_alu_shifter_N167, dp_ex_stage_alu_shifter_N166, 
      dp_ex_stage_alu_shifter_N165, dp_ex_stage_alu_shifter_N164, 
      dp_ex_stage_alu_shifter_N163, dp_ex_stage_alu_shifter_N162, 
      dp_ex_stage_alu_shifter_N161, dp_ex_stage_alu_shifter_N160, 
      dp_ex_stage_alu_shifter_N159, dp_ex_stage_alu_shifter_N158, 
      dp_ex_stage_alu_shifter_N157, dp_ex_stage_alu_shifter_N156, 
      dp_ex_stage_alu_shifter_N155, dp_ex_stage_alu_shifter_N154, 
      dp_ex_stage_alu_shifter_N153, dp_ex_stage_alu_shifter_N152, 
      dp_ex_stage_alu_shifter_N151, dp_ex_stage_alu_shifter_N150, 
      dp_ex_stage_alu_shifter_N149, dp_ex_stage_alu_shifter_N148, 
      dp_ex_stage_alu_shifter_N147, dp_ex_stage_alu_shifter_N146, 
      dp_ex_stage_alu_shifter_N145, dp_ex_stage_alu_shifter_N144, 
      dp_ex_stage_alu_shifter_N143, dp_ex_stage_alu_shifter_N142, 
      dp_ex_stage_alu_shifter_N141, dp_ex_stage_alu_shifter_N140, 
      dp_ex_stage_alu_shifter_N139, dp_ex_stage_alu_shifter_N138, 
      dp_ex_stage_alu_shifter_N137, dp_ex_stage_alu_shifter_N136, 
      dp_ex_stage_alu_shifter_N135, dp_ex_stage_alu_shifter_N134, 
      dp_ex_stage_alu_shifter_N133, dp_ex_stage_alu_shifter_N132, 
      dp_ex_stage_alu_shifter_N131, dp_ex_stage_alu_shifter_N130, 
      dp_ex_stage_alu_shifter_N129, dp_ex_stage_alu_shifter_N128, 
      dp_ex_stage_alu_shifter_N127, dp_ex_stage_alu_shifter_N126, 
      dp_ex_stage_alu_shifter_N125, dp_ex_stage_alu_shifter_N124, 
      dp_ex_stage_alu_shifter_N123, dp_ex_stage_alu_shifter_N122, 
      dp_ex_stage_alu_shifter_N121, dp_ex_stage_alu_shifter_N120, 
      dp_ex_stage_alu_shifter_N119, dp_ex_stage_alu_shifter_N118_port, 
      dp_ex_stage_alu_shifter_N117_port, dp_ex_stage_alu_shifter_N116_port, 
      dp_ex_stage_alu_shifter_N115_port, dp_ex_stage_alu_shifter_N114_port, 
      dp_ex_stage_alu_shifter_N113_port, dp_ex_stage_alu_shifter_N112_port, 
      dp_ex_stage_alu_shifter_N111_port, dp_ex_stage_alu_shifter_N110_port, 
      dp_ex_stage_alu_shifter_N109_port, dp_ex_stage_alu_shifter_N108_port, 
      dp_ex_stage_alu_shifter_N107_port, dp_ex_stage_alu_shifter_N106_port, 
      dp_ex_stage_alu_shifter_N105_port, dp_ex_stage_alu_shifter_N70_port, 
      dp_ex_stage_alu_shifter_N69_port, dp_ex_stage_alu_shifter_N68_port, 
      dp_ex_stage_alu_shifter_N67_port, dp_ex_stage_alu_shifter_N66_port, 
      dp_ex_stage_alu_shifter_N65_port, dp_ex_stage_alu_shifter_N64_port, 
      dp_ex_stage_alu_shifter_N63_port, dp_ex_stage_alu_shifter_N62_port, 
      dp_ex_stage_alu_shifter_N61_port, dp_ex_stage_alu_shifter_N60_port, 
      dp_ex_stage_alu_shifter_N59_port, dp_ex_stage_alu_shifter_N58_port, 
      dp_ex_stage_alu_shifter_N57_port, dp_ex_stage_alu_shifter_N56_port, 
      dp_ex_stage_alu_shifter_N55_port, dp_ex_stage_alu_shifter_N54_port, 
      dp_ex_stage_alu_shifter_N53_port, dp_ex_stage_alu_shifter_N52_port, 
      dp_ex_stage_alu_shifter_N51_port, dp_ex_stage_alu_shifter_N50_port, 
      dp_ex_stage_alu_shifter_N49_port, dp_ex_stage_alu_shifter_N48_port, 
      dp_ex_stage_alu_shifter_N47_port, dp_ex_stage_alu_shifter_N46_port, 
      dp_ex_stage_alu_shifter_N45_port, dp_ex_stage_alu_shifter_N44_port, 
      dp_ex_stage_alu_shifter_N43_port, dp_ex_stage_alu_shifter_N42_port, 
      dp_ex_stage_alu_shifter_N41_port, dp_ex_stage_alu_shifter_N40_port, 
      dp_ex_stage_alu_shifter_N39_port, dp_ex_stage_alu_shifter_N38_port, 
      dp_ex_stage_alu_shifter_N37_port, dp_ex_stage_alu_shifter_N36_port, 
      dp_ex_stage_alu_shifter_N35_port, dp_ex_stage_alu_shifter_N34_port, 
      dp_ex_stage_alu_shifter_N33_port, dp_ex_stage_alu_shifter_N32_port, 
      dp_ex_stage_alu_shifter_N31_port, dp_ex_stage_alu_shifter_N30_port, 
      dp_ex_stage_alu_shifter_N29_port, dp_ex_stage_alu_shifter_N28_port, 
      dp_ex_stage_alu_shifter_N27_port, dp_ex_stage_alu_shifter_N26_port, 
      dp_ex_stage_alu_shifter_N25_port, dp_ex_stage_alu_shifter_N24_port, 
      dp_ex_stage_alu_shifter_N23_port, dp_ex_stage_alu_shifter_N22_port, 
      dp_ex_stage_alu_shifter_N21_port, dp_ex_stage_alu_shifter_N20_port, 
      dp_ex_stage_alu_shifter_N19_port, dp_ex_stage_alu_shifter_N18_port, 
      dp_ex_stage_alu_shifter_N17_port, dp_ex_stage_alu_shifter_N16_port, 
      dp_ex_stage_alu_shifter_N15_port, dp_ex_stage_alu_shifter_N14_port, 
      dp_ex_stage_alu_shifter_N13_port, dp_ex_stage_alu_shifter_N12_port, 
      dp_ex_stage_alu_shifter_N11_port, dp_ex_stage_alu_shifter_N10_port, 
      dp_ex_stage_alu_shifter_N9_port, dp_ex_stage_alu_shifter_N8_port, 
      dp_ex_stage_alu_shifter_N7_port, dp_ex_stage_alu_shifter_sll_48_n34, 
      dp_ex_stage_alu_shifter_sll_48_n33, dp_ex_stage_alu_shifter_sll_48_n32, 
      dp_ex_stage_alu_shifter_sll_48_n31, dp_ex_stage_alu_shifter_sll_48_n30, 
      dp_ex_stage_alu_shifter_sll_48_n29, dp_ex_stage_alu_shifter_sll_48_n28, 
      dp_ex_stage_alu_shifter_sll_48_n27, dp_ex_stage_alu_shifter_sll_48_n26, 
      dp_ex_stage_alu_shifter_sll_48_n25, dp_ex_stage_alu_shifter_sll_48_n24, 
      dp_ex_stage_alu_shifter_sll_48_n23, dp_ex_stage_alu_shifter_sll_48_n22, 
      dp_ex_stage_alu_shifter_sll_48_n21, dp_ex_stage_alu_shifter_sll_48_n20, 
      dp_ex_stage_alu_shifter_sll_48_n19, dp_ex_stage_alu_shifter_sll_48_n18, 
      dp_ex_stage_alu_shifter_sll_48_n17, dp_ex_stage_alu_shifter_sll_48_n16, 
      dp_ex_stage_alu_shifter_sll_48_n15, dp_ex_stage_alu_shifter_sll_48_n14, 
      dp_ex_stage_alu_shifter_sll_48_n13, dp_ex_stage_alu_shifter_sll_48_n12, 
      dp_ex_stage_alu_shifter_sll_48_n11, dp_ex_stage_alu_shifter_sll_48_n10, 
      dp_ex_stage_alu_shifter_sll_48_n9, dp_ex_stage_alu_shifter_sll_48_n8, 
      dp_ex_stage_alu_shifter_sll_48_n7, dp_ex_stage_alu_shifter_sll_48_n6, 
      dp_ex_stage_alu_shifter_sll_48_n5, dp_ex_stage_alu_shifter_sll_48_n4, 
      dp_ex_stage_alu_shifter_sll_48_n3, dp_ex_stage_alu_shifter_sll_48_n2, 
      dp_ex_stage_alu_shifter_sll_48_n1, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_8_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_9_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_10_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_11_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_12_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_13_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_14_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_15_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_16_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_17_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_18_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_19_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_20_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_21_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_22_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_23_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_24_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_25_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_26_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_27_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_28_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_29_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_30_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_4_31_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_0_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_1_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_2_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_3_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_4_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_5_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_6_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_7_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_8_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_9_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_10_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_11_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_12_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_13_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_14_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_15_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_16_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_17_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_18_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_19_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_20_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_21_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_22_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_23_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_24_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_25_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_26_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_27_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_28_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_29_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_30_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_3_31_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_0_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_1_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_2_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_3_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_4_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_5_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_6_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_7_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_8_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_9_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_10_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_11_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_12_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_13_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_14_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_15_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_16_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_17_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_18_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_19_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_20_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_21_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_22_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_23_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_24_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_25_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_26_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_27_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_28_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_29_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_30_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_2_31_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_0_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_1_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_2_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_3_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_4_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_5_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_6_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_7_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_8_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_9_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_10_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_11_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_12_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_13_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_14_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_15_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_16_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_17_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_18_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_19_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_20_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_21_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_22_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_23_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_24_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_25_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_26_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_27_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_28_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_29_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_30_port, 
      dp_ex_stage_alu_shifter_sll_48_ML_int_1_31_port, 
      dp_ex_stage_alu_shifter_sla_46_n193, dp_ex_stage_alu_shifter_sla_46_n192,
      dp_ex_stage_alu_shifter_sla_46_n191, dp_ex_stage_alu_shifter_sla_46_n190,
      dp_ex_stage_alu_shifter_sla_46_n189, dp_ex_stage_alu_shifter_sla_46_n188,
      dp_ex_stage_alu_shifter_sla_46_n187, dp_ex_stage_alu_shifter_sla_46_n186,
      dp_ex_stage_alu_shifter_sla_46_n185, dp_ex_stage_alu_shifter_sla_46_n184,
      dp_ex_stage_alu_shifter_sla_46_n183, dp_ex_stage_alu_shifter_sla_46_n182,
      dp_ex_stage_alu_shifter_sla_46_n181, dp_ex_stage_alu_shifter_sla_46_n180,
      dp_ex_stage_alu_shifter_sla_46_n179, dp_ex_stage_alu_shifter_sla_46_n178,
      dp_ex_stage_alu_shifter_sla_46_n177, dp_ex_stage_alu_shifter_sla_46_n176,
      dp_ex_stage_alu_shifter_sla_46_n175, dp_ex_stage_alu_shifter_sla_46_n174,
      dp_ex_stage_alu_shifter_sla_46_n173, dp_ex_stage_alu_shifter_sla_46_n172,
      dp_ex_stage_alu_shifter_sla_46_n171, dp_ex_stage_alu_shifter_sla_46_n170,
      dp_ex_stage_alu_shifter_sla_46_n169, dp_ex_stage_alu_shifter_sla_46_n168,
      dp_ex_stage_alu_shifter_sla_46_n167, dp_ex_stage_alu_shifter_sla_46_n166,
      dp_ex_stage_alu_shifter_sla_46_n165, dp_ex_stage_alu_shifter_sla_46_n164,
      dp_ex_stage_alu_shifter_sla_46_n163, dp_ex_stage_alu_shifter_sla_46_n162,
      dp_ex_stage_alu_shifter_sla_46_n161, dp_ex_stage_alu_shifter_sla_46_n160,
      dp_ex_stage_alu_shifter_sla_46_n159, dp_ex_stage_alu_shifter_sla_46_n158,
      dp_ex_stage_alu_shifter_sla_46_n157, dp_ex_stage_alu_shifter_sla_46_n156,
      dp_ex_stage_alu_shifter_sla_46_n155, dp_ex_stage_alu_shifter_sla_46_n154,
      dp_ex_stage_alu_shifter_sla_46_n153, dp_ex_stage_alu_shifter_sla_46_n152,
      dp_ex_stage_alu_shifter_sla_46_n151, dp_ex_stage_alu_shifter_sla_46_n150,
      dp_ex_stage_alu_shifter_sla_46_n149, dp_ex_stage_alu_shifter_sla_46_n148,
      dp_ex_stage_alu_shifter_sla_46_n147, dp_ex_stage_alu_shifter_sla_46_n146,
      dp_ex_stage_alu_shifter_sla_46_n145, dp_ex_stage_alu_shifter_sla_46_n144,
      dp_ex_stage_alu_shifter_sla_46_n143, dp_ex_stage_alu_shifter_sla_46_n142,
      dp_ex_stage_alu_shifter_sla_46_n141, dp_ex_stage_alu_shifter_sla_46_n140,
      dp_ex_stage_alu_shifter_sla_46_n139, dp_ex_stage_alu_shifter_sla_46_n138,
      dp_ex_stage_alu_shifter_sla_46_n137, dp_ex_stage_alu_shifter_sla_46_n136,
      dp_ex_stage_alu_shifter_sla_46_n135, dp_ex_stage_alu_shifter_sla_46_n134,
      dp_ex_stage_alu_shifter_sla_46_n133, dp_ex_stage_alu_shifter_sla_46_n132,
      dp_ex_stage_alu_shifter_sla_46_n131, dp_ex_stage_alu_shifter_sla_46_n130,
      dp_ex_stage_alu_shifter_sla_46_n129, dp_ex_stage_alu_shifter_sla_46_n128,
      dp_ex_stage_alu_shifter_sla_46_n127, dp_ex_stage_alu_shifter_sla_46_n126,
      dp_ex_stage_alu_shifter_sla_46_n125, dp_ex_stage_alu_shifter_sla_46_n124,
      dp_ex_stage_alu_shifter_sla_46_n123, dp_ex_stage_alu_shifter_sla_46_n122,
      dp_ex_stage_alu_shifter_sla_46_n121, dp_ex_stage_alu_shifter_sla_46_n120,
      dp_ex_stage_alu_shifter_sla_46_n119, dp_ex_stage_alu_shifter_sla_46_n118,
      dp_ex_stage_alu_shifter_sla_46_n117, dp_ex_stage_alu_shifter_sla_46_n116,
      dp_ex_stage_alu_shifter_sla_46_n115, dp_ex_stage_alu_shifter_sla_46_n114,
      dp_ex_stage_alu_shifter_sla_46_n113, dp_ex_stage_alu_shifter_sla_46_n112,
      dp_ex_stage_alu_shifter_sla_46_n111, dp_ex_stage_alu_shifter_sla_46_n110,
      dp_ex_stage_alu_shifter_sla_46_n109, dp_ex_stage_alu_shifter_sla_46_n108,
      dp_ex_stage_alu_shifter_sla_46_n107, dp_ex_stage_alu_shifter_sla_46_n106,
      dp_ex_stage_alu_shifter_sla_46_n105, dp_ex_stage_alu_shifter_sla_46_n104,
      dp_ex_stage_alu_shifter_sla_46_n103, dp_ex_stage_alu_shifter_sla_46_n102,
      dp_ex_stage_alu_shifter_sla_46_n101, dp_ex_stage_alu_shifter_sla_46_n100,
      dp_ex_stage_alu_shifter_sla_46_n99, dp_ex_stage_alu_shifter_sla_46_n98, 
      dp_ex_stage_alu_shifter_sla_46_n97, dp_ex_stage_alu_shifter_sla_46_n96, 
      dp_ex_stage_alu_shifter_sla_46_n95, dp_ex_stage_alu_shifter_sla_46_n94, 
      dp_ex_stage_alu_shifter_sla_46_n93, dp_ex_stage_alu_shifter_sla_46_n92, 
      dp_ex_stage_alu_shifter_sla_46_n91, dp_ex_stage_alu_shifter_sla_46_n90, 
      dp_ex_stage_alu_shifter_sla_46_n89, dp_ex_stage_alu_shifter_sla_46_n88, 
      dp_ex_stage_alu_shifter_sla_46_n87, dp_ex_stage_alu_shifter_sla_46_n86, 
      dp_ex_stage_alu_shifter_sla_46_n85, dp_ex_stage_alu_shifter_sla_46_n84, 
      dp_ex_stage_alu_shifter_sla_46_n83, dp_ex_stage_alu_shifter_sla_46_n82, 
      dp_ex_stage_alu_shifter_sla_46_n81, dp_ex_stage_alu_shifter_sla_46_n80, 
      dp_ex_stage_alu_shifter_sla_46_n79, dp_ex_stage_alu_shifter_sla_46_n78, 
      dp_ex_stage_alu_shifter_sla_46_n77, dp_ex_stage_alu_shifter_sla_46_n76, 
      dp_ex_stage_alu_shifter_sla_46_n75, dp_ex_stage_alu_shifter_sla_46_n74, 
      dp_ex_stage_alu_shifter_sla_46_n73, dp_ex_stage_alu_shifter_sla_46_n72, 
      dp_ex_stage_alu_shifter_sla_46_n71, dp_ex_stage_alu_shifter_sla_46_n70, 
      dp_ex_stage_alu_shifter_sla_46_n69, dp_ex_stage_alu_shifter_sla_46_n68, 
      dp_ex_stage_alu_shifter_sla_46_n67, dp_ex_stage_alu_shifter_sla_46_n66, 
      dp_ex_stage_alu_shifter_sla_46_n65, dp_ex_stage_alu_shifter_sla_46_n64, 
      dp_ex_stage_alu_shifter_sla_46_n63, dp_ex_stage_alu_shifter_sla_46_n62, 
      dp_ex_stage_alu_shifter_sla_46_n61, dp_ex_stage_alu_shifter_sla_46_n60, 
      dp_ex_stage_alu_shifter_sla_46_n59, dp_ex_stage_alu_shifter_sla_46_n58, 
      dp_ex_stage_alu_shifter_sla_46_n57, dp_ex_stage_alu_shifter_sla_46_n56, 
      dp_ex_stage_alu_shifter_sla_46_n55, dp_ex_stage_alu_shifter_sla_46_n54, 
      dp_ex_stage_alu_shifter_sla_46_n53, dp_ex_stage_alu_shifter_sla_46_n52, 
      dp_ex_stage_alu_shifter_sla_46_n51, dp_ex_stage_alu_shifter_sla_46_n50, 
      dp_ex_stage_alu_shifter_sla_46_n49, dp_ex_stage_alu_shifter_sla_46_n48, 
      dp_ex_stage_alu_shifter_sla_46_n47, dp_ex_stage_alu_shifter_sla_46_n46, 
      dp_ex_stage_alu_shifter_sla_46_n45, dp_ex_stage_alu_shifter_sla_46_n44, 
      dp_ex_stage_alu_shifter_sla_46_n43, dp_ex_stage_alu_shifter_sla_46_n42, 
      dp_ex_stage_alu_shifter_sla_46_n41, dp_ex_stage_alu_shifter_sla_46_n40, 
      dp_ex_stage_alu_shifter_sla_46_n39, dp_ex_stage_alu_shifter_sla_46_n38, 
      dp_ex_stage_alu_shifter_sla_46_n37, dp_ex_stage_alu_shifter_sla_46_n36, 
      dp_ex_stage_alu_shifter_sla_46_n35, dp_ex_stage_alu_shifter_sla_46_n34, 
      dp_ex_stage_alu_shifter_sla_46_n33, dp_ex_stage_alu_shifter_sla_46_n32, 
      dp_ex_stage_alu_shifter_sla_46_n31, dp_ex_stage_alu_shifter_sla_46_n30, 
      dp_ex_stage_alu_shifter_sla_46_n29, dp_ex_stage_alu_shifter_sla_46_n28, 
      dp_ex_stage_alu_shifter_sla_46_n27, dp_ex_stage_alu_shifter_sla_46_n26, 
      dp_ex_stage_alu_shifter_sla_46_n25, dp_ex_stage_alu_shifter_sla_46_n24, 
      dp_ex_stage_alu_shifter_sla_46_n23, dp_ex_stage_alu_shifter_sla_46_n22, 
      dp_ex_stage_alu_shifter_sla_46_n21, dp_ex_stage_alu_shifter_sla_46_n20, 
      dp_ex_stage_alu_shifter_sla_46_n19, dp_ex_stage_alu_shifter_sla_46_n18, 
      dp_ex_stage_alu_shifter_sla_46_n17, dp_ex_stage_alu_shifter_sla_46_n16, 
      dp_ex_stage_alu_shifter_sla_46_n15, dp_ex_stage_alu_shifter_sla_46_n14, 
      dp_ex_stage_alu_shifter_sla_46_n13, dp_ex_stage_alu_shifter_sla_46_n12, 
      dp_ex_stage_alu_shifter_sla_46_n11, dp_ex_stage_alu_shifter_sla_46_n10, 
      dp_ex_stage_alu_shifter_sla_46_n9, dp_ex_stage_alu_shifter_sla_46_n8, 
      dp_ex_stage_alu_shifter_sla_46_n7, dp_ex_stage_alu_shifter_sla_46_n6, 
      dp_ex_stage_alu_shifter_sla_46_n5, dp_ex_stage_alu_shifter_sla_46_n4, 
      dp_ex_stage_alu_shifter_sla_46_n3, dp_ex_stage_alu_shifter_sla_46_n2, 
      dp_ex_stage_alu_shifter_sla_46_n1, dp_ex_stage_alu_shifter_srl_41_n189, 
      dp_ex_stage_alu_shifter_srl_41_n188, dp_ex_stage_alu_shifter_srl_41_n187,
      dp_ex_stage_alu_shifter_srl_41_n186, dp_ex_stage_alu_shifter_srl_41_n185,
      dp_ex_stage_alu_shifter_srl_41_n184, dp_ex_stage_alu_shifter_srl_41_n183,
      dp_ex_stage_alu_shifter_srl_41_n182, dp_ex_stage_alu_shifter_srl_41_n181,
      dp_ex_stage_alu_shifter_srl_41_n180, dp_ex_stage_alu_shifter_srl_41_n179,
      dp_ex_stage_alu_shifter_srl_41_n178, dp_ex_stage_alu_shifter_srl_41_n177,
      dp_ex_stage_alu_shifter_srl_41_n176, dp_ex_stage_alu_shifter_srl_41_n175,
      dp_ex_stage_alu_shifter_srl_41_n174, dp_ex_stage_alu_shifter_srl_41_n173,
      dp_ex_stage_alu_shifter_srl_41_n172, dp_ex_stage_alu_shifter_srl_41_n171,
      dp_ex_stage_alu_shifter_srl_41_n170, dp_ex_stage_alu_shifter_srl_41_n169,
      dp_ex_stage_alu_shifter_srl_41_n168, dp_ex_stage_alu_shifter_srl_41_n167,
      dp_ex_stage_alu_shifter_srl_41_n166, dp_ex_stage_alu_shifter_srl_41_n165,
      dp_ex_stage_alu_shifter_srl_41_n164, dp_ex_stage_alu_shifter_srl_41_n163,
      dp_ex_stage_alu_shifter_srl_41_n162, dp_ex_stage_alu_shifter_srl_41_n161,
      dp_ex_stage_alu_shifter_srl_41_n160, dp_ex_stage_alu_shifter_srl_41_n159,
      dp_ex_stage_alu_shifter_srl_41_n158, dp_ex_stage_alu_shifter_srl_41_n157,
      dp_ex_stage_alu_shifter_srl_41_n156, dp_ex_stage_alu_shifter_srl_41_n155,
      dp_ex_stage_alu_shifter_srl_41_n154, dp_ex_stage_alu_shifter_srl_41_n153,
      dp_ex_stage_alu_shifter_srl_41_n152, dp_ex_stage_alu_shifter_srl_41_n151,
      dp_ex_stage_alu_shifter_srl_41_n150, dp_ex_stage_alu_shifter_srl_41_n149,
      dp_ex_stage_alu_shifter_srl_41_n148, dp_ex_stage_alu_shifter_srl_41_n147,
      dp_ex_stage_alu_shifter_srl_41_n146, dp_ex_stage_alu_shifter_srl_41_n145,
      dp_ex_stage_alu_shifter_srl_41_n144, dp_ex_stage_alu_shifter_srl_41_n143,
      dp_ex_stage_alu_shifter_srl_41_n142, dp_ex_stage_alu_shifter_srl_41_n141,
      dp_ex_stage_alu_shifter_srl_41_n140, dp_ex_stage_alu_shifter_srl_41_n139,
      dp_ex_stage_alu_shifter_srl_41_n138, dp_ex_stage_alu_shifter_srl_41_n137,
      dp_ex_stage_alu_shifter_srl_41_n136, dp_ex_stage_alu_shifter_srl_41_n135,
      dp_ex_stage_alu_shifter_srl_41_n134, dp_ex_stage_alu_shifter_srl_41_n133,
      dp_ex_stage_alu_shifter_srl_41_n132, dp_ex_stage_alu_shifter_srl_41_n131,
      dp_ex_stage_alu_shifter_srl_41_n130, dp_ex_stage_alu_shifter_srl_41_n129,
      dp_ex_stage_alu_shifter_srl_41_n128, dp_ex_stage_alu_shifter_srl_41_n127,
      dp_ex_stage_alu_shifter_srl_41_n126, dp_ex_stage_alu_shifter_srl_41_n125,
      dp_ex_stage_alu_shifter_srl_41_n124, dp_ex_stage_alu_shifter_srl_41_n123,
      dp_ex_stage_alu_shifter_srl_41_n122, dp_ex_stage_alu_shifter_srl_41_n121,
      dp_ex_stage_alu_shifter_srl_41_n120, dp_ex_stage_alu_shifter_srl_41_n119,
      dp_ex_stage_alu_shifter_srl_41_n118, dp_ex_stage_alu_shifter_srl_41_n117,
      dp_ex_stage_alu_shifter_srl_41_n116, dp_ex_stage_alu_shifter_srl_41_n115,
      dp_ex_stage_alu_shifter_srl_41_n114, dp_ex_stage_alu_shifter_srl_41_n113,
      dp_ex_stage_alu_shifter_srl_41_n112, dp_ex_stage_alu_shifter_srl_41_n111,
      dp_ex_stage_alu_shifter_srl_41_n110, dp_ex_stage_alu_shifter_srl_41_n109,
      dp_ex_stage_alu_shifter_srl_41_n108, dp_ex_stage_alu_shifter_srl_41_n107,
      dp_ex_stage_alu_shifter_srl_41_n106, dp_ex_stage_alu_shifter_srl_41_n105,
      dp_ex_stage_alu_shifter_srl_41_n104, dp_ex_stage_alu_shifter_srl_41_n103,
      dp_ex_stage_alu_shifter_srl_41_n102, dp_ex_stage_alu_shifter_srl_41_n101,
      dp_ex_stage_alu_shifter_srl_41_n100, dp_ex_stage_alu_shifter_srl_41_n99, 
      dp_ex_stage_alu_shifter_srl_41_n98, dp_ex_stage_alu_shifter_srl_41_n97, 
      dp_ex_stage_alu_shifter_srl_41_n96, dp_ex_stage_alu_shifter_srl_41_n95, 
      dp_ex_stage_alu_shifter_srl_41_n94, dp_ex_stage_alu_shifter_srl_41_n93, 
      dp_ex_stage_alu_shifter_srl_41_n92, dp_ex_stage_alu_shifter_srl_41_n91, 
      dp_ex_stage_alu_shifter_srl_41_n90, dp_ex_stage_alu_shifter_srl_41_n89, 
      dp_ex_stage_alu_shifter_srl_41_n88, dp_ex_stage_alu_shifter_srl_41_n87, 
      dp_ex_stage_alu_shifter_srl_41_n86, dp_ex_stage_alu_shifter_srl_41_n85, 
      dp_ex_stage_alu_shifter_srl_41_n84, dp_ex_stage_alu_shifter_srl_41_n83, 
      dp_ex_stage_alu_shifter_srl_41_n82, dp_ex_stage_alu_shifter_srl_41_n81, 
      dp_ex_stage_alu_shifter_srl_41_n80, dp_ex_stage_alu_shifter_srl_41_n79, 
      dp_ex_stage_alu_shifter_srl_41_n78, dp_ex_stage_alu_shifter_srl_41_n77, 
      dp_ex_stage_alu_shifter_srl_41_n76, dp_ex_stage_alu_shifter_srl_41_n75, 
      dp_ex_stage_alu_shifter_srl_41_n74, dp_ex_stage_alu_shifter_srl_41_n73, 
      dp_ex_stage_alu_shifter_srl_41_n72, dp_ex_stage_alu_shifter_srl_41_n71, 
      dp_ex_stage_alu_shifter_srl_41_n70, dp_ex_stage_alu_shifter_srl_41_n69, 
      dp_ex_stage_alu_shifter_srl_41_n68, dp_ex_stage_alu_shifter_srl_41_n67, 
      dp_ex_stage_alu_shifter_srl_41_n66, dp_ex_stage_alu_shifter_srl_41_n65, 
      dp_ex_stage_alu_shifter_srl_41_n64, dp_ex_stage_alu_shifter_srl_41_n63, 
      dp_ex_stage_alu_shifter_srl_41_n62, dp_ex_stage_alu_shifter_srl_41_n60, 
      dp_ex_stage_alu_shifter_srl_41_n59, dp_ex_stage_alu_shifter_srl_41_n58, 
      dp_ex_stage_alu_shifter_srl_41_n57, dp_ex_stage_alu_shifter_srl_41_n56, 
      dp_ex_stage_alu_shifter_srl_41_n55, dp_ex_stage_alu_shifter_srl_41_n54, 
      dp_ex_stage_alu_shifter_srl_41_n53, dp_ex_stage_alu_shifter_srl_41_n52, 
      dp_ex_stage_alu_shifter_srl_41_n51, dp_ex_stage_alu_shifter_srl_41_n50, 
      dp_ex_stage_alu_shifter_srl_41_n49, dp_ex_stage_alu_shifter_srl_41_n48, 
      dp_ex_stage_alu_shifter_srl_41_n47, dp_ex_stage_alu_shifter_srl_41_n46, 
      dp_ex_stage_alu_shifter_srl_41_n45, dp_ex_stage_alu_shifter_srl_41_n44, 
      dp_ex_stage_alu_shifter_srl_41_n43, dp_ex_stage_alu_shifter_srl_41_n42, 
      dp_ex_stage_alu_shifter_srl_41_n41, dp_ex_stage_alu_shifter_srl_41_n40, 
      dp_ex_stage_alu_shifter_srl_41_n39, dp_ex_stage_alu_shifter_srl_41_n38, 
      dp_ex_stage_alu_shifter_srl_41_n37, dp_ex_stage_alu_shifter_srl_41_n36, 
      dp_ex_stage_alu_shifter_srl_41_n35, dp_ex_stage_alu_shifter_srl_41_n34, 
      dp_ex_stage_alu_shifter_srl_41_n33, dp_ex_stage_alu_shifter_srl_41_n32, 
      dp_ex_stage_alu_shifter_srl_41_n31, dp_ex_stage_alu_shifter_srl_41_n30, 
      dp_ex_stage_alu_shifter_srl_41_n29, dp_ex_stage_alu_shifter_srl_41_n28, 
      dp_ex_stage_alu_shifter_srl_41_n27, dp_ex_stage_alu_shifter_srl_41_n26, 
      dp_ex_stage_alu_shifter_srl_41_n25, dp_ex_stage_alu_shifter_srl_41_n24, 
      dp_ex_stage_alu_shifter_srl_41_n23, dp_ex_stage_alu_shifter_srl_41_n22, 
      dp_ex_stage_alu_shifter_srl_41_n21, dp_ex_stage_alu_shifter_srl_41_n20, 
      dp_ex_stage_alu_shifter_srl_41_n19, dp_ex_stage_alu_shifter_srl_41_n18, 
      dp_ex_stage_alu_shifter_srl_41_n17, dp_ex_stage_alu_shifter_srl_41_n16, 
      dp_ex_stage_alu_shifter_srl_41_n15, dp_ex_stage_alu_shifter_srl_41_n14, 
      dp_ex_stage_alu_shifter_srl_41_n13, dp_ex_stage_alu_shifter_srl_41_n12, 
      dp_ex_stage_alu_shifter_srl_41_n11, dp_ex_stage_alu_shifter_srl_41_n10, 
      dp_ex_stage_alu_shifter_srl_41_n9, dp_ex_stage_alu_shifter_srl_41_n8, 
      dp_ex_stage_alu_shifter_srl_41_n7, dp_ex_stage_alu_shifter_srl_41_n6, 
      dp_ex_stage_alu_shifter_srl_41_n5, dp_ex_stage_alu_shifter_srl_41_n4, 
      dp_ex_stage_alu_shifter_srl_41_n3, dp_ex_stage_alu_shifter_srl_41_n2, 
      dp_ex_stage_alu_shifter_srl_41_n1, dp_ex_stage_alu_shifter_sra_39_n193, 
      dp_ex_stage_alu_shifter_sra_39_n192, dp_ex_stage_alu_shifter_sra_39_n191,
      dp_ex_stage_alu_shifter_sra_39_n190, dp_ex_stage_alu_shifter_sra_39_n189,
      dp_ex_stage_alu_shifter_sra_39_n188, dp_ex_stage_alu_shifter_sra_39_n187,
      dp_ex_stage_alu_shifter_sra_39_n186, dp_ex_stage_alu_shifter_sra_39_n185,
      dp_ex_stage_alu_shifter_sra_39_n184, dp_ex_stage_alu_shifter_sra_39_n183,
      dp_ex_stage_alu_shifter_sra_39_n182, dp_ex_stage_alu_shifter_sra_39_n181,
      dp_ex_stage_alu_shifter_sra_39_n180, dp_ex_stage_alu_shifter_sra_39_n179,
      dp_ex_stage_alu_shifter_sra_39_n178, dp_ex_stage_alu_shifter_sra_39_n177,
      dp_ex_stage_alu_shifter_sra_39_n176, dp_ex_stage_alu_shifter_sra_39_n175,
      dp_ex_stage_alu_shifter_sra_39_n174, dp_ex_stage_alu_shifter_sra_39_n173,
      dp_ex_stage_alu_shifter_sra_39_n172, dp_ex_stage_alu_shifter_sra_39_n171,
      dp_ex_stage_alu_shifter_sra_39_n170, dp_ex_stage_alu_shifter_sra_39_n169,
      dp_ex_stage_alu_shifter_sra_39_n168, dp_ex_stage_alu_shifter_sra_39_n167,
      dp_ex_stage_alu_shifter_sra_39_n166, dp_ex_stage_alu_shifter_sra_39_n165,
      dp_ex_stage_alu_shifter_sra_39_n164, dp_ex_stage_alu_shifter_sra_39_n163,
      dp_ex_stage_alu_shifter_sra_39_n162, dp_ex_stage_alu_shifter_sra_39_n161,
      dp_ex_stage_alu_shifter_sra_39_n160, dp_ex_stage_alu_shifter_sra_39_n159,
      dp_ex_stage_alu_shifter_sra_39_n158, dp_ex_stage_alu_shifter_sra_39_n157,
      dp_ex_stage_alu_shifter_sra_39_n156, dp_ex_stage_alu_shifter_sra_39_n155,
      dp_ex_stage_alu_shifter_sra_39_n154, dp_ex_stage_alu_shifter_sra_39_n153,
      dp_ex_stage_alu_shifter_sra_39_n152, dp_ex_stage_alu_shifter_sra_39_n151,
      dp_ex_stage_alu_shifter_sra_39_n150, dp_ex_stage_alu_shifter_sra_39_n149,
      dp_ex_stage_alu_shifter_sra_39_n148, dp_ex_stage_alu_shifter_sra_39_n147,
      dp_ex_stage_alu_shifter_sra_39_n146, dp_ex_stage_alu_shifter_sra_39_n145,
      dp_ex_stage_alu_shifter_sra_39_n144, dp_ex_stage_alu_shifter_sra_39_n143,
      dp_ex_stage_alu_shifter_sra_39_n142, dp_ex_stage_alu_shifter_sra_39_n141,
      dp_ex_stage_alu_shifter_sra_39_n140, dp_ex_stage_alu_shifter_sra_39_n139,
      dp_ex_stage_alu_shifter_sra_39_n138, dp_ex_stage_alu_shifter_sra_39_n137,
      dp_ex_stage_alu_shifter_sra_39_n136, dp_ex_stage_alu_shifter_sra_39_n135,
      dp_ex_stage_alu_shifter_sra_39_n134, dp_ex_stage_alu_shifter_sra_39_n133,
      dp_ex_stage_alu_shifter_sra_39_n132, dp_ex_stage_alu_shifter_sra_39_n131,
      dp_ex_stage_alu_shifter_sra_39_n130, dp_ex_stage_alu_shifter_sra_39_n129,
      dp_ex_stage_alu_shifter_sra_39_n128, dp_ex_stage_alu_shifter_sra_39_n127,
      dp_ex_stage_alu_shifter_sra_39_n126, dp_ex_stage_alu_shifter_sra_39_n125,
      dp_ex_stage_alu_shifter_sra_39_n124, dp_ex_stage_alu_shifter_sra_39_n123,
      dp_ex_stage_alu_shifter_sra_39_n122, dp_ex_stage_alu_shifter_sra_39_n121,
      dp_ex_stage_alu_shifter_sra_39_n120, dp_ex_stage_alu_shifter_sra_39_n119,
      dp_ex_stage_alu_shifter_sra_39_n118, dp_ex_stage_alu_shifter_sra_39_n117,
      dp_ex_stage_alu_shifter_sra_39_n116, dp_ex_stage_alu_shifter_sra_39_n115,
      dp_ex_stage_alu_shifter_sra_39_n114, dp_ex_stage_alu_shifter_sra_39_n113,
      dp_ex_stage_alu_shifter_sra_39_n112, dp_ex_stage_alu_shifter_sra_39_n111,
      dp_ex_stage_alu_shifter_sra_39_n110, dp_ex_stage_alu_shifter_sra_39_n109,
      dp_ex_stage_alu_shifter_sra_39_n108, dp_ex_stage_alu_shifter_sra_39_n107,
      dp_ex_stage_alu_shifter_sra_39_n106, dp_ex_stage_alu_shifter_sra_39_n105,
      dp_ex_stage_alu_shifter_sra_39_n104, dp_ex_stage_alu_shifter_sra_39_n103,
      dp_ex_stage_alu_shifter_sra_39_n102, dp_ex_stage_alu_shifter_sra_39_n101,
      dp_ex_stage_alu_shifter_sra_39_n100, dp_ex_stage_alu_shifter_sra_39_n99, 
      dp_ex_stage_alu_shifter_sra_39_n98, dp_ex_stage_alu_shifter_sra_39_n97, 
      dp_ex_stage_alu_shifter_sra_39_n96, dp_ex_stage_alu_shifter_sra_39_n95, 
      dp_ex_stage_alu_shifter_sra_39_n94, dp_ex_stage_alu_shifter_sra_39_n93, 
      dp_ex_stage_alu_shifter_sra_39_n92, dp_ex_stage_alu_shifter_sra_39_n91, 
      dp_ex_stage_alu_shifter_sra_39_n90, dp_ex_stage_alu_shifter_sra_39_n89, 
      dp_ex_stage_alu_shifter_sra_39_n88, dp_ex_stage_alu_shifter_sra_39_n87, 
      dp_ex_stage_alu_shifter_sra_39_n86, dp_ex_stage_alu_shifter_sra_39_n85, 
      dp_ex_stage_alu_shifter_sra_39_n84, dp_ex_stage_alu_shifter_sra_39_n83, 
      dp_ex_stage_alu_shifter_sra_39_n82, dp_ex_stage_alu_shifter_sra_39_n81, 
      dp_ex_stage_alu_shifter_sra_39_n80, dp_ex_stage_alu_shifter_sra_39_n79, 
      dp_ex_stage_alu_shifter_sra_39_n78, dp_ex_stage_alu_shifter_sra_39_n77, 
      dp_ex_stage_alu_shifter_sra_39_n76, dp_ex_stage_alu_shifter_sra_39_n75, 
      dp_ex_stage_alu_shifter_sra_39_n74, dp_ex_stage_alu_shifter_sra_39_n73, 
      dp_ex_stage_alu_shifter_sra_39_n72, dp_ex_stage_alu_shifter_sra_39_n71, 
      dp_ex_stage_alu_shifter_sra_39_n70, dp_ex_stage_alu_shifter_sra_39_n69, 
      dp_ex_stage_alu_shifter_sra_39_n68, dp_ex_stage_alu_shifter_sra_39_n67, 
      dp_ex_stage_alu_shifter_sra_39_n66, dp_ex_stage_alu_shifter_sra_39_n65, 
      dp_ex_stage_alu_shifter_sra_39_n64, dp_ex_stage_alu_shifter_sra_39_n63, 
      dp_ex_stage_alu_shifter_sra_39_n62, dp_ex_stage_alu_shifter_sra_39_n61, 
      dp_ex_stage_alu_shifter_sra_39_n60, dp_ex_stage_alu_shifter_sra_39_n59, 
      dp_ex_stage_alu_shifter_sra_39_n58, dp_ex_stage_alu_shifter_sra_39_n57, 
      dp_ex_stage_alu_shifter_sra_39_n56, dp_ex_stage_alu_shifter_sra_39_n55, 
      dp_ex_stage_alu_shifter_sra_39_n54, dp_ex_stage_alu_shifter_sra_39_n53, 
      dp_ex_stage_alu_shifter_sra_39_n52, dp_ex_stage_alu_shifter_sra_39_n51, 
      dp_ex_stage_alu_shifter_sra_39_n50, dp_ex_stage_alu_shifter_sra_39_n49, 
      dp_ex_stage_alu_shifter_sra_39_n48, dp_ex_stage_alu_shifter_sra_39_n47, 
      dp_ex_stage_alu_shifter_sra_39_n46, dp_ex_stage_alu_shifter_sra_39_n45, 
      dp_ex_stage_alu_shifter_sra_39_n43, dp_ex_stage_alu_shifter_sra_39_n42, 
      dp_ex_stage_alu_shifter_sra_39_n41, dp_ex_stage_alu_shifter_sra_39_n40, 
      dp_ex_stage_alu_shifter_sra_39_n39, dp_ex_stage_alu_shifter_sra_39_n38, 
      dp_ex_stage_alu_shifter_sra_39_n37, dp_ex_stage_alu_shifter_sra_39_n36, 
      dp_ex_stage_alu_shifter_sra_39_n35, dp_ex_stage_alu_shifter_sra_39_n34, 
      dp_ex_stage_alu_shifter_sra_39_n33, dp_ex_stage_alu_shifter_sra_39_n32, 
      dp_ex_stage_alu_shifter_sra_39_n31, dp_ex_stage_alu_shifter_sra_39_n30, 
      dp_ex_stage_alu_shifter_sra_39_n29, dp_ex_stage_alu_shifter_sra_39_n28, 
      dp_ex_stage_alu_shifter_sra_39_n27, dp_ex_stage_alu_shifter_sra_39_n26, 
      dp_ex_stage_alu_shifter_sra_39_n25, dp_ex_stage_alu_shifter_sra_39_n24, 
      dp_ex_stage_alu_shifter_sra_39_n23, dp_ex_stage_alu_shifter_sra_39_n22, 
      dp_ex_stage_alu_shifter_sra_39_n21, dp_ex_stage_alu_shifter_sra_39_n20, 
      dp_ex_stage_alu_shifter_sra_39_n19, dp_ex_stage_alu_shifter_sra_39_n18, 
      dp_ex_stage_alu_shifter_sra_39_n17, dp_ex_stage_alu_shifter_sra_39_n16, 
      dp_ex_stage_alu_shifter_sra_39_n15, dp_ex_stage_alu_shifter_sra_39_n14, 
      dp_ex_stage_alu_shifter_sra_39_n13, dp_ex_stage_alu_shifter_sra_39_n12, 
      dp_ex_stage_alu_shifter_sra_39_n11, dp_ex_stage_alu_shifter_sra_39_n10, 
      dp_ex_stage_alu_shifter_sra_39_n9, dp_ex_stage_alu_shifter_sra_39_n8, 
      dp_ex_stage_alu_shifter_sra_39_n7, dp_ex_stage_alu_shifter_sra_39_n6, 
      dp_ex_stage_alu_shifter_sra_39_n5, dp_ex_stage_alu_shifter_sra_39_n4, 
      dp_ex_stage_alu_shifter_sra_39_n3, dp_ex_stage_alu_shifter_sra_39_n2, 
      dp_ex_stage_alu_shifter_sra_39_n1, dp_ex_stage_alu_shifter_rol_32_n15, 
      dp_ex_stage_alu_shifter_rol_32_n14, dp_ex_stage_alu_shifter_rol_32_n13, 
      dp_ex_stage_alu_shifter_rol_32_n12, dp_ex_stage_alu_shifter_rol_32_n11, 
      dp_ex_stage_alu_shifter_rol_32_n10, dp_ex_stage_alu_shifter_rol_32_n9, 
      dp_ex_stage_alu_shifter_rol_32_n8, dp_ex_stage_alu_shifter_rol_32_n7, 
      dp_ex_stage_alu_shifter_rol_32_n6, dp_ex_stage_alu_shifter_rol_32_n5, 
      dp_ex_stage_alu_shifter_rol_32_n4, dp_ex_stage_alu_shifter_rol_32_n3, 
      dp_ex_stage_alu_shifter_rol_32_n2, dp_ex_stage_alu_shifter_rol_32_n1, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_0_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_1_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_2_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_3_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_4_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_5_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_6_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_7_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_8_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_9_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_10_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_11_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_12_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_13_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_14_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_15_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_16_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_17_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_18_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_19_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_20_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_21_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_22_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_23_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_24_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_25_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_26_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_27_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_28_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_29_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_30_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_4_31_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_0_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_1_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_2_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_3_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_4_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_5_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_6_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_7_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_8_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_9_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_10_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_11_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_12_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_13_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_14_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_15_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_16_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_17_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_18_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_19_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_20_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_21_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_22_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_23_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_24_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_25_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_26_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_27_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_28_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_29_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_30_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_3_31_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_0_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_1_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_2_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_3_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_4_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_5_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_6_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_7_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_8_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_9_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_10_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_11_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_12_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_13_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_14_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_15_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_16_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_17_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_18_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_19_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_20_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_21_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_22_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_23_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_24_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_25_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_26_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_27_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_28_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_29_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_30_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_2_31_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_0_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_1_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_2_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_3_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_4_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_5_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_6_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_7_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_8_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_9_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_10_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_11_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_12_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_13_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_14_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_15_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_16_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_17_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_18_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_19_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_20_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_21_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_22_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_23_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_24_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_25_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_26_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_27_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_28_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_29_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_30_port, 
      dp_ex_stage_alu_shifter_rol_32_ML_int_1_31_port, 
      dp_ex_stage_alu_shifter_ror_30_n15, dp_ex_stage_alu_shifter_ror_30_n14, 
      dp_ex_stage_alu_shifter_ror_30_n13, dp_ex_stage_alu_shifter_ror_30_n12, 
      dp_ex_stage_alu_shifter_ror_30_n11, dp_ex_stage_alu_shifter_ror_30_n10, 
      dp_ex_stage_alu_shifter_ror_30_n9, dp_ex_stage_alu_shifter_ror_30_n8, 
      dp_ex_stage_alu_shifter_ror_30_n7, dp_ex_stage_alu_shifter_ror_30_n6, 
      dp_ex_stage_alu_shifter_ror_30_n5, dp_ex_stage_alu_shifter_ror_30_n4, 
      dp_ex_stage_alu_shifter_ror_30_n3, dp_ex_stage_alu_shifter_ror_30_n2, 
      dp_ex_stage_alu_shifter_ror_30_n1, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_0_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_1_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_2_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_3_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_4_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_5_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_6_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_7_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_8_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_9_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_10_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_11_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_12_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_13_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_14_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_15_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_16_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_17_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_18_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_19_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_20_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_21_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_22_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_23_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_24_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_25_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_26_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_27_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_28_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_29_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_30_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_4_31_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_0_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_1_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_2_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_3_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_4_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_5_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_6_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_7_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_8_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_9_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_10_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_11_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_12_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_13_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_14_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_15_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_16_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_17_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_18_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_19_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_20_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_21_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_22_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_23_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_24_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_25_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_26_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_27_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_28_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_29_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_30_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_3_31_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_0_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_1_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_2_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_3_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_4_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_5_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_6_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_7_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_8_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_9_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_10_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_11_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_12_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_13_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_14_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_15_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_16_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_17_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_18_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_19_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_20_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_21_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_22_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_23_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_24_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_25_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_26_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_27_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_28_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_29_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_30_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_2_31_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_0_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_1_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_2_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_3_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_4_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_5_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_6_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_7_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_8_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_9_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_10_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_11_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_12_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_13_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_14_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_15_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_16_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_17_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_18_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_19_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_20_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_21_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_22_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_23_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_24_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_25_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_26_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_27_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_28_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_29_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_30_port, 
      dp_ex_stage_alu_shifter_ror_30_MR_int_1_31_port, dp_ex_stage_alu_r61_n222
      , dp_ex_stage_alu_r61_n221, dp_ex_stage_alu_r61_n220, 
      dp_ex_stage_alu_r61_n219, dp_ex_stage_alu_r61_n218, 
      dp_ex_stage_alu_r61_n217, dp_ex_stage_alu_r61_n216, 
      dp_ex_stage_alu_r61_n215, dp_ex_stage_alu_r61_n214, 
      dp_ex_stage_alu_r61_n213, dp_ex_stage_alu_r61_n212, 
      dp_ex_stage_alu_r61_n211, dp_ex_stage_alu_r61_n210, 
      dp_ex_stage_alu_r61_n209, dp_ex_stage_alu_r61_n208, 
      dp_ex_stage_alu_r61_n207, dp_ex_stage_alu_r61_n206, 
      dp_ex_stage_alu_r61_n205, dp_ex_stage_alu_r61_n204, 
      dp_ex_stage_alu_r61_n203, dp_ex_stage_alu_r61_n202, 
      dp_ex_stage_alu_r61_n201, dp_ex_stage_alu_r61_n200, 
      dp_ex_stage_alu_r61_n199, dp_ex_stage_alu_r61_n198, 
      dp_ex_stage_alu_r61_n197, dp_ex_stage_alu_r61_n196, 
      dp_ex_stage_alu_r61_n195, dp_ex_stage_alu_r61_n194, 
      dp_ex_stage_alu_r61_n193, dp_ex_stage_alu_r61_n192, 
      dp_ex_stage_alu_r61_n191, dp_ex_stage_alu_r61_n190, 
      dp_ex_stage_alu_r61_n189, dp_ex_stage_alu_r61_n188, 
      dp_ex_stage_alu_r61_n187, dp_ex_stage_alu_r61_n186, 
      dp_ex_stage_alu_r61_n185, dp_ex_stage_alu_r61_n184, 
      dp_ex_stage_alu_r61_n183, dp_ex_stage_alu_r61_n182, 
      dp_ex_stage_alu_r61_n181, dp_ex_stage_alu_r61_n180, 
      dp_ex_stage_alu_r61_n179, dp_ex_stage_alu_r61_n178, 
      dp_ex_stage_alu_r61_n177, dp_ex_stage_alu_r61_n176, 
      dp_ex_stage_alu_r61_n175, dp_ex_stage_alu_r61_n174, 
      dp_ex_stage_alu_r61_n173, dp_ex_stage_alu_r61_n172, 
      dp_ex_stage_alu_r61_n171, dp_ex_stage_alu_r61_n170, 
      dp_ex_stage_alu_r61_n169, dp_ex_stage_alu_r61_n168, 
      dp_ex_stage_alu_r61_n167, dp_ex_stage_alu_r61_n166, 
      dp_ex_stage_alu_r61_n165, dp_ex_stage_alu_r61_n164, 
      dp_ex_stage_alu_r61_n163, dp_ex_stage_alu_r61_n162, 
      dp_ex_stage_alu_r61_n161, dp_ex_stage_alu_r61_n160, 
      dp_ex_stage_alu_r61_n159, dp_ex_stage_alu_r61_n158, 
      dp_ex_stage_alu_r61_n157, dp_ex_stage_alu_r61_n156, 
      dp_ex_stage_alu_r61_n155, dp_ex_stage_alu_r61_n154, 
      dp_ex_stage_alu_r61_n153, dp_ex_stage_alu_r61_n152, 
      dp_ex_stage_alu_r61_n151, dp_ex_stage_alu_r61_n150, 
      dp_ex_stage_alu_r61_n149, dp_ex_stage_alu_r61_n148, 
      dp_ex_stage_alu_r61_n147, dp_ex_stage_alu_r61_n146, 
      dp_ex_stage_alu_r61_n145, dp_ex_stage_alu_r61_n144, 
      dp_ex_stage_alu_r61_n143, dp_ex_stage_alu_r61_n142, 
      dp_ex_stage_alu_r61_n141, dp_ex_stage_alu_r61_n140, 
      dp_ex_stage_alu_r61_n139, dp_ex_stage_alu_r61_n138, 
      dp_ex_stage_alu_r61_n137, dp_ex_stage_alu_r61_n136, 
      dp_ex_stage_alu_r61_n135, dp_ex_stage_alu_r61_n134, 
      dp_ex_stage_alu_r61_n133, dp_ex_stage_alu_r61_n132, 
      dp_ex_stage_alu_r61_n131, dp_ex_stage_alu_r61_n130, 
      dp_ex_stage_alu_r61_n129, dp_ex_stage_alu_r61_n128, 
      dp_ex_stage_alu_r61_n127, dp_ex_stage_alu_r61_n126, 
      dp_ex_stage_alu_r61_n125, dp_ex_stage_alu_r61_n124, 
      dp_ex_stage_alu_r61_n123, dp_ex_stage_alu_r61_n122, 
      dp_ex_stage_alu_r61_n121, dp_ex_stage_alu_r61_n120, 
      dp_ex_stage_alu_r61_n119, dp_ex_stage_alu_r61_n118, 
      dp_ex_stage_alu_r61_n117, dp_ex_stage_alu_r61_n116, 
      dp_ex_stage_alu_r61_n115, dp_ex_stage_alu_r61_n114, 
      dp_ex_stage_alu_r61_n113, dp_ex_stage_alu_r61_n112, 
      dp_ex_stage_alu_r61_n111, dp_ex_stage_alu_r61_n110, 
      dp_ex_stage_alu_r61_n109, dp_ex_stage_alu_r61_n108, 
      dp_ex_stage_alu_r61_n107, dp_ex_stage_alu_r61_n106, 
      dp_ex_stage_alu_r61_n105, dp_ex_stage_alu_r61_n104, 
      dp_ex_stage_alu_r61_n103, dp_ex_stage_alu_r61_n102, 
      dp_ex_stage_alu_r61_n101, dp_ex_stage_alu_r61_n100, 
      dp_ex_stage_alu_r61_n99, dp_ex_stage_alu_r61_n98, dp_ex_stage_alu_r61_n97
      , dp_ex_stage_alu_r61_n96, dp_ex_stage_alu_r61_n95, 
      dp_ex_stage_alu_r61_n94, dp_ex_stage_alu_r61_n93, dp_ex_stage_alu_r61_n92
      , dp_ex_stage_alu_r61_n91, dp_ex_stage_alu_r61_n90, 
      dp_ex_stage_alu_r61_n89, dp_ex_stage_alu_r61_n88, dp_ex_stage_alu_r61_n87
      , dp_ex_stage_alu_r61_n86, dp_ex_stage_alu_r61_n85, 
      dp_ex_stage_alu_r61_n84, dp_ex_stage_alu_r61_n83, dp_ex_stage_alu_r61_n82
      , dp_ex_stage_alu_r61_n81, dp_ex_stage_alu_r61_n80, 
      dp_ex_stage_alu_r61_n79, dp_ex_stage_alu_r61_n78, dp_ex_stage_alu_r61_n77
      , dp_ex_stage_alu_r61_n76, dp_ex_stage_alu_r61_n75, 
      dp_ex_stage_alu_r61_n74, dp_ex_stage_alu_r61_n73, dp_ex_stage_alu_r61_n72
      , dp_ex_stage_alu_r61_n71, dp_ex_stage_alu_r61_n70, 
      dp_ex_stage_alu_r61_n69, dp_ex_stage_alu_r61_n68, dp_ex_stage_alu_r61_n67
      , dp_ex_stage_alu_r61_n66, dp_ex_stage_alu_r61_n65, 
      dp_ex_stage_alu_r61_n64, dp_ex_stage_alu_r61_n63, dp_ex_stage_alu_r61_n62
      , dp_ex_stage_alu_r61_n61, dp_ex_stage_alu_r61_n60, 
      dp_ex_stage_alu_r61_n59, dp_ex_stage_alu_r61_n58, dp_ex_stage_alu_r61_n57
      , dp_ex_stage_alu_r61_n56, dp_ex_stage_alu_r61_n55, 
      dp_ex_stage_alu_r61_n54, dp_ex_stage_alu_r61_n53, dp_ex_stage_alu_r61_n52
      , dp_ex_stage_alu_r61_n51, dp_ex_stage_alu_r61_n50, 
      dp_ex_stage_alu_r61_n49, dp_ex_stage_alu_r61_n48, dp_ex_stage_alu_r61_n47
      , dp_ex_stage_alu_r61_n46, dp_ex_stage_alu_r61_n45, 
      dp_ex_stage_alu_r61_n44, dp_ex_stage_alu_r61_n43, dp_ex_stage_alu_r61_n42
      , dp_ex_stage_alu_r61_n41, dp_ex_stage_alu_r61_n40, 
      dp_ex_stage_alu_r61_n39, dp_ex_stage_alu_r61_n38, dp_ex_stage_alu_r61_n37
      , dp_ex_stage_alu_r61_n36, dp_ex_stage_alu_r61_n35, 
      dp_ex_stage_alu_r61_n34, dp_ex_stage_alu_r61_n33, dp_ex_stage_alu_r61_n32
      , dp_ex_stage_alu_r61_n31, dp_ex_stage_alu_r61_n30, 
      dp_ex_stage_alu_r61_n29, dp_ex_stage_alu_r61_n28, dp_ex_stage_alu_r61_n27
      , dp_ex_stage_alu_r61_n26, dp_ex_stage_alu_r61_n25, 
      dp_ex_stage_alu_r61_n24, dp_ex_stage_alu_r61_n23, dp_ex_stage_alu_r61_n22
      , dp_ex_stage_alu_r61_n21, dp_ex_stage_alu_r61_n20, 
      dp_ex_stage_alu_r61_n19, dp_ex_stage_alu_r61_n18, dp_ex_stage_alu_r61_n17
      , dp_ex_stage_alu_r61_n16, dp_ex_stage_alu_r61_n15, 
      dp_ex_stage_alu_r61_n14, dp_ex_stage_alu_r61_n13, dp_ex_stage_alu_r61_n12
      , dp_ex_stage_alu_r61_n11, dp_ex_stage_alu_r61_n10, 
      dp_ex_stage_alu_r61_n9, dp_ex_stage_alu_r61_n8, dp_ex_stage_alu_r61_n7, 
      dp_ex_stage_alu_r61_n6, dp_ex_stage_alu_r61_n5, dp_ex_stage_alu_r61_n4, 
      dp_ex_stage_alu_r61_n3, dp_ex_stage_alu_r61_n2, dp_ex_stage_alu_r61_n1, 
      dp_ex_stage_alu_r60_n315, dp_ex_stage_alu_r60_n314, 
      dp_ex_stage_alu_r60_n313, dp_ex_stage_alu_r60_n312, 
      dp_ex_stage_alu_r60_n311, dp_ex_stage_alu_r60_n310, 
      dp_ex_stage_alu_r60_n309, dp_ex_stage_alu_r60_n308, 
      dp_ex_stage_alu_r60_n307, dp_ex_stage_alu_r60_n306, 
      dp_ex_stage_alu_r60_n305, dp_ex_stage_alu_r60_n304, 
      dp_ex_stage_alu_r60_n303, dp_ex_stage_alu_r60_n302, 
      dp_ex_stage_alu_r60_n301, dp_ex_stage_alu_r60_n300, 
      dp_ex_stage_alu_r60_n299, dp_ex_stage_alu_r60_n298, 
      dp_ex_stage_alu_r60_n297, dp_ex_stage_alu_r60_n296, 
      dp_ex_stage_alu_r60_n295, dp_ex_stage_alu_r60_n294, 
      dp_ex_stage_alu_r60_n293, dp_ex_stage_alu_r60_n292, 
      dp_ex_stage_alu_r60_n291, dp_ex_stage_alu_r60_n290, 
      dp_ex_stage_alu_r60_n289, dp_ex_stage_alu_r60_n288, 
      dp_ex_stage_alu_r60_n287, dp_ex_stage_alu_r60_n286, 
      dp_ex_stage_alu_r60_n285, dp_ex_stage_alu_r60_n284, 
      dp_ex_stage_alu_r60_n283, dp_ex_stage_alu_r60_n282, 
      dp_ex_stage_alu_r60_n281, dp_ex_stage_alu_r60_n280, 
      dp_ex_stage_alu_r60_n279, dp_ex_stage_alu_r60_n278, 
      dp_ex_stage_alu_r60_n277, dp_ex_stage_alu_r60_n276, 
      dp_ex_stage_alu_r60_n275, dp_ex_stage_alu_r60_n274, 
      dp_ex_stage_alu_r60_n273, dp_ex_stage_alu_r60_n272, 
      dp_ex_stage_alu_r60_n271, dp_ex_stage_alu_r60_n270, 
      dp_ex_stage_alu_r60_n269, dp_ex_stage_alu_r60_n268, 
      dp_ex_stage_alu_r60_n267, dp_ex_stage_alu_r60_n266, 
      dp_ex_stage_alu_r60_n265, dp_ex_stage_alu_r60_n264, 
      dp_ex_stage_alu_r60_n263, dp_ex_stage_alu_r60_n262, 
      dp_ex_stage_alu_r60_n261, dp_ex_stage_alu_r60_n260, 
      dp_ex_stage_alu_r60_n259, dp_ex_stage_alu_r60_n258, 
      dp_ex_stage_alu_r60_n257, dp_ex_stage_alu_r60_n256, 
      dp_ex_stage_alu_r60_n255, dp_ex_stage_alu_r60_n254, 
      dp_ex_stage_alu_r60_n253, dp_ex_stage_alu_r60_n252, 
      dp_ex_stage_alu_r60_n251, dp_ex_stage_alu_r60_n250, 
      dp_ex_stage_alu_r60_n249, dp_ex_stage_alu_r60_n248, 
      dp_ex_stage_alu_r60_n247, dp_ex_stage_alu_r60_n246, 
      dp_ex_stage_alu_r60_n245, dp_ex_stage_alu_r60_n244, 
      dp_ex_stage_alu_r60_n243, dp_ex_stage_alu_r60_n242, 
      dp_ex_stage_alu_r60_n241, dp_ex_stage_alu_r60_n240, 
      dp_ex_stage_alu_r60_n239, dp_ex_stage_alu_r60_n238, 
      dp_ex_stage_alu_r60_n237, dp_ex_stage_alu_r60_n236, 
      dp_ex_stage_alu_r60_n235, dp_ex_stage_alu_r60_n234, 
      dp_ex_stage_alu_r60_n233, dp_ex_stage_alu_r60_n232, 
      dp_ex_stage_alu_r60_n231, dp_ex_stage_alu_r60_n230, 
      dp_ex_stage_alu_r60_n229, dp_ex_stage_alu_r60_n228, 
      dp_ex_stage_alu_r60_n227, dp_ex_stage_alu_r60_n226, 
      dp_ex_stage_alu_r60_n225, dp_ex_stage_alu_r60_n224, 
      dp_ex_stage_alu_r60_n223, dp_ex_stage_alu_r60_n222, 
      dp_ex_stage_alu_r60_n221, dp_ex_stage_alu_r60_n220, 
      dp_ex_stage_alu_r60_n219, dp_ex_stage_alu_r60_n218, 
      dp_ex_stage_alu_r60_n217, dp_ex_stage_alu_r60_n216, 
      dp_ex_stage_alu_r60_n215, dp_ex_stage_alu_r60_n214, 
      dp_ex_stage_alu_r60_n213, dp_ex_stage_alu_r60_n212, 
      dp_ex_stage_alu_r60_n211, dp_ex_stage_alu_r60_n210, 
      dp_ex_stage_alu_r60_n209, dp_ex_stage_alu_r60_n208, 
      dp_ex_stage_alu_r60_n207, dp_ex_stage_alu_r60_n206, 
      dp_ex_stage_alu_r60_n205, dp_ex_stage_alu_r60_n204, 
      dp_ex_stage_alu_r60_n203, dp_ex_stage_alu_r60_n202, 
      dp_ex_stage_alu_r60_n201, dp_ex_stage_alu_r60_n200, 
      dp_ex_stage_alu_r60_n199, dp_ex_stage_alu_r60_n198, 
      dp_ex_stage_alu_r60_n197, dp_ex_stage_alu_r60_n196, 
      dp_ex_stage_alu_r60_n195, dp_ex_stage_alu_r60_n194, 
      dp_ex_stage_alu_r60_n193, dp_ex_stage_alu_r60_n192, 
      dp_ex_stage_alu_r60_n191, dp_ex_stage_alu_r60_n190, 
      dp_ex_stage_alu_r60_n189, dp_ex_stage_alu_r60_n188, 
      dp_ex_stage_alu_r60_n187, dp_ex_stage_alu_r60_n186, 
      dp_ex_stage_alu_r60_n185, dp_ex_stage_alu_r60_n184, 
      dp_ex_stage_alu_r60_n183, dp_ex_stage_alu_r60_n182, 
      dp_ex_stage_alu_r60_n181, dp_ex_stage_alu_r60_n180, 
      dp_ex_stage_alu_r60_n179, dp_ex_stage_alu_r60_n178, 
      dp_ex_stage_alu_r60_n177, dp_ex_stage_alu_r60_n176, 
      dp_ex_stage_alu_r60_n175, dp_ex_stage_alu_r60_n174, 
      dp_ex_stage_alu_r60_n173, dp_ex_stage_alu_r60_n172, 
      dp_ex_stage_alu_r60_n171, dp_ex_stage_alu_r60_n170, 
      dp_ex_stage_alu_r60_n169, dp_ex_stage_alu_r60_n168, 
      dp_ex_stage_alu_r60_n167, dp_ex_stage_alu_r60_n166, 
      dp_ex_stage_alu_r60_n165, dp_ex_stage_alu_r60_n164, 
      dp_ex_stage_alu_r60_n163, dp_ex_stage_alu_r60_n162, 
      dp_ex_stage_alu_r60_n161, dp_ex_stage_alu_r60_n160, 
      dp_ex_stage_alu_r60_n159, dp_ex_stage_alu_r60_n158, 
      dp_ex_stage_alu_r60_n157, dp_ex_stage_alu_r60_n156, 
      dp_ex_stage_alu_r60_n155, dp_ex_stage_alu_r60_n154, 
      dp_ex_stage_alu_r60_n153, dp_ex_stage_alu_r60_n152, 
      dp_ex_stage_alu_r60_n151, dp_ex_stage_alu_r60_n150, 
      dp_ex_stage_alu_r60_n149, dp_ex_stage_alu_r60_n148, 
      dp_ex_stage_alu_r60_n147, dp_ex_stage_alu_r60_n146, 
      dp_ex_stage_alu_r60_n145, dp_ex_stage_alu_r60_n144, 
      dp_ex_stage_alu_r60_n143, dp_ex_stage_alu_r60_n142, 
      dp_ex_stage_alu_r60_n141, dp_ex_stage_alu_r60_n140, 
      dp_ex_stage_alu_r60_n139, dp_ex_stage_alu_r60_n138, 
      dp_ex_stage_alu_r60_n137, dp_ex_stage_alu_r60_n136, 
      dp_ex_stage_alu_r60_n135, dp_ex_stage_alu_r60_n134, 
      dp_ex_stage_alu_r60_n133, dp_ex_stage_alu_r60_n132, 
      dp_ex_stage_alu_r60_n131, dp_ex_stage_alu_r60_n130, 
      dp_ex_stage_alu_r60_n129, dp_ex_stage_alu_r60_n128, 
      dp_ex_stage_alu_r60_n127, dp_ex_stage_alu_r60_n126, 
      dp_ex_stage_alu_r60_n125, dp_ex_stage_alu_r60_n124, 
      dp_ex_stage_alu_r60_n123, dp_ex_stage_alu_r60_n122, 
      dp_ex_stage_alu_r60_n121, dp_ex_stage_alu_r60_n120, 
      dp_ex_stage_alu_r60_n119, dp_ex_stage_alu_r60_n118, 
      dp_ex_stage_alu_r60_n117, dp_ex_stage_alu_r60_n116, 
      dp_ex_stage_alu_r60_n115, dp_ex_stage_alu_r60_n114, 
      dp_ex_stage_alu_r60_n113, dp_ex_stage_alu_r60_n112, 
      dp_ex_stage_alu_r60_n111, dp_ex_stage_alu_r60_n110, 
      dp_ex_stage_alu_r60_n109, dp_ex_stage_alu_r60_n108, 
      dp_ex_stage_alu_r60_n107, dp_ex_stage_alu_r60_n106, 
      dp_ex_stage_alu_r60_n105, dp_ex_stage_alu_r60_n104, 
      dp_ex_stage_alu_r60_n103, dp_ex_stage_alu_r60_n102, 
      dp_ex_stage_alu_r60_n101, dp_ex_stage_alu_r60_n100, 
      dp_ex_stage_alu_r60_n99, dp_ex_stage_alu_r60_n98, dp_ex_stage_alu_r60_n97
      , dp_ex_stage_alu_r60_n96, dp_ex_stage_alu_r60_n95, 
      dp_ex_stage_alu_r60_n94, dp_ex_stage_alu_r60_n93, dp_ex_stage_alu_r60_n92
      , dp_ex_stage_alu_r60_n91, dp_ex_stage_alu_r60_n90, 
      dp_ex_stage_alu_r60_n89, dp_ex_stage_alu_r60_n88, dp_ex_stage_alu_r60_n87
      , dp_ex_stage_alu_r60_n86, dp_ex_stage_alu_r60_n85, 
      dp_ex_stage_alu_r60_n84, dp_ex_stage_alu_r60_n83, dp_ex_stage_alu_r60_n82
      , dp_ex_stage_alu_r60_n81, dp_ex_stage_alu_r60_n80, 
      dp_ex_stage_alu_r60_n79, dp_ex_stage_alu_r60_n78, dp_ex_stage_alu_r60_n77
      , dp_ex_stage_alu_r60_n76, dp_ex_stage_alu_r60_n75, 
      dp_ex_stage_alu_r60_n74, dp_ex_stage_alu_r60_n73, dp_ex_stage_alu_r60_n72
      , dp_ex_stage_alu_r60_n71, dp_ex_stage_alu_r60_n70, 
      dp_ex_stage_alu_r60_n69, dp_ex_stage_alu_r60_n68, dp_ex_stage_alu_r60_n67
      , dp_ex_stage_alu_r60_n66, dp_ex_stage_alu_r60_n65, 
      dp_ex_stage_alu_r60_n64, dp_ex_stage_alu_r60_n63, dp_ex_stage_alu_r60_n62
      , dp_ex_stage_alu_r60_n61, dp_ex_stage_alu_r60_n60, 
      dp_ex_stage_alu_r60_n59, dp_ex_stage_alu_r60_n58, dp_ex_stage_alu_r60_n57
      , dp_ex_stage_alu_r60_n56, dp_ex_stage_alu_r60_n55, 
      dp_ex_stage_alu_r60_n54, dp_ex_stage_alu_r60_n53, dp_ex_stage_alu_r60_n52
      , dp_ex_stage_alu_r60_n51, dp_ex_stage_alu_r60_n50, 
      dp_ex_stage_alu_r60_n49, dp_ex_stage_alu_r60_n48, dp_ex_stage_alu_r60_n47
      , dp_ex_stage_alu_r60_n46, dp_ex_stage_alu_r60_n45, 
      dp_ex_stage_alu_r60_n44, dp_ex_stage_alu_r60_n43, dp_ex_stage_alu_r60_n42
      , dp_ex_stage_alu_r60_n41, dp_ex_stage_alu_r60_n40, 
      dp_ex_stage_alu_r60_n39, dp_ex_stage_alu_r60_n38, dp_ex_stage_alu_r60_n37
      , dp_ex_stage_alu_r60_n36, dp_ex_stage_alu_r60_n35, 
      dp_ex_stage_alu_r60_n34, dp_ex_stage_alu_r60_n33, dp_ex_stage_alu_r60_n32
      , dp_ex_stage_alu_r60_n31, dp_ex_stage_alu_r60_n30, 
      dp_ex_stage_alu_r60_n29, dp_ex_stage_alu_r60_n28, dp_ex_stage_alu_r60_n27
      , dp_ex_stage_alu_r60_n26, dp_ex_stage_alu_r60_n25, 
      dp_ex_stage_alu_r60_n24, dp_ex_stage_alu_r60_n23, dp_ex_stage_alu_r60_n22
      , dp_ex_stage_alu_r60_n21, dp_ex_stage_alu_r60_n20, 
      dp_ex_stage_alu_r60_n19, dp_ex_stage_alu_r60_n17, dp_ex_stage_alu_r60_n16
      , dp_ex_stage_alu_r60_n15, dp_ex_stage_alu_r60_n14, 
      dp_ex_stage_alu_r60_n13, dp_ex_stage_alu_r60_n12, dp_ex_stage_alu_r60_n11
      , dp_ex_stage_alu_r60_n10, dp_ex_stage_alu_r60_n9, dp_ex_stage_alu_r60_n8
      , dp_ex_stage_alu_r60_n7, dp_ex_stage_alu_r60_n6, dp_ex_stage_alu_r60_n5,
      dp_ex_stage_alu_r60_n4, dp_ex_stage_alu_r60_n3, dp_ex_stage_alu_r60_n2, 
      dp_ex_stage_alu_r60_n1, n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, 
      n_1006, n_1007, n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, 
      n_1015, n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023, 
      n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, 
      n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, n_1055, n_1056, n_1057, n_1058, n_1059, 
      n_1060, n_1061, n_1062, n_1063, n_1064, n_1065, n_1066, n_1067, n_1068, 
      n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, 
      n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, 
      n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, 
      n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, 
      n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, 
      n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, 
      n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, 
      n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, 
      n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, 
      n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, 
      n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, 
      n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, 
      n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, 
      n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, 
      n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, 
      n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, 
      n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, 
      n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, 
      n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, 
      n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, 
      n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, 
      n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, 
      n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, 
      n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, 
      n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, 
      n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, 
      n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, 
      n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, 
      n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, 
      n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, 
      n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, 
      n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, 
      n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, 
      n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, 
      n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, 
      n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, 
      n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, 
      n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, 
      n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, 
      n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, 
      n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, 
      n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, 
      n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, 
      n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, 
      n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, 
      n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, 
      n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, 
      n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, 
      n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, 
      n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, 
      n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, 
      n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, 
      n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, 
      n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, 
      n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, 
      n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, 
      n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, 
      n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, 
      n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, 
      n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, 
      n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, 
      n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, 
      n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, 
      n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, 
      n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, 
      n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, 
      n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, 
      n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, 
      n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, 
      n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, 
      n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, 
      n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, 
      n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, 
      n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, 
      n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, 
      n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, 
      n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, 
      n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, 
      n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, 
      n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, 
      n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, 
      n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, 
      n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, 
      n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, 
      n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, 
      n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, 
      n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, 
      n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, 
      n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, 
      n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, 
      n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, 
      n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, 
      n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, 
      n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, 
      n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, 
      n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, 
      n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, 
      n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, 
      n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, 
      n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, 
      n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, 
      n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, 
      n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, 
      n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, 
      n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, 
      n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, 
      n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, 
      n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, 
      n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, 
      n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, 
      n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, 
      n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, 
      n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, 
      n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, 
      n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, 
      n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, 
      n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, 
      n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, 
      n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, 
      n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, 
      n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, 
      n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, 
      n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, 
      n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, 
      n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, 
      n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, 
      n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, 
      n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, 
      n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, 
      n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, 
      n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, 
      n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, 
      n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, 
      n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, 
      n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, 
      n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, 
      n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, 
      n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, 
      n_2311, n_2312 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, dp_if_stage_NPC_4_i_1_port, 
      dp_if_stage_NPC_4_i_0_port );
   IRAM_ISSUE <= IRAM_ISSUE_port;
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, DRAM_ADDRESS_0_port );
   DRAM_ISSUE <= DRAM_ISSUE_port;
   DRAM_READNOTWRITE <= DRAM_READNOTWRITE_port;
   
   rf_en_i <= '1';
   rf_ret_i <= '0';
   rf_call_i <= '0';
   CU_I_U264 : INV_X2 port map( A => IRAM_DATA(0), ZN => CU_I_n291);
   CU_I_U263 : NAND2_X1 port map( A1 => alu_op_i_1_port, A2 => CU_I_n63, ZN => 
                           CU_I_n79);
   CU_I_U262 : NAND2_X1 port map( A1 => alu_op_i_3_port, A2 => CU_I_n63, ZN => 
                           CU_I_n82);
   CU_I_U261 : NAND2_X1 port map( A1 => CU_I_n293, A2 => CU_I_n66, ZN => 
                           CU_I_n167);
   CU_I_U260 : NAND2_X1 port map( A1 => alu_op_i_2_port, A2 => CU_I_n63, ZN => 
                           CU_I_n81);
   CU_I_U259 : OAI211_X1 port map( C1 => CU_I_n69, C2 => CU_I_n35, A => 
                           CU_I_n80, B => CU_I_n81, ZN => CU_I_n213);
   CU_I_U258 : NAND2_X1 port map( A1 => CU_I_n180, A2 => CU_I_n132, ZN => 
                           CU_I_n102);
   CU_I_U257 : AND2_X1 port map( A1 => CU_I_n102, A2 => CU_I_n127, ZN => 
                           CU_I_n206);
   CU_I_U256 : AOI21_X1 port map( B1 => CU_I_n117, B2 => CU_I_n180, A => 
                           CU_I_n75, ZN => CU_I_n145);
   CU_I_U255 : INV_X1 port map( A => CU_I_n47, ZN => CU_I_n261);
   CU_I_U254 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n8, B1 => 
                           CU_I_n175, B2 => CU_I_n67, ZN => CU_I_n241);
   CU_I_U253 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n36, A => CU_I_n79
                           , ZN => CU_I_n212);
   CU_I_U252 : NOR3_X1 port map( A1 => CU_I_n157, A2 => IRAM_DATA(30), A3 => 
                           CU_I_n276, ZN => CU_I_n152);
   CU_I_U251 : AND2_X1 port map( A1 => CU_I_n202, A2 => CU_I_n276, ZN => 
                           CU_I_n176);
   CU_I_U250 : NOR3_X1 port map( A1 => CU_I_n276, A2 => CU_I_n157, A3 => 
                           CU_I_n274, ZN => CU_I_n207);
   CU_I_U249 : NOR4_X1 port map( A1 => IRAM_DATA(30), A2 => IRAM_DATA(29), A3 
                           => CU_I_n276, A4 => CU_I_n279, ZN => CU_I_n150);
   CU_I_U248 : AOI21_X1 port map( B1 => CU_I_n278, B2 => CU_I_n276, A => 
                           IRAM_DATA(30), ZN => CU_I_n162);
   CU_I_U247 : NAND4_X1 port map( A1 => CU_I_n161, A2 => CU_I_n154, A3 => 
                           IRAM_DATA(29), A4 => CU_I_n276, ZN => CU_I_n187);
   CU_I_U246 : AOI22_X1 port map( A1 => CU_I_n259, A2 => CU_I_n276, B1 => 
                           IRAM_DATA(30), B2 => CU_I_n156, ZN => CU_I_n147);
   CU_I_U245 : NOR3_X1 port map( A1 => IRAM_DATA(28), A2 => IRAM_DATA(30), A3 
                           => CU_I_n157, ZN => CU_I_n133);
   CU_I_U244 : NAND2_X1 port map( A1 => CU_I_n154, A2 => CU_I_n133, ZN => 
                           CU_I_n101);
   CU_I_U243 : NAND2_X1 port map( A1 => CU_I_n38, A2 => CU_I_n117, ZN => 
                           CU_I_n155);
   CU_I_U242 : AOI21_X1 port map( B1 => CU_I_n132, B2 => CU_I_n38, A => 
                           CU_I_n264, ZN => CU_I_n131);
   CU_I_U241 : NOR2_X1 port map( A1 => CU_I_n267, A2 => CU_I_n194, ZN => 
                           CU_I_n192);
   CU_I_U240 : OAI211_X1 port map( C1 => CU_I_n48, C2 => CU_I_n281, A => 
                           CU_I_n130, B => CU_I_n206, ZN => CU_I_n111);
   CU_I_U239 : AOI211_X1 port map( C1 => CU_I_n152, C2 => CU_I_n160, A => 
                           CU_I_n111, B => CU_I_n204, ZN => CU_I_n87);
   CU_I_U238 : NOR3_X1 port map( A1 => CU_I_n110, A2 => CU_I_n41, A3 => 
                           CU_I_n112, ZN => CU_I_n109);
   CU_I_U237 : NAND2_X1 port map( A1 => CU_I_n292, A2 => CU_I_n64, ZN => 
                           CU_I_n166);
   CU_I_U236 : OAI211_X1 port map( C1 => CU_I_n69, C2 => CU_I_n33, A => 
                           CU_I_n80, B => CU_I_n83, ZN => CU_I_n215);
   CU_I_U235 : AOI22_X1 port map( A1 => CU_I_n68, A2 => CU_I_cw1_1_port, B1 => 
                           CU_I_n171, B2 => CU_I_n172, ZN => CU_I_n170);
   CU_I_U234 : INV_X1 port map( A => CU_I_n170, ZN => CU_I_n74);
   CU_I_U233 : AOI22_X1 port map( A1 => CU_I_n291, A2 => IRAM_DATA(2), B1 => 
                           CU_I_n289, B2 => CU_I_n94, ZN => CU_I_n93);
   CU_I_U232 : OR2_X1 port map( A1 => CU_I_n93, A2 => IRAM_DATA(3), ZN => 
                           CU_I_n88);
   CU_I_U223 : NAND2_X1 port map( A1 => pipe_clear_n_i, A2 => CU_I_n30, ZN => 
                           jump_en_i);
   CU_I_U215 : INV_X1 port map( A => IRAM_DATA(26), ZN => CU_I_n282);
   CU_I_U214 : INV_X1 port map( A => IRAM_DATA(4), ZN => CU_I_n286);
   CU_I_U213 : NAND2_X1 port map( A1 => IRAM_READY, A2 => IRAM_ISSUE_port, ZN 
                           => CU_I_n78);
   CU_I_U212 : INV_X1 port map( A => IRAM_DATA(27), ZN => CU_I_n279);
   CU_I_U211 : INV_X1 port map( A => IRAM_DATA(31), ZN => CU_I_n266);
   CU_I_U210 : INV_X1 port map( A => CU_I_n126, ZN => CU_I_n285);
   CU_I_U209 : INV_X1 port map( A => CU_I_n185, ZN => CU_I_n260);
   CU_I_U208 : NAND2_X1 port map( A1 => regrd_sel_i, A2 => CU_I_n65, ZN => 
                           CU_I_n190);
   CU_I_U207 : OAI21_X1 port map( B1 => CU_I_n260, B2 => CU_I_n49, A => 
                           CU_I_n190, ZN => CU_I_n247);
   CU_I_U206 : AND3_X1 port map( A1 => CU_I_n114, A2 => CU_I_n196, A3 => 
                           CU_I_n187, ZN => CU_I_n197);
   CU_I_U205 : NAND2_X1 port map( A1 => rf_rs2_en_i, A2 => CU_I_n66, ZN => 
                           CU_I_n198);
   CU_I_U204 : OAI21_X1 port map( B1 => CU_I_n197, B2 => CU_I_n49, A => 
                           CU_I_n198, ZN => CU_I_n251);
   CU_I_U203 : NAND2_X1 port map( A1 => imm_isoff_i, A2 => CU_I_n66, ZN => 
                           CU_I_n195);
   CU_I_U202 : OAI21_X1 port map( B1 => CU_I_n268, B2 => CU_I_n49, A => 
                           CU_I_n195, ZN => CU_I_n250);
   CU_I_U201 : NAND2_X1 port map( A1 => imm_uns_i, A2 => CU_I_n66, ZN => 
                           CU_I_n193);
   CU_I_U200 : OAI21_X1 port map( B1 => CU_I_n192, B2 => CU_I_n49, A => 
                           CU_I_n193, ZN => CU_I_n249);
   CU_I_U199 : NOR4_X1 port map( A1 => CU_I_n267, A2 => CU_I_n179, A3 => 
                           CU_I_n184, A4 => CU_I_n181, ZN => CU_I_n199);
   CU_I_U198 : NAND2_X1 port map( A1 => rf_rs1_en_i, A2 => CU_I_n67, ZN => 
                           CU_I_n200);
   CU_I_U197 : OAI21_X1 port map( B1 => CU_I_n199, B2 => CU_I_n49, A => 
                           CU_I_n200, ZN => CU_I_n252);
   CU_I_U196 : OR3_X1 port map( A1 => CU_I_n157, A2 => IRAM_DATA(28), A3 => 
                           CU_I_n274, ZN => CU_I_n116);
   CU_I_U195 : OAI21_X1 port map( B1 => CU_I_n2, B2 => pipe_ex_mem_en_i, A => 
                           CU_I_n182, ZN => CU_I_n248);
   CU_I_U194 : NAND2_X1 port map( A1 => CU_I_n91, A2 => CU_I_n92, ZN => 
                           CU_I_n90);
   CU_I_U193 : OAI21_X1 port map( B1 => pipe_if_id_en_i, B2 => CU_I_n6, A => 
                           CU_I_n182, ZN => CU_I_n243);
   CU_I_U192 : NAND4_X1 port map( A1 => CU_I_n91, A2 => IRAM_DATA(1), A3 => 
                           IRAM_DATA(0), A4 => CU_I_n289, ZN => CU_I_n128);
   CU_I_U191 : NAND2_X1 port map( A1 => CU_I_n127, A2 => CU_I_n128, ZN => 
                           CU_I_n105);
   CU_I_U190 : INV_X1 port map( A => IRAM_DATA(5), ZN => CU_I_n284);
   CU_I_U189 : NOR2_X1 port map( A1 => IRAM_DATA(2), A2 => CU_I_n291, ZN => 
                           CU_I_n144);
   CU_I_U188 : NAND2_X1 port map( A1 => DRAM_READNOTWRITE_port, A2 => CU_I_n67,
                           ZN => CU_I_n209);
   CU_I_U187 : OAI211_X1 port map( C1 => CU_I_n69, C2 => CU_I_n16, A => 
                           CU_I_n80, B => CU_I_n209, ZN => CU_I_n253);
   CU_I_U186 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n3, A => CU_I_n166
                           , ZN => CU_I_n226);
   CU_I_U185 : NAND2_X1 port map( A1 => mem_in_en_i, A2 => CU_I_n65, ZN => 
                           CU_I_n168);
   CU_I_U184 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n5, A => CU_I_n168
                           , ZN => CU_I_n228);
   CU_I_U183 : NAND2_X1 port map( A1 => npc_wb_en_i, A2 => CU_I_n65, ZN => 
                           CU_I_n169);
   CU_I_U182 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n6, A => CU_I_n169
                           , ZN => CU_I_n229);
   CU_I_U181 : NAND2_X1 port map( A1 => wb_mux_sel_i, A2 => CU_I_n64, ZN => 
                           CU_I_n165);
   CU_I_U180 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n31, A => 
                           CU_I_n165, ZN => CU_I_n222);
   CU_I_U179 : NAND2_X1 port map( A1 => rf_we_i, A2 => CU_I_n64, ZN => 
                           CU_I_n164);
   CU_I_U178 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n32, A => 
                           CU_I_n164, ZN => CU_I_n221);
   CU_I_U177 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n34, A => CU_I_n82
                           , ZN => CU_I_n214);
   CU_I_U176 : NAND2_X1 port map( A1 => CU_I_n294, A2 => CU_I_n65, ZN => 
                           CU_I_n77);
   CU_I_U175 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n37, A => CU_I_n77
                           , ZN => CU_I_n211);
   CU_I_U174 : OAI21_X1 port map( B1 => CU_I_n51, B2 => CU_I_n4, A => CU_I_n167
                           , ZN => CU_I_n227);
   CU_I_U173 : OAI22_X1 port map( A1 => IRAM_DATA(0), A2 => CU_I_n290, B1 => 
                           CU_I_n291, B2 => CU_I_n119, ZN => CU_I_n135);
   CU_I_U172 : NAND4_X1 port map( A1 => CU_I_n107, A2 => IRAM_DATA(5), A3 => 
                           CU_I_n135, A4 => CU_I_n288, ZN => CU_I_n129);
   CU_I_U171 : NAND4_X1 port map( A1 => CU_I_n107, A2 => IRAM_DATA(5), A3 => 
                           IRAM_DATA(0), A4 => CU_I_n108, ZN => CU_I_n103);
   CU_I_U170 : INV_X1 port map( A => IRAM_DATA(1), ZN => CU_I_n290);
   CU_I_U169 : NAND2_X1 port map( A1 => IRAM_DATA(2), A2 => IRAM_DATA(1), ZN =>
                           CU_I_n108);
   CU_I_U168 : NAND2_X1 port map( A1 => CU_I_n25, A2 => CU_I_n64, ZN => 
                           CU_I_n83);
   CU_I_U167 : NOR2_X1 port map( A1 => IRAM_DATA(28), A2 => IRAM_DATA(29), ZN 
                           => CU_I_n201);
   CU_I_U166 : AOI21_X1 port map( B1 => IRAM_DATA(29), B2 => CU_I_n281, A => 
                           CU_I_n274, ZN => CU_I_n163);
   CU_I_U165 : INV_X1 port map( A => IRAM_DATA(2), ZN => CU_I_n289);
   CU_I_U164 : NOR4_X1 port map( A1 => CU_I_n96, A2 => CU_I_n97, A3 => CU_I_n98
                           , A4 => CU_I_n99, ZN => CU_I_n95);
   CU_I_U163 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n36, B1 =>
                           CU_I_n95, B2 => CU_I_n49, ZN => CU_I_n217);
   CU_I_U162 : INV_X1 port map( A => CU_I_n187, ZN => CU_I_n257);
   CU_I_U161 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n4, B1 => 
                           CU_I_n183, B2 => CU_I_n49, ZN => CU_I_n245);
   CU_I_U160 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n23, B1 => 
                           CU_I_n50, B2 => CU_I_n13, ZN => CU_I_n236);
   CU_I_U159 : OAI211_X1 port map( C1 => CU_I_n271, C2 => CU_I_n88, A => 
                           CU_I_n89, B => CU_I_n90, ZN => CU_I_n86);
   CU_I_U158 : AOI211_X1 port map( C1 => CU_I_n85, C2 => CU_I_n291, A => 
                           CU_I_n86, B => CU_I_n261, ZN => CU_I_n84);
   CU_I_U157 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n37, B1 =>
                           CU_I_n84, B2 => CU_I_n49, ZN => CU_I_n216);
   CU_I_U156 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n11, B1 => 
                           CU_I_n268, B2 => CU_I_n49, ZN => CU_I_n238);
   CU_I_U155 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n12, B1 => 
                           CU_I_n26, B2 => CU_I_n49, ZN => CU_I_n237);
   CU_I_U154 : INV_X1 port map( A => CU_I_n181, ZN => CU_I_n258);
   CU_I_U153 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n7, B1 => 
                           CU_I_n258, B2 => CU_I_n49, ZN => CU_I_n242);
   CU_I_U152 : NOR4_X1 port map( A1 => CU_I_n263, A2 => CU_I_n149, A3 => 
                           CU_I_n150, A4 => CU_I_n265, ZN => CU_I_n148);
   CU_I_U151 : OAI21_X1 port map( B1 => CU_I_n162, B2 => CU_I_n163, A => 
                           IRAM_DATA(31), ZN => CU_I_n146);
   CU_I_U150 : NAND4_X1 port map( A1 => CU_I_n145, A2 => CU_I_n146, A3 => 
                           CU_I_n147, A4 => CU_I_n148, ZN => CU_I_n112);
   CU_I_U149 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n27, B1 => 
                           CU_I_n50, B2 => CU_I_n15, ZN => CU_I_n254);
   CU_I_U148 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n22, B1 =>
                           CU_I_n50, B2 => CU_I_n12, ZN => CU_I_n235);
   CU_I_U147 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n21, B1 => 
                           CU_I_n50, B2 => CU_I_n11, ZN => CU_I_n234);
   CU_I_U146 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n19, B1 => 
                           CU_I_n50, B2 => CU_I_n10, ZN => CU_I_n233);
   CU_I_U145 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n17, B1 => 
                           CU_I_n50, B2 => CU_I_n9, ZN => CU_I_n232);
   CU_I_U144 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n15, B1 => 
                           CU_I_n50, B2 => CU_I_n7, ZN => CU_I_n230);
   CU_I_U143 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n30, B1 =>
                           CU_I_n50, B2 => CU_I_n21, ZN => CU_I_n225);
   CU_I_U142 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n31, B1 =>
                           CU_I_n50, B2 => CU_I_n22, ZN => CU_I_n224);
   CU_I_U141 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n32, B1 =>
                           CU_I_n50, B2 => CU_I_n23, ZN => CU_I_n223);
   CU_I_U140 : INV_X1 port map( A => CU_I_n99, ZN => CU_I_n262);
   CU_I_U139 : OAI211_X1 port map( C1 => CU_I_n113, C2 => CU_I_n114, A => 
                           CU_I_n115, B => CU_I_n262, ZN => CU_I_n110);
   CU_I_U138 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n35, B1 =>
                           CU_I_n109, B2 => CU_I_n68, ZN => CU_I_n218);
   CU_I_U137 : OAI21_X1 port map( B1 => CU_I_n139, B2 => CU_I_n114, A => 
                           CU_I_n140, ZN => CU_I_n138);
   CU_I_U136 : OAI211_X1 port map( C1 => CU_I_n278, C2 => CU_I_n116, A => 
                           CU_I_n101, B => CU_I_n269, ZN => CU_I_n137);
   CU_I_U135 : NOR3_X1 port map( A1 => CU_I_n137, A2 => CU_I_n112, A3 => 
                           CU_I_n138, ZN => CU_I_n136);
   CU_I_U134 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n33, B1 =>
                           CU_I_n136, B2 => CU_I_n67, ZN => CU_I_n220);
   CU_I_U133 : NOR3_X1 port map( A1 => CU_I_n124, A2 => CU_I_n105, A3 => 
                           CU_I_n125, ZN => CU_I_n123);
   CU_I_U132 : OAI22_X1 port map( A1 => pipe_ex_mem_en_i, A2 => CU_I_n34, B1 =>
                           CU_I_n123, B2 => CU_I_n49, ZN => CU_I_n219);
   CU_I_U131 : AOI22_X1 port map( A1 => CU_I_n69, A2 => CU_I_cw3_4_port, B1 => 
                           CU_I_n172, B2 => CU_I_cw2_4_port, ZN => CU_I_n210);
   CU_I_U130 : INV_X1 port map( A => CU_I_n210, ZN => CU_I_n72);
   CU_I_U129 : AOI22_X1 port map( A1 => CU_I_n68, A2 => CU_I_cw3_5_port, B1 => 
                           CU_I_n172, B2 => CU_I_cw2_5_port, ZN => CU_I_n208);
   CU_I_U128 : INV_X1 port map( A => CU_I_n208, ZN => CU_I_n73);
   CU_I_U127 : NOR2_X1 port map( A1 => CU_I_n266, A2 => IRAM_DATA(30), ZN => 
                           CU_I_n161);
   CU_I_U126 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n9, B1 => 
                           CU_I_n50, B2 => CU_I_n174, ZN => CU_I_n240);
   CU_I_U125 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n10, B1 => 
                           CU_I_n50, B2 => CU_I_n173, ZN => CU_I_n239);
   CU_I_U124 : OAI22_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n5, B1 => 
                           CU_I_n50, B2 => CU_I_n178, ZN => CU_I_n244);
   CU_I_U123 : INV_X1 port map( A => CU_I_n145, ZN => CU_I_n70);
   CU_I_U122 : INV_X1 port map( A => CU_I_n189, ZN => CU_I_n273);
   CU_I_U121 : NOR2_X1 port map( A1 => CU_I_n273, A2 => CU_I_n184, ZN => 
                           CU_I_n188);
   CU_I_U120 : NOR2_X1 port map( A1 => CU_I_n114, A2 => IRAM_DATA(4), ZN => 
                           CU_I_n107);
   CU_I_U119 : NOR3_X1 port map( A1 => IRAM_DATA(30), A2 => IRAM_DATA(31), A3 
                           => IRAM_DATA(29), ZN => CU_I_n202);
   CU_I_U118 : NOR3_X1 port map( A1 => CU_I_n274, A2 => IRAM_DATA(31), A3 => 
                           CU_I_n275, ZN => CU_I_n153);
   CU_I_U117 : OAI22_X1 port map( A1 => IRAM_DATA(3), A2 => CU_I_n291, B1 => 
                           CU_I_n144, B2 => CU_I_n283, ZN => CU_I_n142);
   CU_I_U116 : AOI21_X1 port map( B1 => CU_I_n106, B2 => CU_I_n119, A => 
                           CU_I_n286, ZN => CU_I_n143);
   CU_I_U115 : OAI211_X1 port map( C1 => IRAM_DATA(1), C2 => CU_I_n288, A => 
                           CU_I_n291, B => IRAM_DATA(2), ZN => CU_I_n141);
   CU_I_U114 : AOI221_X1 port map( B1 => CU_I_n141, B2 => CU_I_n284, C1 => 
                           IRAM_DATA(1), C2 => CU_I_n142, A => CU_I_n143, ZN =>
                           CU_I_n139);
   CU_I_U113 : AOI211_X1 port map( C1 => CU_I_n122, C2 => CU_I_n291, A => 
                           IRAM_DATA(4), B => CU_I_n94, ZN => CU_I_n121);
   CU_I_U112 : AOI21_X1 port map( B1 => CU_I_n291, B2 => CU_I_n288, A => 
                           CU_I_n108, ZN => CU_I_n120);
   CU_I_U111 : OAI222_X1 port map( A1 => CU_I_n288, A2 => CU_I_n119, B1 => 
                           IRAM_DATA(5), B2 => CU_I_n120, C1 => CU_I_n121, C2 
                           => CU_I_n289, ZN => CU_I_n118);
   CU_I_U110 : AOI221_X1 port map( B1 => CU_I_n106, B2 => IRAM_DATA(1), C1 => 
                           IRAM_DATA(4), C2 => CU_I_n288, A => CU_I_n118, ZN =>
                           CU_I_n113);
   CU_I_U109 : NOR2_X1 port map( A1 => IRAM_DATA(27), A2 => IRAM_DATA(26), ZN 
                           => CU_I_n160);
   CU_I_U108 : NOR3_X1 port map( A1 => CU_I_n271, A2 => IRAM_DATA(5), A3 => 
                           CU_I_n108, ZN => CU_I_n85);
   CU_I_U107 : NOR2_X1 port map( A1 => CU_I_n279, A2 => IRAM_DATA(26), ZN => 
                           CU_I_n132);
   CU_I_U106 : NOR2_X1 port map( A1 => CU_I_n282, A2 => IRAM_DATA(27), ZN => 
                           CU_I_n117);
   CU_I_U105 : INV_X1 port map( A => is_zero_i, ZN => CU_I_n76);
   CU_I_U104 : AOI22_X1 port map( A1 => is_zero_i, A2 => CU_I_cw3_4_port, B1 =>
                           CU_I_n76, B2 => CU_I_cw3_5_port, ZN => 
                           pipe_clear_n_i);
   CU_I_U103 : BUF_X1 port map( A => CU_I_n256, Z => CU_I_n57);
   CU_I_U102 : BUF_X1 port map( A => CU_I_n256, Z => CU_I_n56);
   CU_I_U101 : BUF_X1 port map( A => CU_I_n78, Z => CU_I_n60);
   CU_I_U100 : AOI22_X1 port map( A1 => CU_I_n157, A2 => CU_I_n117, B1 => 
                           CU_I_n160, B2 => CU_I_n161, ZN => CU_I_n159);
   CU_I_U99 : INV_X1 port map( A => CU_I_n159, ZN => CU_I_n259);
   CU_I_U98 : INV_X1 port map( A => CU_I_n201, ZN => CU_I_n275);
   CU_I_U97 : INV_X1 port map( A => CU_I_n85, ZN => CU_I_n270);
   CU_I_U96 : OAI21_X1 port map( B1 => CU_I_n152, B2 => CU_I_n153, A => 
                           CU_I_n154, ZN => CU_I_n151);
   CU_I_U95 : INV_X1 port map( A => CU_I_n151, ZN => CU_I_n265);
   CU_I_U94 : INV_X1 port map( A => CU_I_n107, ZN => CU_I_n271);
   CU_I_U93 : INV_X1 port map( A => DRAM_ISSUE_port, ZN => IRAM_ISSUE_port);
   CU_I_U92 : INV_X1 port map( A => CU_I_n132, ZN => CU_I_n278);
   CU_I_U91 : NAND2_X1 port map( A1 => CU_I_n176, A2 => CU_I_n132, ZN => 
                           CU_I_n189);
   CU_I_U90 : INV_X1 port map( A => CU_I_n160, ZN => CU_I_n281);
   CU_I_U89 : NOR2_X1 port map( A1 => CU_I_n281, A2 => CU_I_n116, ZN => 
                           CU_I_n149);
   CU_I_U88 : NAND2_X1 port map( A1 => CU_I_n153, A2 => CU_I_n132, ZN => 
                           CU_I_n196);
   CU_I_U87 : NAND2_X1 port map( A1 => CU_I_n160, A2 => CU_I_n207, ZN => 
                           CU_I_n115);
   CU_I_U86 : NAND2_X1 port map( A1 => CU_I_n290, A2 => CU_I_n289, ZN => 
                           CU_I_n119);
   CU_I_U85 : INV_X1 port map( A => CU_I_n106, ZN => CU_I_n287);
   CU_I_U84 : AOI21_X1 port map( B1 => CU_I_n85, B2 => CU_I_n287, A => 
                           CU_I_n105, ZN => CU_I_n104);
   CU_I_U83 : INV_X1 port map( A => pipe_clear_n_i, ZN => CU_I_n75);
   CU_I_U82 : NAND2_X1 port map( A1 => CU_I_n178, A2 => CU_I_n187, ZN => 
                           CU_I_n181);
   CU_I_U81 : NAND2_X1 port map( A1 => CU_I_n132, A2 => CU_I_n152, ZN => 
                           CU_I_n134);
   CU_I_U80 : NAND2_X1 port map( A1 => CU_I_n174, A2 => CU_I_n173, ZN => 
                           CU_I_n184);
   CU_I_U79 : NAND2_X1 port map( A1 => CU_I_n207, A2 => CU_I_n117, ZN => 
                           CU_I_n89);
   CU_I_U78 : INV_X1 port map( A => CU_I_n134, ZN => CU_I_n264);
   CU_I_U77 : NOR2_X1 port map( A1 => CU_I_n288, A2 => CU_I_n284, ZN => 
                           CU_I_n122);
   CU_I_U76 : NAND2_X1 port map( A1 => CU_I_n152, A2 => CU_I_n117, ZN => 
                           CU_I_n100);
   CU_I_U75 : INV_X1 port map( A => CU_I_n117, ZN => CU_I_n280);
   CU_I_U74 : NOR2_X1 port map( A1 => CU_I_n116, A2 => CU_I_n280, ZN => 
                           CU_I_n99);
   CU_I_U73 : NAND2_X1 port map( A1 => CU_I_n176, A2 => CU_I_n160, ZN => 
                           CU_I_n114);
   CU_I_U72 : NOR2_X1 port map( A1 => CU_I_n288, A2 => CU_I_n291, ZN => 
                           CU_I_n106);
   CU_I_U71 : NOR3_X1 port map( A1 => CU_I_n290, A2 => CU_I_n291, A3 => 
                           CU_I_n284, ZN => CU_I_n94);
   CU_I_U70 : BUF_X1 port map( A => CU_I_n56, Z => CU_I_n55);
   CU_I_U69 : BUF_X1 port map( A => CU_I_n57, Z => CU_I_n52);
   CU_I_U68 : BUF_X1 port map( A => CU_I_n56, Z => CU_I_n54);
   CU_I_U67 : BUF_X1 port map( A => CU_I_n57, Z => CU_I_n53);
   CU_I_U66 : INV_X1 port map( A => CU_I_n155, ZN => CU_I_n263);
   CU_I_U65 : INV_X1 port map( A => CU_I_n122, ZN => CU_I_n283);
   CU_I_U64 : BUF_X1 port map( A => CU_I_n58, Z => CU_I_n63);
   CU_I_U63 : INV_X1 port map( A => CU_I_n196, ZN => CU_I_n267);
   CU_I_U62 : NAND2_X1 port map( A1 => CU_I_n176, A2 => CU_I_n154, ZN => 
                           CU_I_n177);
   CU_I_U61 : BUF_X1 port map( A => CU_I_n59, Z => CU_I_n67);
   CU_I_U60 : BUF_X1 port map( A => CU_I_n59, Z => CU_I_n64);
   CU_I_U59 : BUF_X1 port map( A => CU_I_n59, Z => CU_I_n66);
   CU_I_U58 : INV_X1 port map( A => CU_I_n154, ZN => CU_I_n277);
   CU_I_U57 : BUF_X1 port map( A => CU_I_n58, Z => CU_I_n68);
   CU_I_U56 : BUF_X1 port map( A => CU_I_n58, Z => CU_I_n65);
   CU_I_U55 : NAND2_X1 port map( A1 => CU_I_n191, A2 => CU_I_n114, ZN => 
                           CU_I_n179);
   CU_I_U54 : NAND2_X1 port map( A1 => CU_I_n191, A2 => CU_I_n178, ZN => 
                           CU_I_n185);
   CU_I_U53 : NAND2_X1 port map( A1 => pipe_if_id_en_i, A2 => CU_I_n75, ZN => 
                           CU_I_n80);
   CU_I_U52 : NOR2_X1 port map( A1 => CU_I_n48, A2 => CU_I_n277, ZN => CU_I_n98
                           );
   CU_I_U51 : NOR2_X1 port map( A1 => CU_I_n283, A2 => CU_I_n114, ZN => 
                           CU_I_n91);
   CU_I_U50 : NOR2_X1 port map( A1 => CU_I_n68, A2 => CU_I_n75, ZN => CU_I_n172
                           );
   CU_I_U49 : INV_X1 port map( A => CU_I_n91, ZN => CU_I_n272);
   CU_I_U48 : INV_X1 port map( A => CU_I_n98, ZN => CU_I_n269);
   CU_I_U47 : INV_X1 port map( A => CU_I_n186, ZN => CU_I_n268);
   CU_I_U46 : INV_X1 port map( A => CU_I_n172, ZN => CU_I_n71);
   CU_I_U45 : OR2_X1 port map( A1 => CU_I_n177, A2 => CU_I_n51, ZN => CU_I_n182
                           );
   CU_I_U44 : BUF_X1 port map( A => CU_I_n71, Z => CU_I_n49);
   CU_I_U43 : BUF_X1 port map( A => CU_I_n71, Z => CU_I_n50);
   CU_I_U42 : BUF_X1 port map( A => CU_I_n71, Z => CU_I_n51);
   CU_I_U41 : CLKBUF_X1 port map( A => CU_I_n78, Z => CU_I_n59);
   CU_I_U40 : BUF_X2 port map( A => CU_I_n60, Z => CU_I_n69);
   CU_I_U39 : INV_X2 port map( A => CU_I_n58, ZN => pipe_if_id_en_i);
   CU_I_U38 : INV_X2 port map( A => IRAM_DATA(28), ZN => CU_I_n276);
   CU_I_U37 : OR4_X1 port map( A1 => CU_I_n274, A2 => CU_I_n276, A3 => 
                           IRAM_DATA(29), A4 => IRAM_DATA(31), ZN => CU_I_n48);
   CU_I_U36 : AOI211_X1 port map( C1 => CU_I_n152, C2 => CU_I_n160, A => 
                           CU_I_n41, B => CU_I_n204, ZN => CU_I_n47);
   CU_I_U35 : INV_X1 port map( A => IRAM_DATA(30), ZN => CU_I_n274);
   CU_I_U34 : AND3_X1 port map( A1 => IRAM_DATA(30), A2 => IRAM_DATA(29), A3 =>
                           IRAM_DATA(31), ZN => CU_I_n205);
   CU_I_U33 : NOR2_X1 port map( A1 => CU_I_n171, A2 => CU_I_n1, ZN => CU_I_n175
                           );
   CU_I_U32 : INV_X1 port map( A => CU_I_n43, ZN => muxA_sel_i);
   CU_I_U31 : NOR2_X1 port map( A1 => IRAM_DATA(29), A2 => IRAM_DATA(31), ZN =>
                           CU_I_n42);
   CU_I_U30 : CLKBUF_X1 port map( A => CU_I_n111, Z => CU_I_n41);
   CU_I_U29 : AND3_X1 port map( A1 => IRAM_DATA(28), A2 => IRAM_DATA(30), A3 =>
                           CU_I_n42, ZN => CU_I_n180);
   CU_I_U28 : NAND2_X2 port map( A1 => IRAM_DATA(29), A2 => CU_I_n266, ZN => 
                           CU_I_n157);
   CU_I_U27 : NAND2_X1 port map( A1 => CU_I_n26, A2 => CU_I_n14, ZN => 
                           CU_I_n171);
   CU_I_U26 : INV_X1 port map( A => CU_I_n39, ZN => alu_op_i_0_port);
   CU_I_U25 : INV_X2 port map( A => CU_I_n69, ZN => pipe_ex_mem_en_i);
   CU_I_U24 : NOR3_X1 port map( A1 => IRAM_DATA(28), A2 => IRAM_DATA(30), A3 =>
                           CU_I_n157, ZN => CU_I_n38);
   CU_I_U23 : INV_X1 port map( A => CU_I_n28, ZN => CU_I_n29);
   CU_I_U22 : NAND2_X1 port map( A1 => CU_I_n87, A2 => CU_I_n29, ZN => 
                           CU_I_n194);
   CU_I_U21 : NAND3_X1 port map( A1 => CU_I_n100, A2 => CU_I_n155, A3 => 
                           CU_I_n269, ZN => CU_I_n28);
   CU_I_U20 : OAI221_X4 port map( B1 => CU_I_n63, B2 => CU_I_n8, C1 => 
                           pipe_if_id_en_i, C2 => CU_I_n16, A => CU_I_n80, ZN 
                           => CU_I_n231);
   CU_I_U19 : AND2_X2 port map( A1 => IRAM_DATA(27), A2 => IRAM_DATA(26), ZN =>
                           CU_I_n154);
   CU_I_U18 : INV_X1 port map( A => CU_I_n45, ZN => muxB_sel_i);
   CU_I_U17 : NOR3_X1 port map( A1 => CU_I_n185, A2 => CU_I_n186, A3 => 
                           CU_I_n18, ZN => CU_I_n183);
   CU_I_U16 : INV_X1 port map( A => CU_I_n24, ZN => CU_I_n25);
   CU_I_U15 : NOR2_X1 port map( A1 => CU_I_n133, A2 => CU_I_n28, ZN => CU_I_n20
                           );
   CU_I_U14 : AND2_X1 port map( A1 => CU_I_n20, A2 => CU_I_n87, ZN => CU_I_n203
                           );
   CU_I_U13 : INV_X2 port map( A => RST, ZN => CU_I_n256);
   CU_I_U12 : OR2_X1 port map( A1 => CU_I_n184, A2 => CU_I_n257, ZN => CU_I_n18
                           );
   CU_I_U11 : AND2_X1 port map( A1 => CU_I_n178, A2 => CU_I_n177, ZN => 
                           CU_I_n14);
   CU_I_U10 : OR3_X1 port map( A1 => CU_I_n267, A2 => CU_I_n70, A3 => CU_I_n176
                           , ZN => CU_I_n1);
   CU_I_U9 : BUF_X1 port map( A => CU_I_n78, Z => CU_I_n58);
   CU_I_U8 : OAI221_X1 port map( B1 => CU_I_n188, B2 => CU_I_n51, C1 => 
                           pipe_if_id_en_i, C2 => CU_I_n3, A => CU_I_n182, ZN 
                           => CU_I_n246);
   CU_I_U7 : NOR2_X1 port map( A1 => DRAM_READY, A2 => CU_I_n27, ZN => 
                           DRAM_ISSUE_port);
   CU_I_U6 : INV_X1 port map( A => IRAM_DATA(3), ZN => CU_I_n288);
   CU_I_U5 : AND2_X1 port map( A1 => CU_I_n191, A2 => CU_I_n114, ZN => CU_I_n26
                           );
   CU_I_U4 : AND4_X1 port map( A1 => CU_I_n89, A2 => CU_I_n115, A3 => CU_I_n116
                           , A4 => CU_I_n203, ZN => CU_I_n191);
   CU_I_U3 : OAI221_X1 port map( B1 => IRAM_DATA(27), B2 => CU_I_n275, C1 => 
                           CU_I_n157, C2 => CU_I_n277, A => CU_I_n158, ZN => 
                           CU_I_n156);
   CU_I_cw1_reg_17_inst : DFFR_X1 port map( D => CU_I_n252, CK => CLK, RN => 
                           CU_I_n256, Q => rf_rs1_en_i, QN => n_1000);
   CU_I_cw1_reg_12_inst : DFFR_X1 port map( D => CU_I_n247, CK => CLK, RN => 
                           CU_I_n256, Q => regrd_sel_i, QN => n_1001);
   CU_I_cw1_reg_14_inst : DFFR_X1 port map( D => CU_I_n249, CK => CLK, RN => 
                           CU_I_n256, Q => imm_uns_i, QN => n_1002);
   CU_I_cw1_reg_15_inst : DFFR_X1 port map( D => CU_I_n250, CK => CLK, RN => 
                           CU_I_n256, Q => imm_isoff_i, QN => n_1003);
   CU_I_cw1_reg_16_inst : DFFR_X1 port map( D => CU_I_n251, CK => CLK, RN => 
                           CU_I_n256, Q => rf_rs2_en_i, QN => n_1004);
   CU_I_aluOpcode2_reg_1_inst : DFFR_X1 port map( D => CU_I_n212, CK => CLK, RN
                           => CU_I_n256, Q => alu_op_i_1_port, QN => n_1005);
   CU_I_cw2_reg_8_inst : DFFR_X1 port map( D => CU_I_n229, CK => CLK, RN => 
                           CU_I_n256, Q => npc_wb_en_i, QN => n_1006);
   CU_I_cw2_reg_9_inst : DFFR_X1 port map( D => CU_I_n228, CK => CLK, RN => 
                           CU_I_n256, Q => mem_in_en_i, QN => n_1007);
   CU_I_cw4_reg_1_inst : DFFR_X1 port map( D => CU_I_n221, CK => CLK, RN => 
                           CU_I_n256, Q => rf_we_i, QN => n_1008);
   CU_I_cw4_reg_2_inst : DFFR_X1 port map( D => CU_I_n222, CK => CLK, RN => 
                           CU_I_n256, Q => wb_mux_sel_i, QN => n_1009);
   CU_I_cw3_reg_4_inst : DFFR_X1 port map( D => CU_I_n72, CK => CLK, RN => 
                           CU_I_n256, Q => CU_I_cw3_4_port, QN => n_1010);
   CU_I_cw3_reg_5_inst : DFFR_X1 port map( D => CU_I_n73, CK => CLK, RN => 
                           CU_I_n256, Q => CU_I_cw3_5_port, QN => n_1011);
   CU_I_cw1_reg_2_inst : DFFR_X1 port map( D => CU_I_n237, CK => CLK, RN => 
                           CU_I_n256, Q => n_1012, QN => CU_I_n12);
   CU_I_cw1_reg_11_inst : DFFR_X1 port map( D => CU_I_n246, CK => CLK, RN => 
                           CU_I_n256, Q => n_1013, QN => CU_I_n3);
   CU_I_aluOpcode1_reg_0_inst : DFFR_X1 port map( D => CU_I_n216, CK => CLK, RN
                           => CU_I_n256, Q => n_1014, QN => CU_I_n37);
   CU_I_cw1_reg_8_inst : DFFR_X1 port map( D => CU_I_n243, CK => CLK, RN => 
                           CU_I_n256, Q => n_1015, QN => CU_I_n6);
   CU_I_cw1_reg_4_inst : DFFR_X1 port map( D => CU_I_n239, CK => CLK, RN => 
                           CU_I_n256, Q => n_1016, QN => CU_I_n10);
   CU_I_cw1_reg_5_inst : DFFR_X1 port map( D => CU_I_n240, CK => CLK, RN => 
                           CU_I_n256, Q => n_1017, QN => CU_I_n9);
   CU_I_cw1_reg_9_inst : DFFR_X1 port map( D => CU_I_n244, CK => CLK, RN => 
                           CU_I_n256, Q => n_1018, QN => CU_I_n5);
   CU_I_cw2_reg_1_inst : DFFR_X1 port map( D => CU_I_n236, CK => CLK, RN => 
                           CU_I_n256, Q => n_1019, QN => CU_I_n23);
   CU_I_cw2_reg_2_inst : DFFR_X1 port map( D => CU_I_n235, CK => CLK, RN => 
                           CU_I_n256, Q => n_1020, QN => CU_I_n22);
   CU_I_cw2_reg_3_inst : DFFR_X1 port map( D => CU_I_n234, CK => CLK, RN => 
                           CU_I_n256, Q => n_1021, QN => CU_I_n21);
   CU_I_cw2_reg_7_inst : DFFR_X1 port map( D => CU_I_n230, CK => CLK, RN => 
                           CU_I_n256, Q => n_1022, QN => CU_I_n15);
   CU_I_cw3_reg_1_inst : DFFR_X1 port map( D => CU_I_n223, CK => CLK, RN => 
                           CU_I_n256, Q => n_1023, QN => CU_I_n32);
   CU_I_cw3_reg_2_inst : DFFR_X1 port map( D => CU_I_n224, CK => CLK, RN => 
                           CU_I_n256, Q => n_1024, QN => CU_I_n31);
   CU_I_cw3_reg_3_inst : DFFR_X1 port map( D => CU_I_n225, CK => CLK, RN => 
                           CU_I_n256, Q => n_1025, QN => CU_I_n30);
   CU_I_cw3_reg_7_inst : DFFR_X1 port map( D => CU_I_n254, CK => CLK, RN => 
                           CU_I_n256, Q => n_1026, QN => CU_I_n27);
   CU_I_cw1_reg_3_inst : DFFR_X1 port map( D => CU_I_n238, CK => CLK, RN => 
                           CU_I_n256, Q => n_1027, QN => CU_I_n11);
   CU_I_cw1_reg_7_inst : DFFR_X1 port map( D => CU_I_n242, CK => CLK, RN => 
                           CU_I_n256, Q => n_1028, QN => CU_I_n7);
   CU_I_aluOpcode2_reg_2_inst : DFFS_X1 port map( D => CU_I_n213, CK => CLK, SN
                           => CU_I_n256, Q => alu_op_i_2_port, QN => n_1029);
   CU_I_aluOpcode2_reg_4_inst : DFFS_X2 port map( D => CU_I_n215, CK => CLK, SN
                           => CU_I_n55, Q => alu_op_i_4_port, QN => CU_I_n24);
   CU_I_U231 : NAND3_X1 port map( A1 => CU_I_n117, A2 => IRAM_DATA(28), A3 => 
                           CU_I_n205, ZN => CU_I_n130);
   CU_I_U230 : NAND3_X1 port map( A1 => CU_I_n154, A2 => CU_I_n276, A3 => 
                           CU_I_n205, ZN => CU_I_n127);
   CU_I_U229 : NAND3_X1 port map( A1 => CU_I_n132, A2 => CU_I_n276, A3 => 
                           CU_I_n205, ZN => CU_I_n140);
   CU_I_U228 : NAND3_X1 port map( A1 => CU_I_n134, A2 => CU_I_n101, A3 => 
                           CU_I_n140, ZN => CU_I_n204);
   CU_I_U227 : NAND3_X1 port map( A1 => CU_I_n160, A2 => IRAM_DATA(28), A3 => 
                           CU_I_n202, ZN => CU_I_n174);
   CU_I_U226 : NAND3_X1 port map( A1 => CU_I_n117, A2 => IRAM_DATA(28), A3 => 
                           CU_I_n202, ZN => CU_I_n173);
   CU_I_U225 : NAND3_X1 port map( A1 => CU_I_n201, A2 => CU_I_n154, A3 => 
                           CU_I_n161, ZN => CU_I_n178);
   CU_I_U224 : NAND3_X1 port map( A1 => CU_I_n189, A2 => CU_I_n196, A3 => 
                           CU_I_n177, ZN => CU_I_n186);
   CU_I_U222 : NAND3_X1 port map( A1 => IRAM_DATA(28), A2 => IRAM_DATA(29), A3 
                           => IRAM_DATA(27), ZN => CU_I_n158);
   CU_I_U221 : NAND3_X1 port map( A1 => CU_I_n129, A2 => CU_I_n130, A3 => 
                           CU_I_n131, ZN => CU_I_n124);
   CU_I_U220 : OAI33_X1 port map( A1 => CU_I_n286, A2 => CU_I_n291, A3 => 
                           CU_I_n289, B1 => IRAM_DATA(0), B2 => IRAM_DATA(4), 
                           B3 => IRAM_DATA(2), ZN => CU_I_n126);
   CU_I_U219 : OAI33_X1 port map( A1 => CU_I_n270, A2 => IRAM_DATA(0), A3 => 
                           CU_I_n288, B1 => CU_I_n272, B2 => IRAM_DATA(1), B3 
                           => CU_I_n285, ZN => CU_I_n125);
   CU_I_U218 : NAND3_X1 port map( A1 => CU_I_n103, A2 => CU_I_n89, A3 => 
                           CU_I_n104, ZN => CU_I_n96);
   CU_I_U217 : NAND3_X1 port map( A1 => CU_I_n100, A2 => CU_I_n101, A3 => 
                           CU_I_n102, ZN => CU_I_n97);
   CU_I_U216 : OAI33_X1 port map( A1 => CU_I_n286, A2 => IRAM_DATA(2), A3 => 
                           CU_I_n290, B1 => CU_I_n289, B2 => IRAM_DATA(1), B3 
                           => CU_I_n291, ZN => CU_I_n92);
   CU_I_aluOpcode2_reg_0_inst : DFFR_X1 port map( D => CU_I_n211, CK => CLK, RN
                           => CU_I_n53, Q => CU_I_n294, QN => CU_I_n39);
   CU_I_aluOpcode2_reg_3_inst : DFFR_X1 port map( D => CU_I_n214, CK => CLK, RN
                           => CU_I_n52, Q => alu_op_i_3_port, QN => n_1030);
   CU_I_aluOpcode1_reg_1_inst : DFFR_X1 port map( D => CU_I_n217, CK => CLK, RN
                           => CU_I_n52, Q => n_1031, QN => CU_I_n36);
   CU_I_aluOpcode1_reg_2_inst : DFFS_X1 port map( D => CU_I_n218, CK => CLK, SN
                           => CU_I_n55, Q => n_1032, QN => CU_I_n35);
   CU_I_aluOpcode1_reg_3_inst : DFFR_X1 port map( D => CU_I_n219, CK => CLK, RN
                           => CU_I_n52, Q => n_1033, QN => CU_I_n34);
   CU_I_aluOpcode1_reg_4_inst : DFFS_X1 port map( D => CU_I_n220, CK => CLK, SN
                           => CU_I_n55, Q => n_1034, QN => CU_I_n33);
   CU_I_cw1_reg_1_inst : DFFR_X1 port map( D => CU_I_n74, CK => CLK, RN => 
                           CU_I_n53, Q => CU_I_cw1_1_port, QN => CU_I_n13);
   CU_I_cw3_reg_6_inst : DFFS_X1 port map( D => CU_I_n253, CK => CLK, SN => 
                           CU_I_n55, Q => DRAM_READNOTWRITE_port, QN => n_1035)
                           ;
   CU_I_cw2_reg_6_inst : DFFS_X1 port map( D => CU_I_n231, CK => CLK, SN => 
                           CU_I_n55, Q => n_1036, QN => CU_I_n16);
   CU_I_cw1_reg_6_inst : DFFS_X1 port map( D => CU_I_n241, CK => CLK, SN => 
                           CU_I_n55, Q => n_1037, QN => CU_I_n8);
   CU_I_cw2_reg_10_inst : DFFR_X1 port map( D => CU_I_n227, CK => CLK, RN => 
                           CU_I_n53, Q => CU_I_n293, QN => CU_I_n45);
   CU_I_cw2_reg_11_inst : DFFR_X1 port map( D => CU_I_n226, CK => CLK, RN => 
                           CU_I_n54, Q => CU_I_n292, QN => CU_I_n43);
   CU_I_cw1_reg_13_inst : DFFR_X1 port map( D => CU_I_n248, CK => CLK, RN => 
                           CU_I_n53, Q => reg31_sel_i, QN => CU_I_n2);
   CU_I_cw1_reg_10_inst : DFFR_X1 port map( D => CU_I_n245, CK => CLK, RN => 
                           CU_I_n54, Q => n_1038, QN => CU_I_n4);
   CU_I_cw2_reg_5_inst : DFFR_X1 port map( D => CU_I_n232, CK => CLK, RN => 
                           CU_I_n54, Q => CU_I_cw2_5_port, QN => CU_I_n17);
   CU_I_cw2_reg_4_inst : DFFR_X1 port map( D => CU_I_n233, CK => CLK, RN => 
                           CU_I_n54, Q => CU_I_cw2_4_port, QN => CU_I_n19);
   CU_I_Logic0_port <= '0';
   CU_I_Logic1_port <= '1';
   dp_U792 : INV_X1 port map( A => dp_n141, ZN => dp_n941);
   dp_U791 : AOI22_X1 port map( A1 => dp_alu_out_ex_o_0_port, A2 => dp_n15, B1 
                           => dp_n17, B2 => DRAM_ADDRESS_0_port, ZN => dp_n141)
                           ;
   dp_U790 : OAI21_X1 port map( B1 => dp_n558, B2 => dp_n110, A => dp_n140, ZN 
                           => dp_n691);
   dp_U789 : NAND2_X1 port map( A1 => dp_npc_if_o_16_port, A2 => dp_n104, ZN =>
                           dp_n140);
   dp_U788 : OAI21_X1 port map( B1 => dp_n559, B2 => dp_n110, A => dp_n139, ZN 
                           => dp_n692);
   dp_U787 : NAND2_X1 port map( A1 => dp_npc_if_o_17_port, A2 => dp_n104, ZN =>
                           dp_n139);
   dp_U786 : OAI21_X1 port map( B1 => dp_n560, B2 => dp_n110, A => dp_n138, ZN 
                           => dp_n693);
   dp_U785 : NAND2_X1 port map( A1 => dp_npc_if_o_18_port, A2 => dp_n104, ZN =>
                           dp_n138);
   dp_U784 : OAI21_X1 port map( B1 => dp_n561, B2 => dp_n110, A => dp_n137, ZN 
                           => dp_n694);
   dp_U783 : NAND2_X1 port map( A1 => dp_npc_if_o_19_port, A2 => dp_n104, ZN =>
                           dp_n137);
   dp_U782 : OAI21_X1 port map( B1 => dp_n562, B2 => dp_n110, A => dp_n136, ZN 
                           => dp_n695);
   dp_U781 : NAND2_X1 port map( A1 => dp_npc_if_o_20_port, A2 => dp_n104, ZN =>
                           dp_n136);
   dp_U780 : OAI21_X1 port map( B1 => dp_n563, B2 => dp_n110, A => dp_n135, ZN 
                           => dp_n696);
   dp_U779 : NAND2_X1 port map( A1 => dp_npc_if_o_21_port, A2 => dp_n104, ZN =>
                           dp_n135);
   dp_U778 : OAI21_X1 port map( B1 => dp_n564, B2 => dp_n110, A => dp_n134, ZN 
                           => dp_n697);
   dp_U777 : NAND2_X1 port map( A1 => dp_npc_if_o_22_port, A2 => dp_n104, ZN =>
                           dp_n134);
   dp_U776 : OAI21_X1 port map( B1 => dp_n565, B2 => dp_n110, A => dp_n133, ZN 
                           => dp_n698);
   dp_U775 : NAND2_X1 port map( A1 => dp_npc_if_o_23_port, A2 => dp_n104, ZN =>
                           dp_n133);
   dp_U774 : OAI21_X1 port map( B1 => dp_n566, B2 => dp_n110, A => dp_n130, ZN 
                           => dp_n699);
   dp_U773 : NAND2_X1 port map( A1 => dp_npc_if_o_24_port, A2 => dp_n104, ZN =>
                           dp_n130);
   dp_U772 : OAI21_X1 port map( B1 => dp_n567, B2 => dp_n111, A => dp_n129, ZN 
                           => dp_n700);
   dp_U771 : NAND2_X1 port map( A1 => dp_npc_if_o_25_port, A2 => dp_n104, ZN =>
                           dp_n129);
   dp_U770 : OAI21_X1 port map( B1 => dp_n568, B2 => dp_n110, A => dp_n128, ZN 
                           => dp_n701);
   dp_U769 : NAND2_X1 port map( A1 => dp_npc_if_o_26_port, A2 => dp_n104, ZN =>
                           dp_n128);
   dp_U768 : OAI21_X1 port map( B1 => dp_n569, B2 => dp_n110, A => dp_n127, ZN 
                           => dp_n702);
   dp_U767 : NAND2_X1 port map( A1 => dp_npc_if_o_27_port, A2 => dp_n104, ZN =>
                           dp_n127);
   dp_U766 : OAI21_X1 port map( B1 => dp_n570, B2 => dp_n111, A => dp_n126, ZN 
                           => dp_n703);
   dp_U765 : NAND2_X1 port map( A1 => dp_npc_if_o_28_port, A2 => dp_n104, ZN =>
                           dp_n126);
   dp_U764 : OAI21_X1 port map( B1 => dp_n571, B2 => dp_n111, A => dp_n125, ZN 
                           => dp_n704);
   dp_U763 : NAND2_X1 port map( A1 => dp_npc_if_o_29_port, A2 => dp_n104, ZN =>
                           dp_n125);
   dp_U762 : OAI21_X1 port map( B1 => dp_n572, B2 => dp_n111, A => dp_n124, ZN 
                           => dp_n705);
   dp_U761 : NAND2_X1 port map( A1 => dp_npc_if_o_30_port, A2 => dp_n104, ZN =>
                           dp_n124);
   dp_U760 : OAI21_X1 port map( B1 => dp_n573, B2 => dp_n111, A => dp_n123, ZN 
                           => dp_n706);
   dp_U759 : NAND2_X1 port map( A1 => dp_npc_if_o_31_port, A2 => dp_n103, ZN =>
                           dp_n123);
   dp_U758 : OR2_X1 port map( A1 => pipe_if_id_en_i, A2 => dp_n142, ZN => 
                           dp_n68);
   dp_U757 : INV_X1 port map( A => pipe_clear_n_i, ZN => dp_n142);
   dp_U756 : INV_X1 port map( A => dp_n121, ZN => dp_n114);
   dp_U755 : INV_X1 port map( A => pipe_ex_mem_en_i, ZN => dp_n112);
   dp_U754 : INV_X1 port map( A => dp_n103, ZN => dp_n102);
   dp_U751 : CLKBUF_X1 port map( A => dp_n89, Z => dp_n99);
   dp_U750 : CLKBUF_X1 port map( A => dp_n22, Z => dp_n45);
   dp_U749 : CLKBUF_X1 port map( A => dp_n22, Z => dp_n44);
   dp_U748 : CLKBUF_X1 port map( A => dp_n21, Z => dp_n43);
   dp_U747 : CLKBUF_X1 port map( A => dp_n21, Z => dp_n42);
   dp_U746 : CLKBUF_X1 port map( A => dp_n21, Z => dp_n41);
   dp_U745 : CLKBUF_X1 port map( A => dp_n21, Z => dp_n40);
   dp_U744 : CLKBUF_X1 port map( A => dp_n21, Z => dp_n39);
   dp_U743 : CLKBUF_X1 port map( A => dp_n21, Z => dp_n38);
   dp_U742 : CLKBUF_X1 port map( A => dp_n20, Z => dp_n37);
   dp_U741 : CLKBUF_X1 port map( A => dp_n20, Z => dp_n36);
   dp_U740 : CLKBUF_X1 port map( A => dp_n20, Z => dp_n35);
   dp_U739 : CLKBUF_X1 port map( A => dp_n19, Z => dp_n34);
   dp_U738 : CLKBUF_X1 port map( A => dp_n19, Z => dp_n33);
   dp_U737 : CLKBUF_X1 port map( A => dp_n19, Z => dp_n32);
   dp_U736 : CLKBUF_X1 port map( A => dp_n19, Z => dp_n31);
   dp_U735 : CLKBUF_X1 port map( A => dp_n18, Z => dp_n30);
   dp_U734 : CLKBUF_X1 port map( A => dp_n18, Z => dp_n29);
   dp_U733 : CLKBUF_X1 port map( A => dp_n18, Z => dp_n28);
   dp_U732 : CLKBUF_X1 port map( A => dp_n18, Z => dp_n27);
   dp_U731 : CLKBUF_X1 port map( A => dp_n18, Z => dp_n26);
   dp_U730 : CLKBUF_X1 port map( A => dp_n18, Z => dp_n25);
   dp_U729 : OAI22_X1 port map( A1 => dp_n857, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n169, ZN => dp_n921);
   dp_U728 : OAI22_X1 port map( A1 => dp_n851, A2 => dp_n71, B1 => dp_n163, B2 
                           => dp_n67, ZN => dp_n915);
   dp_U727 : INV_X1 port map( A => dp_alu_out_ex_o_25_port, ZN => dp_n164);
   dp_U726 : OAI22_X1 port map( A1 => dp_n852, A2 => dp_n71, B1 => dp_n164, B2 
                           => dp_n67, ZN => dp_n916);
   dp_U725 : INV_X1 port map( A => dp_alu_out_ex_o_30_port, ZN => dp_n159);
   dp_U724 : OAI22_X1 port map( A1 => dp_n853, A2 => dp_n71, B1 => dp_n67, B2 
                           => dp_n165, ZN => dp_n917);
   dp_U723 : INV_X1 port map( A => dp_alu_out_ex_o_21_port, ZN => dp_n168);
   dp_U722 : INV_X1 port map( A => dp_alu_out_ex_o_29_port, ZN => dp_n160);
   dp_U721 : OAI22_X1 port map( A1 => dp_n848, A2 => dp_n71, B1 => dp_n160, B2 
                           => dp_n67, ZN => dp_n912);
   dp_U720 : INV_X1 port map( A => dp_alu_out_ex_o_28_port, ZN => dp_n161);
   dp_U719 : INV_X1 port map( A => dp_alu_out_ex_o_22_port, ZN => dp_n167);
   dp_U718 : INV_X1 port map( A => dp_alu_out_ex_o_24_port, ZN => dp_n165);
   dp_U717 : INV_X1 port map( A => dp_alu_out_ex_o_27_port, ZN => dp_n162);
   dp_U716 : OAI22_X1 port map( A1 => dp_n850, A2 => dp_n71, B1 => dp_n67, B2 
                           => dp_n162, ZN => dp_n914);
   dp_U715 : INV_X1 port map( A => dp_alu_out_ex_o_26_port, ZN => dp_n163);
   dp_U714 : OAI22_X1 port map( A1 => dp_n847, A2 => dp_n71, B1 => dp_n159, B2 
                           => dp_n67, ZN => dp_n911);
   dp_U713 : OAI22_X1 port map( A1 => dp_n856, A2 => dp_n71, B1 => dp_n67, B2 
                           => dp_n168, ZN => dp_n920);
   dp_U712 : INV_X1 port map( A => dp_alu_out_ex_o_20_port, ZN => dp_n169);
   dp_U711 : INV_X1 port map( A => dp_alu_out_ex_o_31_port, ZN => dp_n158);
   dp_U710 : INV_X1 port map( A => dp_alu_out_ex_o_23_port, ZN => dp_n166);
   dp_U709 : OAI22_X1 port map( A1 => dp_n854, A2 => dp_n71, B1 => dp_n67, B2 
                           => dp_n166, ZN => dp_n918);
   dp_U708 : OAI22_X1 port map( A1 => dp_n849, A2 => dp_n71, B1 => dp_n161, B2 
                           => dp_n67, ZN => dp_n913);
   dp_U707 : OAI22_X1 port map( A1 => dp_n855, A2 => dp_n71, B1 => dp_n167, B2 
                           => dp_n67, ZN => dp_n919);
   dp_U706 : OAI22_X1 port map( A1 => dp_n846, A2 => dp_n71, B1 => dp_n158, B2 
                           => dp_n67, ZN => dp_n910);
   dp_U705 : INV_X1 port map( A => dp_alu_out_ex_o_5_port, ZN => dp_n184);
   dp_U704 : INV_X1 port map( A => dp_alu_out_ex_o_4_port, ZN => dp_n185);
   dp_U703 : INV_X1 port map( A => wb_mux_sel_i, ZN => dp_n122);
   dp_U702 : INV_X1 port map( A => mem_in_en_i, ZN => dp_n1027);
   dp_U701 : INV_X1 port map( A => DRAM_DATA(0), ZN => dp_n400);
   dp_U700 : INV_X1 port map( A => DRAM_DATA(1), ZN => dp_n365);
   dp_U699 : INV_X1 port map( A => DRAM_DATA(2), ZN => dp_n364);
   dp_U698 : INV_X1 port map( A => DRAM_DATA(3), ZN => dp_n363);
   dp_U697 : INV_X1 port map( A => DRAM_DATA(4), ZN => dp_n362);
   dp_U696 : INV_X1 port map( A => DRAM_DATA(5), ZN => dp_n361);
   dp_U695 : INV_X1 port map( A => DRAM_DATA(6), ZN => dp_n360);
   dp_U694 : INV_X1 port map( A => DRAM_DATA(7), ZN => dp_n359);
   dp_U693 : INV_X1 port map( A => DRAM_DATA(8), ZN => dp_n358);
   dp_U692 : INV_X1 port map( A => DRAM_DATA(9), ZN => dp_n357);
   dp_U691 : INV_X1 port map( A => DRAM_DATA(10), ZN => dp_n356);
   dp_U690 : INV_X1 port map( A => DRAM_DATA(11), ZN => dp_n355);
   dp_U689 : INV_X1 port map( A => DRAM_DATA(12), ZN => dp_n354);
   dp_U688 : INV_X1 port map( A => DRAM_DATA(13), ZN => dp_n353);
   dp_U687 : INV_X1 port map( A => DRAM_DATA(14), ZN => dp_n352);
   dp_U686 : INV_X1 port map( A => DRAM_DATA(15), ZN => dp_n351);
   dp_U685 : INV_X1 port map( A => DRAM_DATA(16), ZN => dp_n350);
   dp_U684 : INV_X1 port map( A => DRAM_DATA(17), ZN => dp_n349);
   dp_U683 : INV_X1 port map( A => DRAM_DATA(18), ZN => dp_n348);
   dp_U682 : INV_X1 port map( A => DRAM_DATA(19), ZN => dp_n347);
   dp_U681 : INV_X1 port map( A => DRAM_DATA(20), ZN => dp_n346);
   dp_U680 : INV_X1 port map( A => DRAM_DATA(21), ZN => dp_n345);
   dp_U679 : INV_X1 port map( A => DRAM_DATA(22), ZN => dp_n344);
   dp_U678 : INV_X1 port map( A => DRAM_DATA(23), ZN => dp_n343);
   dp_U677 : INV_X1 port map( A => DRAM_DATA(24), ZN => dp_n342);
   dp_U676 : INV_X1 port map( A => DRAM_DATA(25), ZN => dp_n341);
   dp_U675 : INV_X1 port map( A => DRAM_DATA(26), ZN => dp_n340);
   dp_U674 : INV_X1 port map( A => DRAM_DATA(27), ZN => dp_n339);
   dp_U673 : INV_X1 port map( A => DRAM_DATA(28), ZN => dp_n338);
   dp_U672 : INV_X1 port map( A => DRAM_DATA(29), ZN => dp_n337);
   dp_U671 : INV_X1 port map( A => DRAM_DATA(30), ZN => dp_n336);
   dp_U670 : INV_X1 port map( A => DRAM_DATA(31), ZN => dp_n335);
   dp_U669 : OAI22_X1 port map( A1 => dp_n331, A2 => dp_n63, B1 => dp_n877, B2 
                           => dp_n57, ZN => dp_n909);
   dp_U668 : OAI22_X1 port map( A1 => dp_n525, A2 => dp_n65, B1 => dp_n857, B2 
                           => dp_n55, ZN => dp_n889);
   dp_U667 : OAI22_X1 port map( A1 => dp_n584, A2 => dp_n65, B1 => dp_n856, B2 
                           => dp_n55, ZN => dp_n888);
   dp_U666 : OAI22_X1 port map( A1 => dp_n585, A2 => dp_n65, B1 => dp_n855, B2 
                           => dp_n55, ZN => dp_n887);
   dp_U665 : OAI22_X1 port map( A1 => dp_n586, A2 => dp_n65, B1 => dp_n854, B2 
                           => dp_n55, ZN => dp_n886);
   dp_U664 : OAI22_X1 port map( A1 => dp_n587, A2 => dp_n65, B1 => dp_n853, B2 
                           => dp_n55, ZN => dp_n885);
   dp_U663 : OAI22_X1 port map( A1 => dp_n588, A2 => dp_n65, B1 => dp_n852, B2 
                           => dp_n55, ZN => dp_n884);
   dp_U662 : OAI22_X1 port map( A1 => dp_n589, A2 => dp_n66, B1 => dp_n851, B2 
                           => dp_n55, ZN => dp_n883);
   dp_U661 : OAI22_X1 port map( A1 => dp_n590, A2 => dp_n66, B1 => dp_n850, B2 
                           => dp_n55, ZN => dp_n882);
   dp_U660 : OAI22_X1 port map( A1 => dp_n591, A2 => dp_n66, B1 => dp_n849, B2 
                           => dp_n55, ZN => dp_n881);
   dp_U659 : OAI22_X1 port map( A1 => dp_n592, A2 => dp_n66, B1 => dp_n848, B2 
                           => dp_n55, ZN => dp_n880);
   dp_U658 : OAI22_X1 port map( A1 => dp_n593, A2 => dp_n66, B1 => dp_n847, B2 
                           => dp_n55, ZN => dp_n879);
   dp_U657 : OAI22_X1 port map( A1 => dp_n1025, A2 => dp_n61, B1 => dp_n846, B2
                           => dp_n55, ZN => dp_n878);
   dp_U656 : OAI22_X1 port map( A1 => dp_n444, A2 => dp_n91, B1 => dp_n76, B2 
                           => dp_n624, ZN => dp_n774);
   dp_U655 : OAI22_X1 port map( A1 => dp_n445, A2 => dp_n90, B1 => dp_n78, B2 
                           => dp_n625, ZN => dp_n775);
   dp_U654 : OAI22_X1 port map( A1 => dp_n447, A2 => dp_n90, B1 => dp_n81, B2 
                           => dp_n625, ZN => dp_n777);
   dp_U653 : OAI22_X1 port map( A1 => dp_n446, A2 => dp_n90, B1 => dp_n81, B2 
                           => dp_n624, ZN => dp_n776);
   dp_U652 : OAI22_X1 port map( A1 => dp_n449, A2 => dp_n94, B1 => dp_n81, B2 
                           => dp_n625, ZN => dp_n779);
   dp_U651 : INV_X1 port map( A => dp_imm_id_o_31_port, ZN => dp_n625);
   dp_U650 : OAI22_X1 port map( A1 => dp_n450, A2 => dp_n93, B1 => dp_n79, B2 
                           => dp_n625, ZN => dp_n780);
   dp_U649 : INV_X1 port map( A => dp_imm_id_o_31_port, ZN => dp_n624);
   dp_U648 : OAI22_X1 port map( A1 => dp_n448, A2 => dp_n94, B1 => dp_n80, B2 
                           => dp_n624, ZN => dp_n778);
   dp_U647 : OAI221_X1 port map( B1 => dp_n575, B2 => regrd_sel_i, C1 => 
                           dp_n574, C2 => dp_n1028, A => dp_n1026, ZN => 
                           dp_rd_fwd_id_o_0_port);
   dp_U646 : INV_X1 port map( A => dp_rd_fwd_id_o_0_port, ZN => dp_n605);
   dp_U645 : OAI22_X1 port map( A1 => dp_n93, A2 => dp_n414, B1 => dp_n80, B2 
                           => dp_n605, ZN => dp_n712);
   dp_U644 : INV_X1 port map( A => dp_imm_id_o_22_port, ZN => dp_n621);
   dp_U643 : OAI22_X1 port map( A1 => dp_n441, A2 => dp_n90, B1 => dp_n79, B2 
                           => dp_n621, ZN => dp_n771);
   dp_U642 : INV_X1 port map( A => dp_alu_out_ex_o_19_port, ZN => dp_n170);
   dp_U641 : OAI22_X1 port map( A1 => dp_n858, A2 => dp_n72, B1 => dp_n170, B2 
                           => dp_n67, ZN => dp_n922);
   dp_U640 : INV_X1 port map( A => dp_rf_out2_id_o_3_port, ZN => dp_n245);
   dp_U639 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n454, B1 => dp_n83, B2 
                           => dp_n245, ZN => dp_n784);
   dp_U638 : INV_X1 port map( A => dp_rf_out2_id_o_4_port, ZN => dp_n243);
   dp_U637 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n455, B1 => dp_n82, B2 
                           => dp_n243, ZN => dp_n785);
   dp_U636 : INV_X1 port map( A => dp_rf_out2_id_o_5_port, ZN => dp_n241);
   dp_U635 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n456, B1 => dp_n86, B2 
                           => dp_n241, ZN => dp_n786);
   dp_U634 : INV_X1 port map( A => dp_rf_out2_id_o_6_port, ZN => dp_n239);
   dp_U633 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n457, B1 => dp_n86, B2 
                           => dp_n239, ZN => dp_n787);
   dp_U632 : INV_X1 port map( A => dp_rf_out2_id_o_7_port, ZN => dp_n237);
   dp_U631 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n458, B1 => dp_n86, B2 
                           => dp_n237, ZN => dp_n788);
   dp_U630 : INV_X1 port map( A => dp_rf_out2_id_o_8_port, ZN => dp_n235);
   dp_U629 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n459, B1 => dp_n86, B2 
                           => dp_n235, ZN => dp_n789);
   dp_U628 : INV_X1 port map( A => dp_rf_out2_id_o_9_port, ZN => dp_n233);
   dp_U627 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n460, B1 => dp_n86, B2 
                           => dp_n233, ZN => dp_n790);
   dp_U626 : INV_X1 port map( A => dp_rf_out2_id_o_10_port, ZN => dp_n231);
   dp_U625 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n461, B1 => dp_n86, B2 
                           => dp_n231, ZN => dp_n791);
   dp_U624 : INV_X1 port map( A => dp_rf_out2_id_o_11_port, ZN => dp_n229);
   dp_U623 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n462, B1 => dp_n86, B2 
                           => dp_n229, ZN => dp_n792);
   dp_U622 : INV_X1 port map( A => dp_rf_out2_id_o_12_port, ZN => dp_n227);
   dp_U621 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n463, B1 => dp_n86, B2 
                           => dp_n227, ZN => dp_n793);
   dp_U620 : INV_X1 port map( A => dp_rf_out2_id_o_13_port, ZN => dp_n225);
   dp_U619 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n464, B1 => dp_n86, B2 
                           => dp_n225, ZN => dp_n794);
   dp_U618 : INV_X1 port map( A => dp_rf_out2_id_o_14_port, ZN => dp_n223);
   dp_U617 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n465, B1 => dp_n86, B2 
                           => dp_n223, ZN => dp_n795);
   dp_U616 : INV_X1 port map( A => dp_rf_out2_id_o_15_port, ZN => dp_n221);
   dp_U615 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n466, B1 => dp_n83, B2 
                           => dp_n221, ZN => dp_n796);
   dp_U614 : INV_X1 port map( A => dp_rf_out2_id_o_16_port, ZN => dp_n219);
   dp_U613 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n467, B1 => dp_n82, B2 
                           => dp_n219, ZN => dp_n797);
   dp_U612 : INV_X1 port map( A => dp_rf_out2_id_o_17_port, ZN => dp_n217);
   dp_U611 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n468, B1 => dp_n84, B2 
                           => dp_n217, ZN => dp_n798);
   dp_U610 : INV_X1 port map( A => dp_rf_out2_id_o_18_port, ZN => dp_n215);
   dp_U609 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n469, B1 => dp_n83, B2 
                           => dp_n215, ZN => dp_n799);
   dp_U608 : INV_X1 port map( A => dp_rf_out2_id_o_19_port, ZN => dp_n213);
   dp_U607 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n470, B1 => dp_n82, B2 
                           => dp_n213, ZN => dp_n800);
   dp_U606 : INV_X1 port map( A => dp_rf_out2_id_o_20_port, ZN => dp_n211);
   dp_U605 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n471, B1 => dp_n85, B2 
                           => dp_n211, ZN => dp_n801);
   dp_U604 : INV_X1 port map( A => dp_rf_out2_id_o_21_port, ZN => dp_n209);
   dp_U603 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n472, B1 => dp_n87, B2 
                           => dp_n209, ZN => dp_n802);
   dp_U602 : INV_X1 port map( A => dp_rf_out1_id_o_0_port, ZN => dp_n252);
   dp_U601 : OAI22_X1 port map( A1 => dp_n95, A2 => dp_n483, B1 => dp_n83, B2 
                           => dp_n252, ZN => dp_n813);
   dp_U600 : INV_X1 port map( A => dp_rf_out2_id_o_22_port, ZN => dp_n207);
   dp_U599 : OAI22_X1 port map( A1 => dp_n92, A2 => dp_n473, B1 => dp_n84, B2 
                           => dp_n207, ZN => dp_n803);
   dp_U598 : INV_X1 port map( A => dp_rf_out2_id_o_23_port, ZN => dp_n205);
   dp_U597 : OAI22_X1 port map( A1 => dp_n91, A2 => dp_n474, B1 => dp_n83, B2 
                           => dp_n205, ZN => dp_n804);
   dp_U596 : INV_X1 port map( A => dp_rf_out2_id_o_24_port, ZN => dp_n203);
   dp_U595 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n475, B1 => dp_n82, B2 
                           => dp_n203, ZN => dp_n805);
   dp_U594 : INV_X1 port map( A => dp_rf_out2_id_o_25_port, ZN => dp_n201);
   dp_U593 : OAI22_X1 port map( A1 => dp_n94, A2 => dp_n476, B1 => dp_n85, B2 
                           => dp_n201, ZN => dp_n806);
   dp_U592 : INV_X1 port map( A => dp_rf_out2_id_o_26_port, ZN => dp_n199);
   dp_U591 : OAI22_X1 port map( A1 => dp_n93, A2 => dp_n477, B1 => dp_n87, B2 
                           => dp_n199, ZN => dp_n807);
   dp_U590 : INV_X1 port map( A => dp_rf_out2_id_o_27_port, ZN => dp_n197);
   dp_U589 : OAI22_X1 port map( A1 => dp_n92, A2 => dp_n478, B1 => dp_n82, B2 
                           => dp_n197, ZN => dp_n808);
   dp_U588 : INV_X1 port map( A => dp_rf_out2_id_o_28_port, ZN => dp_n195);
   dp_U587 : OAI22_X1 port map( A1 => dp_n94, A2 => dp_n479, B1 => dp_n84, B2 
                           => dp_n195, ZN => dp_n809);
   dp_U586 : INV_X1 port map( A => dp_rf_out2_id_o_29_port, ZN => dp_n193);
   dp_U585 : OAI22_X1 port map( A1 => dp_n93, A2 => dp_n480, B1 => dp_n87, B2 
                           => dp_n193, ZN => dp_n810);
   dp_U584 : INV_X1 port map( A => dp_rf_out2_id_o_30_port, ZN => dp_n191);
   dp_U583 : OAI22_X1 port map( A1 => dp_n91, A2 => dp_n481, B1 => dp_n85, B2 
                           => dp_n191, ZN => dp_n811);
   dp_U582 : INV_X1 port map( A => dp_rf_out2_id_o_31_port, ZN => dp_n189);
   dp_U581 : OAI22_X1 port map( A1 => dp_n94, A2 => dp_n482, B1 => dp_n83, B2 
                           => dp_n189, ZN => dp_n812);
   dp_U580 : INV_X1 port map( A => dp_rf_out1_id_o_1_port, ZN => dp_n250);
   dp_U579 : OAI22_X1 port map( A1 => dp_n93, A2 => dp_n484, B1 => dp_n82, B2 
                           => dp_n250, ZN => dp_n814);
   dp_U578 : INV_X1 port map( A => dp_rf_out1_id_o_2_port, ZN => dp_n248);
   dp_U577 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n485, B1 => dp_n84, B2 
                           => dp_n248, ZN => dp_n815);
   dp_U576 : INV_X1 port map( A => dp_rf_out1_id_o_3_port, ZN => dp_n246);
   dp_U575 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n486, B1 => dp_n84, B2 
                           => dp_n246, ZN => dp_n816);
   dp_U574 : INV_X1 port map( A => dp_rf_out1_id_o_4_port, ZN => dp_n244);
   dp_U573 : OAI22_X1 port map( A1 => dp_n92, A2 => dp_n487, B1 => dp_n87, B2 
                           => dp_n244, ZN => dp_n817);
   dp_U572 : INV_X1 port map( A => dp_rf_out1_id_o_5_port, ZN => dp_n242);
   dp_U571 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n488, B1 => dp_n85, B2 
                           => dp_n242, ZN => dp_n818);
   dp_U570 : INV_X1 port map( A => dp_rf_out1_id_o_6_port, ZN => dp_n240);
   dp_U569 : OAI22_X1 port map( A1 => dp_n91, A2 => dp_n489, B1 => dp_n82, B2 
                           => dp_n240, ZN => dp_n819);
   dp_U568 : INV_X1 port map( A => dp_rf_out1_id_o_7_port, ZN => dp_n238);
   dp_U567 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n490, B1 => dp_n83, B2 
                           => dp_n238, ZN => dp_n820);
   dp_U566 : INV_X1 port map( A => dp_rf_out1_id_o_8_port, ZN => dp_n236);
   dp_U565 : OAI22_X1 port map( A1 => dp_n93, A2 => dp_n491, B1 => dp_n84, B2 
                           => dp_n236, ZN => dp_n821);
   dp_U564 : INV_X1 port map( A => dp_rf_out1_id_o_9_port, ZN => dp_n234);
   dp_U563 : OAI22_X1 port map( A1 => dp_n92, A2 => dp_n492, B1 => dp_n87, B2 
                           => dp_n234, ZN => dp_n822);
   dp_U562 : INV_X1 port map( A => dp_rf_out1_id_o_10_port, ZN => dp_n232);
   dp_U561 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n493, B1 => dp_n85, B2 
                           => dp_n232, ZN => dp_n823);
   dp_U560 : INV_X1 port map( A => dp_rf_out1_id_o_11_port, ZN => dp_n230);
   dp_U559 : OAI22_X1 port map( A1 => dp_n91, A2 => dp_n494, B1 => dp_n84, B2 
                           => dp_n230, ZN => dp_n824);
   dp_U558 : INV_X1 port map( A => dp_rf_out1_id_o_12_port, ZN => dp_n228);
   dp_U557 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n495, B1 => dp_n83, B2 
                           => dp_n228, ZN => dp_n825);
   dp_U556 : INV_X1 port map( A => dp_rf_out1_id_o_13_port, ZN => dp_n226);
   dp_U555 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n496, B1 => dp_n82, B2 
                           => dp_n226, ZN => dp_n826);
   dp_U554 : INV_X1 port map( A => dp_rf_out1_id_o_14_port, ZN => dp_n224);
   dp_U553 : OAI22_X1 port map( A1 => dp_n94, A2 => dp_n497, B1 => dp_n84, B2 
                           => dp_n224, ZN => dp_n827);
   dp_U552 : INV_X1 port map( A => dp_rf_out1_id_o_15_port, ZN => dp_n222);
   dp_U551 : OAI22_X1 port map( A1 => dp_n94, A2 => dp_n498, B1 => dp_n85, B2 
                           => dp_n222, ZN => dp_n828);
   dp_U550 : INV_X1 port map( A => dp_rf_out1_id_o_16_port, ZN => dp_n220);
   dp_U549 : OAI22_X1 port map( A1 => dp_n93, A2 => dp_n499, B1 => dp_n83, B2 
                           => dp_n220, ZN => dp_n829);
   dp_U548 : INV_X1 port map( A => dp_rf_out1_id_o_17_port, ZN => dp_n218);
   dp_U547 : OAI22_X1 port map( A1 => dp_n93, A2 => dp_n500, B1 => dp_n82, B2 
                           => dp_n218, ZN => dp_n830);
   dp_U546 : INV_X1 port map( A => dp_rf_out1_id_o_18_port, ZN => dp_n216);
   dp_U545 : OAI22_X1 port map( A1 => dp_n92, A2 => dp_n501, B1 => dp_n87, B2 
                           => dp_n216, ZN => dp_n831);
   dp_U544 : INV_X1 port map( A => dp_rf_out1_id_o_19_port, ZN => dp_n214);
   dp_U543 : OAI22_X1 port map( A1 => dp_n92, A2 => dp_n502, B1 => dp_n84, B2 
                           => dp_n214, ZN => dp_n832);
   dp_U542 : INV_X1 port map( A => dp_rf_out1_id_o_20_port, ZN => dp_n212);
   dp_U541 : OAI22_X1 port map( A1 => dp_n91, A2 => dp_n503, B1 => dp_n84, B2 
                           => dp_n212, ZN => dp_n833);
   dp_U540 : INV_X1 port map( A => dp_rf_out1_id_o_21_port, ZN => dp_n210);
   dp_U539 : OAI22_X1 port map( A1 => dp_n91, A2 => dp_n504, B1 => dp_n84, B2 
                           => dp_n210, ZN => dp_n834);
   dp_U538 : INV_X1 port map( A => dp_rf_out1_id_o_22_port, ZN => dp_n208);
   dp_U537 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n505, B1 => dp_n84, B2 
                           => dp_n208, ZN => dp_n835);
   dp_U536 : INV_X1 port map( A => dp_rf_out1_id_o_23_port, ZN => dp_n206);
   dp_U535 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n506, B1 => dp_n87, B2 
                           => dp_n206, ZN => dp_n836);
   dp_U534 : INV_X1 port map( A => dp_rf_out1_id_o_24_port, ZN => dp_n204);
   dp_U533 : OAI22_X1 port map( A1 => dp_n90, A2 => dp_n507, B1 => dp_n83, B2 
                           => dp_n204, ZN => dp_n837);
   dp_U532 : INV_X1 port map( A => dp_npc_id_o_3_port, ZN => dp_n629);
   dp_U531 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n263, B1 => dp_n81, B2 
                           => dp_n629, ZN => dp_n720);
   dp_U530 : INV_X1 port map( A => dp_npc_id_o_4_port, ZN => dp_n630);
   dp_U529 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n264, B1 => dp_n81, B2 
                           => dp_n630, ZN => dp_n721);
   dp_U528 : INV_X1 port map( A => dp_npc_id_o_5_port, ZN => dp_n631);
   dp_U527 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n265, B1 => dp_n76, B2 
                           => dp_n631, ZN => dp_n722);
   dp_U526 : INV_X1 port map( A => dp_npc_id_o_6_port, ZN => dp_n632);
   dp_U525 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n266, B1 => dp_n81, B2 
                           => dp_n632, ZN => dp_n723);
   dp_U524 : INV_X1 port map( A => dp_npc_id_o_7_port, ZN => dp_n633);
   dp_U523 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n267, B1 => dp_n80, B2 
                           => dp_n633, ZN => dp_n724);
   dp_U522 : INV_X1 port map( A => dp_npc_id_o_8_port, ZN => dp_n634);
   dp_U521 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n268, B1 => dp_n76, B2 
                           => dp_n634, ZN => dp_n725);
   dp_U520 : INV_X1 port map( A => dp_npc_id_o_9_port, ZN => dp_n635);
   dp_U519 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n269, B1 => dp_n76, B2 
                           => dp_n635, ZN => dp_n726);
   dp_U518 : INV_X1 port map( A => dp_npc_id_o_10_port, ZN => dp_n636);
   dp_U517 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n270, B1 => dp_n79, B2 
                           => dp_n636, ZN => dp_n727);
   dp_U516 : INV_X1 port map( A => dp_npc_id_o_11_port, ZN => dp_n637);
   dp_U515 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n271, B1 => dp_n81, B2 
                           => dp_n637, ZN => dp_n728);
   dp_U514 : INV_X1 port map( A => dp_npc_id_o_12_port, ZN => dp_n638);
   dp_U513 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n272, B1 => dp_n80, B2 
                           => dp_n638, ZN => dp_n729);
   dp_U512 : INV_X1 port map( A => dp_npc_id_o_13_port, ZN => dp_n639);
   dp_U511 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n273, B1 => dp_n79, B2 
                           => dp_n639, ZN => dp_n730);
   dp_U510 : INV_X1 port map( A => dp_npc_id_o_14_port, ZN => dp_n640);
   dp_U509 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n274, B1 => dp_n78, B2 
                           => dp_n640, ZN => dp_n731);
   dp_U508 : INV_X1 port map( A => dp_npc_id_o_15_port, ZN => dp_n641);
   dp_U507 : OAI22_X1 port map( A1 => dp_n98, A2 => dp_n275, B1 => dp_n80, B2 
                           => dp_n641, ZN => dp_n732);
   dp_U506 : INV_X1 port map( A => dp_npc_id_o_16_port, ZN => dp_n642);
   dp_U505 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n276, B1 => dp_n76, B2 
                           => dp_n642, ZN => dp_n733);
   dp_U504 : INV_X1 port map( A => dp_npc_id_o_17_port, ZN => dp_n643);
   dp_U503 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n277, B1 => dp_n77, B2 
                           => dp_n643, ZN => dp_n734);
   dp_U502 : INV_X1 port map( A => dp_npc_id_o_18_port, ZN => dp_n644);
   dp_U501 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n278, B1 => dp_n81, B2 
                           => dp_n644, ZN => dp_n735);
   dp_U500 : INV_X1 port map( A => dp_npc_id_o_19_port, ZN => dp_n645);
   dp_U499 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n279, B1 => dp_n81, B2 
                           => dp_n645, ZN => dp_n736);
   dp_U498 : INV_X1 port map( A => dp_npc_id_o_20_port, ZN => dp_n646);
   dp_U497 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n280, B1 => dp_n81, B2 
                           => dp_n646, ZN => dp_n737);
   dp_U496 : INV_X1 port map( A => dp_npc_id_o_21_port, ZN => dp_n647);
   dp_U495 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n281, B1 => dp_n76, B2 
                           => dp_n647, ZN => dp_n738);
   dp_U494 : INV_X1 port map( A => dp_npc_id_o_22_port, ZN => dp_n648);
   dp_U493 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n282, B1 => dp_n76, B2 
                           => dp_n648, ZN => dp_n739);
   dp_U492 : INV_X1 port map( A => dp_npc_id_o_23_port, ZN => dp_n1016);
   dp_U491 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n283, B1 => dp_n76, B2 
                           => dp_n1016, ZN => dp_n740);
   dp_U490 : INV_X1 port map( A => dp_npc_id_o_24_port, ZN => dp_n1017);
   dp_U489 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n284, B1 => dp_n81, B2 
                           => dp_n1017, ZN => dp_n741);
   dp_U488 : INV_X1 port map( A => dp_npc_id_o_25_port, ZN => dp_n1018);
   dp_U487 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n285, B1 => dp_n77, B2 
                           => dp_n1018, ZN => dp_n742);
   dp_U486 : INV_X1 port map( A => dp_npc_id_o_26_port, ZN => dp_n1019);
   dp_U485 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n286, B1 => dp_n81, B2 
                           => dp_n1019, ZN => dp_n743);
   dp_U484 : INV_X1 port map( A => dp_npc_id_o_27_port, ZN => dp_n1020);
   dp_U483 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n287, B1 => dp_n78, B2 
                           => dp_n1020, ZN => dp_n744);
   dp_U482 : INV_X1 port map( A => dp_npc_id_o_28_port, ZN => dp_n1021);
   dp_U481 : OAI22_X1 port map( A1 => dp_n97, A2 => dp_n288, B1 => dp_n79, B2 
                           => dp_n1021, ZN => dp_n745);
   dp_U480 : INV_X1 port map( A => dp_npc_id_o_29_port, ZN => dp_n1022);
   dp_U479 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n289, B1 => dp_n77, B2 
                           => dp_n1022, ZN => dp_n746);
   dp_U478 : INV_X1 port map( A => dp_npc_id_o_30_port, ZN => dp_n1023);
   dp_U477 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n290, B1 => dp_n77, B2 
                           => dp_n1023, ZN => dp_n747);
   dp_U476 : INV_X1 port map( A => dp_npc_id_o_31_port, ZN => dp_n1024);
   dp_U475 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n291, B1 => dp_n77, B2 
                           => dp_n1024, ZN => dp_n748);
   dp_U474 : INV_X1 port map( A => dp_imm_id_o_16_port, ZN => dp_n615);
   dp_U473 : OAI22_X1 port map( A1 => dp_n435, A2 => dp_n94, B1 => dp_n81, B2 
                           => dp_n615, ZN => dp_n765);
   dp_U472 : INV_X1 port map( A => dp_imm_id_o_19_port, ZN => dp_n618);
   dp_U471 : OAI22_X1 port map( A1 => dp_n438, A2 => dp_n93, B1 => dp_n79, B2 
                           => dp_n618, ZN => dp_n768);
   dp_U470 : INV_X1 port map( A => dp_imm_id_o_20_port, ZN => dp_n619);
   dp_U469 : OAI22_X1 port map( A1 => dp_n439, A2 => dp_n92, B1 => dp_n80, B2 
                           => dp_n619, ZN => dp_n769);
   dp_U468 : INV_X1 port map( A => dp_imm_id_o_23_port, ZN => dp_n622);
   dp_U467 : OAI22_X1 port map( A1 => dp_n442, A2 => dp_n94, B1 => dp_n80, B2 
                           => dp_n622, ZN => dp_n772);
   dp_U466 : INV_X1 port map( A => dp_imm_id_o_18_port, ZN => dp_n617);
   dp_U465 : OAI22_X1 port map( A1 => dp_n437, A2 => dp_n93, B1 => dp_n80, B2 
                           => dp_n617, ZN => dp_n767);
   dp_U464 : INV_X1 port map( A => dp_imm_id_o_21_port, ZN => dp_n620);
   dp_U463 : OAI22_X1 port map( A1 => dp_n440, A2 => dp_n92, B1 => dp_n79, B2 
                           => dp_n620, ZN => dp_n770);
   dp_U462 : INV_X1 port map( A => dp_imm_id_o_24_port, ZN => dp_n623);
   dp_U461 : OAI22_X1 port map( A1 => dp_n443, A2 => dp_n92, B1 => dp_n81, B2 
                           => dp_n623, ZN => dp_n773);
   dp_U460 : INV_X1 port map( A => dp_imm_id_o_17_port, ZN => dp_n616);
   dp_U459 : OAI22_X1 port map( A1 => dp_n436, A2 => dp_n90, B1 => dp_n80, B2 
                           => dp_n616, ZN => dp_n766);
   dp_U458 : INV_X1 port map( A => dp_rf_out1_id_o_31_port, ZN => dp_n190);
   dp_U457 : OAI22_X1 port map( A1 => dp_n94, A2 => dp_n514, B1 => dp_n85, B2 
                           => dp_n190, ZN => dp_n844);
   dp_U456 : INV_X1 port map( A => dp_rf_out1_id_o_26_port, ZN => dp_n200);
   dp_U455 : OAI22_X1 port map( A1 => dp_n92, A2 => dp_n509, B1 => dp_n82, B2 
                           => dp_n200, ZN => dp_n839);
   dp_U454 : INV_X1 port map( A => dp_rf_out1_id_o_29_port, ZN => dp_n194);
   dp_U453 : OAI22_X1 port map( A1 => dp_n91, A2 => dp_n512, B1 => dp_n85, B2 
                           => dp_n194, ZN => dp_n842);
   dp_U452 : INV_X1 port map( A => dp_rf_out1_id_o_25_port, ZN => dp_n202);
   dp_U451 : OAI22_X1 port map( A1 => dp_n94, A2 => dp_n508, B1 => dp_n85, B2 
                           => dp_n202, ZN => dp_n838);
   dp_U450 : INV_X1 port map( A => dp_rf_out1_id_o_27_port, ZN => dp_n198);
   dp_U449 : OAI22_X1 port map( A1 => dp_n92, A2 => dp_n510, B1 => dp_n84, B2 
                           => dp_n198, ZN => dp_n840);
   dp_U448 : INV_X1 port map( A => dp_rf_out1_id_o_28_port, ZN => dp_n196);
   dp_U447 : OAI22_X1 port map( A1 => dp_n93, A2 => dp_n511, B1 => dp_n87, B2 
                           => dp_n196, ZN => dp_n841);
   dp_U446 : INV_X1 port map( A => dp_rf_out1_id_o_30_port, ZN => dp_n192);
   dp_U445 : OAI22_X1 port map( A1 => dp_n91, A2 => dp_n513, B1 => dp_n84, B2 
                           => dp_n192, ZN => dp_n843);
   dp_U444 : INV_X1 port map( A => dp_rf_out2_id_o_0_port, ZN => dp_n251);
   dp_U443 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n451, B1 => dp_n77, B2 
                           => dp_n251, ZN => dp_n781);
   dp_U442 : INV_X1 port map( A => dp_rf_out2_id_o_1_port, ZN => dp_n249);
   dp_U441 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n452, B1 => dp_n78, B2 
                           => dp_n249, ZN => dp_n782);
   dp_U440 : INV_X1 port map( A => dp_rf_out2_id_o_2_port, ZN => dp_n247);
   dp_U439 : OAI22_X1 port map( A1 => dp_n96, A2 => dp_n453, B1 => dp_n78, B2 
                           => dp_n247, ZN => dp_n783);
   dp_U438 : INV_X1 port map( A => dp_imm_id_o_14_port, ZN => dp_n612);
   dp_U437 : OAI22_X1 port map( A1 => dp_n433, A2 => dp_n91, B1 => dp_n78, B2 
                           => dp_n612, ZN => dp_n763);
   dp_U436 : INV_X1 port map( A => dp_imm_id_o_1_port, ZN => dp_n595);
   dp_U435 : OAI22_X1 port map( A1 => dp_n420, A2 => dp_n93, B1 => dp_n79, B2 
                           => dp_n595, ZN => dp_n750);
   dp_U434 : INV_X1 port map( A => dp_imm_id_o_2_port, ZN => dp_n596);
   dp_U433 : OAI22_X1 port map( A1 => dp_n421, A2 => dp_n92, B1 => dp_n80, B2 
                           => dp_n596, ZN => dp_n751);
   dp_U432 : INV_X1 port map( A => dp_imm_id_o_4_port, ZN => dp_n598);
   dp_U431 : OAI22_X1 port map( A1 => dp_n423, A2 => dp_n91, B1 => dp_n76, B2 
                           => dp_n598, ZN => dp_n753);
   dp_U430 : INV_X1 port map( A => dp_imm_id_o_5_port, ZN => dp_n599);
   dp_U429 : OAI22_X1 port map( A1 => dp_n424, A2 => dp_n90, B1 => dp_n76, B2 
                           => dp_n599, ZN => dp_n754);
   dp_U428 : INV_X1 port map( A => dp_imm_id_o_7_port, ZN => dp_n601);
   dp_U427 : OAI22_X1 port map( A1 => dp_n426, A2 => dp_n94, B1 => dp_n77, B2 
                           => dp_n601, ZN => dp_n756);
   dp_U426 : INV_X1 port map( A => dp_imm_id_o_11_port, ZN => dp_n606);
   dp_U425 : OAI22_X1 port map( A1 => dp_n430, A2 => dp_n91, B1 => dp_n81, B2 
                           => dp_n606, ZN => dp_n760);
   dp_U424 : INV_X1 port map( A => dp_imm_id_o_0_port, ZN => dp_n594);
   dp_U423 : OAI22_X1 port map( A1 => dp_n419, A2 => dp_n90, B1 => dp_n81, B2 
                           => dp_n594, ZN => dp_n749);
   dp_U422 : INV_X1 port map( A => dp_imm_id_o_3_port, ZN => dp_n597);
   dp_U421 : OAI22_X1 port map( A1 => dp_n422, A2 => dp_n93, B1 => dp_n79, B2 
                           => dp_n597, ZN => dp_n752);
   dp_U420 : INV_X1 port map( A => dp_imm_id_o_6_port, ZN => dp_n600);
   dp_U419 : OAI22_X1 port map( A1 => dp_n425, A2 => dp_n92, B1 => dp_n77, B2 
                           => dp_n600, ZN => dp_n755);
   dp_U418 : INV_X1 port map( A => dp_imm_id_o_8_port, ZN => dp_n602);
   dp_U417 : OAI22_X1 port map( A1 => dp_n427, A2 => dp_n91, B1 => dp_n79, B2 
                           => dp_n602, ZN => dp_n757);
   dp_U416 : INV_X1 port map( A => dp_imm_id_o_9_port, ZN => dp_n603);
   dp_U415 : OAI22_X1 port map( A1 => dp_n428, A2 => dp_n94, B1 => dp_n81, B2 
                           => dp_n603, ZN => dp_n758);
   dp_U414 : INV_X1 port map( A => dp_imm_id_o_10_port, ZN => dp_n604);
   dp_U413 : OAI22_X1 port map( A1 => dp_n429, A2 => dp_n90, B1 => dp_n79, B2 
                           => dp_n604, ZN => dp_n759);
   dp_U412 : INV_X1 port map( A => dp_imm_id_o_12_port, ZN => dp_n608);
   dp_U411 : OAI22_X1 port map( A1 => dp_n431, A2 => dp_n90, B1 => dp_n78, B2 
                           => dp_n608, ZN => dp_n761);
   dp_U410 : INV_X1 port map( A => dp_imm_id_o_13_port, ZN => dp_n610);
   dp_U409 : OAI22_X1 port map( A1 => dp_n432, A2 => dp_n90, B1 => dp_n78, B2 
                           => dp_n610, ZN => dp_n762);
   dp_U408 : INV_X1 port map( A => dp_imm_id_o_15_port, ZN => dp_n614);
   dp_U407 : OAI22_X1 port map( A1 => dp_n434, A2 => dp_n94, B1 => dp_n77, B2 
                           => dp_n614, ZN => dp_n764);
   dp_U406 : OAI22_X1 port map( A1 => dp_n332, A2 => dp_n63, B1 => dp_n876, B2 
                           => dp_n57, ZN => dp_n908);
   dp_U405 : OAI22_X1 port map( A1 => dp_n333, A2 => dp_n64, B1 => dp_n875, B2 
                           => dp_n57, ZN => dp_n907);
   dp_U404 : OAI22_X1 port map( A1 => dp_n334, A2 => dp_n64, B1 => dp_n874, B2 
                           => dp_n57, ZN => dp_n906);
   dp_U403 : OAI22_X1 port map( A1 => dp_n402, A2 => dp_n64, B1 => dp_n873, B2 
                           => dp_n57, ZN => dp_n905);
   dp_U402 : OAI22_X1 port map( A1 => dp_n403, A2 => dp_n64, B1 => dp_n872, B2 
                           => dp_n57, ZN => dp_n904);
   dp_U401 : OAI22_X1 port map( A1 => dp_n404, A2 => dp_n64, B1 => dp_n871, B2 
                           => dp_n57, ZN => dp_n903);
   dp_U400 : OAI22_X1 port map( A1 => dp_n405, A2 => dp_n64, B1 => dp_n870, B2 
                           => dp_n57, ZN => dp_n902);
   dp_U399 : OAI22_X1 port map( A1 => dp_n406, A2 => dp_n64, B1 => dp_n869, B2 
                           => dp_n56, ZN => dp_n901);
   dp_U398 : OAI22_X1 port map( A1 => dp_n407, A2 => dp_n64, B1 => dp_n868, B2 
                           => dp_n56, ZN => dp_n900);
   dp_U397 : OAI22_X1 port map( A1 => dp_n408, A2 => dp_n64, B1 => dp_n867, B2 
                           => dp_n56, ZN => dp_n899);
   dp_U396 : OAI22_X1 port map( A1 => dp_n409, A2 => dp_n64, B1 => dp_n866, B2 
                           => dp_n56, ZN => dp_n898);
   dp_U395 : OAI22_X1 port map( A1 => dp_n410, A2 => dp_n64, B1 => dp_n865, B2 
                           => dp_n56, ZN => dp_n897);
   dp_U394 : OAI22_X1 port map( A1 => dp_n411, A2 => dp_n64, B1 => dp_n864, B2 
                           => dp_n56, ZN => dp_n896);
   dp_U393 : OAI22_X1 port map( A1 => dp_n412, A2 => dp_n65, B1 => dp_n863, B2 
                           => dp_n56, ZN => dp_n895);
   dp_U392 : OAI22_X1 port map( A1 => dp_n413, A2 => dp_n65, B1 => dp_n862, B2 
                           => dp_n56, ZN => dp_n894);
   dp_U391 : OAI22_X1 port map( A1 => dp_n517, A2 => dp_n65, B1 => dp_n861, B2 
                           => dp_n56, ZN => dp_n893);
   dp_U390 : OAI22_X1 port map( A1 => dp_n519, A2 => dp_n65, B1 => dp_n860, B2 
                           => dp_n56, ZN => dp_n892);
   dp_U389 : OAI22_X1 port map( A1 => dp_n521, A2 => dp_n65, B1 => dp_n859, B2 
                           => dp_n56, ZN => dp_n891);
   dp_U388 : OAI22_X1 port map( A1 => dp_n523, A2 => dp_n65, B1 => dp_n858, B2 
                           => dp_n56, ZN => dp_n890);
   dp_U387 : INV_X1 port map( A => reg31_sel_i, ZN => dp_n1026);
   dp_U386 : INV_X1 port map( A => regrd_sel_i, ZN => dp_n1028);
   dp_U385 : INV_X1 port map( A => dp_npc_if_o_10_port, ZN => dp_n148);
   dp_U384 : OAI22_X1 port map( A1 => dp_n110, A2 => dp_n552, B1 => dp_n102, B2
                           => dp_n148, ZN => dp_n685);
   dp_U383 : INV_X1 port map( A => dp_npc_if_o_11_port, ZN => dp_n147);
   dp_U382 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n553, B1 => dp_n4, B2 
                           => dp_n147, ZN => dp_n686);
   dp_U381 : INV_X1 port map( A => dp_npc_if_o_12_port, ZN => dp_n146);
   dp_U380 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n554, B1 => dp_n101, B2
                           => dp_n146, ZN => dp_n687);
   dp_U379 : INV_X1 port map( A => dp_npc_if_o_13_port, ZN => dp_n145);
   dp_U378 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n555, B1 => dp_n4, B2 
                           => dp_n145, ZN => dp_n688);
   dp_U377 : INV_X1 port map( A => dp_npc_if_o_14_port, ZN => dp_n144);
   dp_U376 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n556, B1 => dp_n100, B2
                           => dp_n144, ZN => dp_n689);
   dp_U375 : INV_X1 port map( A => dp_npc_if_o_15_port, ZN => dp_n143);
   dp_U374 : OAI22_X1 port map( A1 => dp_n110, A2 => dp_n557, B1 => dp_n102, B2
                           => dp_n143, ZN => dp_n690);
   dp_U373 : INV_X1 port map( A => dp_npc_if_o_0_port, ZN => dp_n253);
   dp_U372 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n542, B1 => dp_n4, B2 
                           => dp_n253, ZN => dp_n675);
   dp_U371 : INV_X1 port map( A => dp_npc_if_o_1_port, ZN => dp_n157);
   dp_U370 : OAI22_X1 port map( A1 => dp_n110, A2 => dp_n543, B1 => dp_n3, B2 
                           => dp_n157, ZN => dp_n676);
   dp_U369 : INV_X1 port map( A => dp_npc_if_o_2_port, ZN => dp_n156);
   dp_U368 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n544, B1 => dp_n4, B2 
                           => dp_n156, ZN => dp_n677);
   dp_U367 : INV_X1 port map( A => dp_npc_if_o_3_port, ZN => dp_n155);
   dp_U366 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n545, B1 => dp_n101, B2
                           => dp_n155, ZN => dp_n678);
   dp_U365 : INV_X1 port map( A => dp_npc_if_o_4_port, ZN => dp_n154);
   dp_U364 : OAI22_X1 port map( A1 => dp_n110, A2 => dp_n546, B1 => dp_n101, B2
                           => dp_n154, ZN => dp_n679);
   dp_U363 : INV_X1 port map( A => dp_npc_if_o_5_port, ZN => dp_n153);
   dp_U362 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n547, B1 => dp_n100, B2
                           => dp_n153, ZN => dp_n680);
   dp_U361 : INV_X1 port map( A => dp_npc_if_o_6_port, ZN => dp_n152);
   dp_U360 : OAI22_X1 port map( A1 => dp_n110, A2 => dp_n548, B1 => dp_n101, B2
                           => dp_n152, ZN => dp_n681);
   dp_U359 : INV_X1 port map( A => dp_npc_if_o_7_port, ZN => dp_n151);
   dp_U358 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n549, B1 => dp_n3, B2 
                           => dp_n151, ZN => dp_n682);
   dp_U357 : INV_X1 port map( A => dp_npc_if_o_8_port, ZN => dp_n150);
   dp_U356 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n550, B1 => dp_n3, B2 
                           => dp_n150, ZN => dp_n683);
   dp_U355 : INV_X1 port map( A => dp_npc_if_o_9_port, ZN => dp_n149);
   dp_U354 : OAI22_X1 port map( A1 => dp_n109, A2 => dp_n551, B1 => dp_n3, B2 
                           => dp_n149, ZN => dp_n684);
   dp_U353 : INV_X1 port map( A => IRAM_DATA(0), ZN => dp_n1055);
   dp_U352 : OAI22_X1 port map( A1 => dp_n526, A2 => dp_n107, B1 => dp_n100, B2
                           => dp_n1055, ZN => dp_n649);
   dp_U351 : INV_X1 port map( A => IRAM_DATA(1), ZN => dp_n1054);
   dp_U350 : OAI22_X1 port map( A1 => dp_n527, A2 => dp_n107, B1 => dp_n101, B2
                           => dp_n1054, ZN => dp_n650);
   dp_U349 : INV_X1 port map( A => IRAM_DATA(2), ZN => dp_n1053);
   dp_U348 : OAI22_X1 port map( A1 => dp_n528, A2 => dp_n107, B1 => dp_n69, B2 
                           => dp_n1053, ZN => dp_n651);
   dp_U347 : INV_X1 port map( A => IRAM_DATA(3), ZN => dp_n1052);
   dp_U346 : OAI22_X1 port map( A1 => dp_n529, A2 => dp_n108, B1 => dp_n3, B2 
                           => dp_n1052, ZN => dp_n652);
   dp_U345 : INV_X1 port map( A => IRAM_DATA(4), ZN => dp_n1051);
   dp_U344 : OAI22_X1 port map( A1 => dp_n530, A2 => dp_n108, B1 => dp_n4, B2 
                           => dp_n1051, ZN => dp_n653);
   dp_U343 : INV_X1 port map( A => IRAM_DATA(5), ZN => dp_n1050);
   dp_U342 : OAI22_X1 port map( A1 => dp_n531, A2 => dp_n107, B1 => dp_n3, B2 
                           => dp_n1050, ZN => dp_n654);
   dp_U341 : INV_X1 port map( A => IRAM_DATA(6), ZN => dp_n1049);
   dp_U340 : OAI22_X1 port map( A1 => dp_n532, A2 => dp_n108, B1 => dp_n100, B2
                           => dp_n1049, ZN => dp_n655);
   dp_U339 : INV_X1 port map( A => IRAM_DATA(7), ZN => dp_n1048);
   dp_U338 : OAI22_X1 port map( A1 => dp_n533, A2 => dp_n107, B1 => dp_n100, B2
                           => dp_n1048, ZN => dp_n656);
   dp_U337 : INV_X1 port map( A => IRAM_DATA(8), ZN => dp_n1047);
   dp_U336 : OAI22_X1 port map( A1 => dp_n534, A2 => dp_n107, B1 => dp_n102, B2
                           => dp_n1047, ZN => dp_n657);
   dp_U335 : INV_X1 port map( A => IRAM_DATA(9), ZN => dp_n1046);
   dp_U334 : OAI22_X1 port map( A1 => dp_n535, A2 => dp_n108, B1 => dp_n4, B2 
                           => dp_n1046, ZN => dp_n658);
   dp_U333 : INV_X1 port map( A => IRAM_DATA(10), ZN => dp_n1045);
   dp_U332 : OAI22_X1 port map( A1 => dp_n536, A2 => dp_n108, B1 => dp_n69, B2 
                           => dp_n1045, ZN => dp_n659);
   dp_U331 : INV_X1 port map( A => IRAM_DATA(11), ZN => dp_n1044);
   dp_U330 : OAI22_X1 port map( A1 => dp_n575, A2 => dp_n107, B1 => dp_n100, B2
                           => dp_n1044, ZN => dp_n660);
   dp_U329 : INV_X1 port map( A => IRAM_DATA(12), ZN => dp_n1043);
   dp_U328 : OAI22_X1 port map( A1 => dp_n577, A2 => dp_n108, B1 => dp_n4, B2 
                           => dp_n1043, ZN => dp_n661);
   dp_U327 : INV_X1 port map( A => IRAM_DATA(13), ZN => dp_n1042);
   dp_U326 : OAI22_X1 port map( A1 => dp_n579, A2 => dp_n108, B1 => dp_n100, B2
                           => dp_n1042, ZN => dp_n662);
   dp_U325 : INV_X1 port map( A => IRAM_DATA(14), ZN => dp_n1041);
   dp_U324 : OAI22_X1 port map( A1 => dp_n581, A2 => dp_n107, B1 => dp_n101, B2
                           => dp_n1041, ZN => dp_n663);
   dp_U323 : INV_X1 port map( A => IRAM_DATA(15), ZN => dp_n1040);
   dp_U322 : OAI22_X1 port map( A1 => dp_n583, A2 => dp_n107, B1 => dp_n69, B2 
                           => dp_n1040, ZN => dp_n664);
   dp_U321 : INV_X1 port map( A => IRAM_DATA(16), ZN => dp_n1039);
   dp_U320 : OAI22_X1 port map( A1 => dp_n574, A2 => dp_n108, B1 => dp_n102, B2
                           => dp_n1039, ZN => dp_n665);
   dp_U319 : INV_X1 port map( A => IRAM_DATA(17), ZN => dp_n1038);
   dp_U318 : OAI22_X1 port map( A1 => dp_n576, A2 => dp_n108, B1 => dp_n102, B2
                           => dp_n1038, ZN => dp_n666);
   dp_U317 : INV_X1 port map( A => IRAM_DATA(18), ZN => dp_n1037);
   dp_U316 : OAI22_X1 port map( A1 => dp_n578, A2 => dp_n108, B1 => dp_n101, B2
                           => dp_n1037, ZN => dp_n667);
   dp_U315 : INV_X1 port map( A => IRAM_DATA(19), ZN => dp_n1036);
   dp_U314 : OAI22_X1 port map( A1 => dp_n580, A2 => dp_n108, B1 => dp_n69, B2 
                           => dp_n1036, ZN => dp_n668);
   dp_U313 : INV_X1 port map( A => IRAM_DATA(20), ZN => dp_n1035);
   dp_U312 : OAI22_X1 port map( A1 => dp_n582, A2 => dp_n108, B1 => dp_n102, B2
                           => dp_n1035, ZN => dp_n669);
   dp_U311 : INV_X1 port map( A => IRAM_DATA(23), ZN => dp_n1032);
   dp_U310 : OAI22_X1 port map( A1 => dp_n539, A2 => dp_n107, B1 => dp_n3, B2 
                           => dp_n1032, ZN => dp_n672);
   dp_U309 : INV_X1 port map( A => IRAM_DATA(24), ZN => dp_n1031);
   dp_U308 : OAI22_X1 port map( A1 => dp_n540, A2 => dp_n107, B1 => dp_n69, B2 
                           => dp_n1031, ZN => dp_n673);
   dp_U307 : INV_X1 port map( A => IRAM_DATA(25), ZN => dp_n1030);
   dp_U306 : OAI22_X1 port map( A1 => dp_n541, A2 => dp_n107, B1 => dp_n102, B2
                           => dp_n1030, ZN => dp_n674);
   dp_U305 : INV_X1 port map( A => IRAM_DATA(21), ZN => dp_n1034);
   dp_U304 : OAI22_X1 port map( A1 => dp_n537, A2 => dp_n109, B1 => dp_n101, B2
                           => dp_n1034, ZN => dp_n670);
   dp_U303 : INV_X1 port map( A => IRAM_DATA(22), ZN => dp_n1033);
   dp_U302 : OAI22_X1 port map( A1 => dp_n538, A2 => dp_n109, B1 => dp_n3, B2 
                           => dp_n1033, ZN => dp_n671);
   dp_U301 : INV_X1 port map( A => dp_alu_out_ex_o_7_port, ZN => dp_n182);
   dp_U300 : OAI22_X1 port map( A1 => dp_n870, A2 => dp_n73, B1 => dp_n67, B2 
                           => dp_n182, ZN => dp_n934);
   dp_U299 : INV_X1 port map( A => dp_alu_out_ex_o_18_port, ZN => dp_n171);
   dp_U298 : OAI22_X1 port map( A1 => dp_n859, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n171, ZN => dp_n923);
   dp_U297 : INV_X1 port map( A => dp_alu_out_ex_o_13_port, ZN => dp_n176);
   dp_U296 : OAI22_X1 port map( A1 => dp_n864, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n176, ZN => dp_n928);
   dp_U295 : INV_X1 port map( A => dp_alu_out_ex_o_14_port, ZN => dp_n175);
   dp_U294 : OAI22_X1 port map( A1 => dp_n863, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n175, ZN => dp_n927);
   dp_U293 : INV_X1 port map( A => dp_alu_out_ex_o_15_port, ZN => dp_n174);
   dp_U292 : OAI22_X1 port map( A1 => dp_n862, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n174, ZN => dp_n926);
   dp_U291 : INV_X1 port map( A => dp_alu_out_ex_o_9_port, ZN => dp_n180);
   dp_U290 : OAI22_X1 port map( A1 => dp_n868, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n180, ZN => dp_n932);
   dp_U289 : INV_X1 port map( A => dp_alu_out_ex_o_8_port, ZN => dp_n181);
   dp_U288 : OAI22_X1 port map( A1 => dp_n869, A2 => dp_n73, B1 => dp_n67, B2 
                           => dp_n181, ZN => dp_n933);
   dp_U287 : INV_X1 port map( A => dp_alu_out_ex_o_10_port, ZN => dp_n179);
   dp_U286 : OAI22_X1 port map( A1 => dp_n867, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n179, ZN => dp_n931);
   dp_U285 : INV_X1 port map( A => dp_alu_out_ex_o_17_port, ZN => dp_n172);
   dp_U284 : OAI22_X1 port map( A1 => dp_n860, A2 => dp_n72, B1 => dp_n172, B2 
                           => dp_n67, ZN => dp_n924);
   dp_U283 : INV_X1 port map( A => dp_alu_out_ex_o_11_port, ZN => dp_n178);
   dp_U282 : OAI22_X1 port map( A1 => dp_n866, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n178, ZN => dp_n930);
   dp_U281 : INV_X1 port map( A => dp_alu_out_ex_o_12_port, ZN => dp_n177);
   dp_U280 : OAI22_X1 port map( A1 => dp_n865, A2 => dp_n72, B1 => dp_n67, B2 
                           => dp_n177, ZN => dp_n929);
   dp_U279 : INV_X1 port map( A => dp_alu_out_ex_o_16_port, ZN => dp_n173);
   dp_U278 : OAI22_X1 port map( A1 => dp_n861, A2 => dp_n72, B1 => dp_n173, B2 
                           => dp_n67, ZN => dp_n925);
   dp_U277 : INV_X1 port map( A => dp_rd_fwd_ex_o_0_port, ZN => dp_n255);
   dp_U276 : OAI22_X1 port map( A1 => dp_n71, A2 => dp_n293, B1 => dp_n67, B2 
                           => dp_n255, ZN => dp_n1014);
   dp_U275 : OAI22_X1 port map( A1 => dp_n872, A2 => dp_n73, B1 => dp_n67, B2 
                           => dp_n184, ZN => dp_n936);
   dp_U274 : INV_X1 port map( A => dp_alu_out_ex_o_3_port, ZN => dp_n186);
   dp_U273 : OAI22_X1 port map( A1 => dp_n874, A2 => dp_n73, B1 => dp_n67, B2 
                           => dp_n186, ZN => dp_n938);
   dp_U272 : INV_X1 port map( A => dp_alu_out_ex_o_2_port, ZN => dp_n187);
   dp_U271 : OAI22_X1 port map( A1 => dp_n875, A2 => dp_n73, B1 => dp_n67, B2 
                           => dp_n187, ZN => dp_n939);
   dp_U270 : INV_X1 port map( A => dp_branch_t_ex_o, ZN => dp_n292);
   dp_U269 : OAI22_X1 port map( A1 => dp_n515, A2 => dp_n71, B1 => dp_n67, B2 
                           => dp_n292, ZN => dp_n845);
   dp_U268 : INV_X1 port map( A => dp_rd_fwd_ex_o_1_port, ZN => dp_n256);
   dp_U267 : OAI22_X1 port map( A1 => dp_n73, A2 => dp_n294, B1 => dp_n67, B2 
                           => dp_n256, ZN => dp_n1013);
   dp_U266 : INV_X1 port map( A => dp_rd_fwd_ex_o_2_port, ZN => dp_n257);
   dp_U265 : OAI22_X1 port map( A1 => dp_n73, A2 => dp_n295, B1 => dp_n67, B2 
                           => dp_n257, ZN => dp_n1012);
   dp_U264 : INV_X1 port map( A => dp_rd_fwd_ex_o_3_port, ZN => dp_n258);
   dp_U263 : OAI22_X1 port map( A1 => dp_n73, A2 => dp_n296, B1 => dp_n67, B2 
                           => dp_n258, ZN => dp_n1011);
   dp_U262 : INV_X1 port map( A => dp_rd_fwd_ex_o_4_port, ZN => dp_n259);
   dp_U261 : OAI22_X1 port map( A1 => dp_n73, A2 => dp_n297, B1 => dp_n67, B2 
                           => dp_n259, ZN => dp_n1010);
   dp_U260 : OAI22_X1 port map( A1 => dp_n873, A2 => dp_n73, B1 => dp_n67, B2 
                           => dp_n185, ZN => dp_n937);
   dp_U259 : INV_X1 port map( A => dp_alu_out_ex_o_1_port, ZN => dp_n188);
   dp_U258 : OAI22_X1 port map( A1 => dp_n876, A2 => dp_n73, B1 => dp_n67, B2 
                           => dp_n188, ZN => dp_n940);
   dp_U257 : INV_X1 port map( A => dp_alu_out_ex_o_6_port, ZN => dp_n183);
   dp_U256 : OAI22_X1 port map( A1 => dp_n871, A2 => dp_n73, B1 => dp_n67, B2 
                           => dp_n183, ZN => dp_n935);
   dp_U255 : OAI221_X1 port map( B1 => dp_n577, B2 => regrd_sel_i, C1 => 
                           dp_n576, C2 => dp_n1028, A => dp_n1026, ZN => 
                           dp_rd_fwd_id_o_1_port);
   dp_U254 : INV_X1 port map( A => dp_rd_fwd_id_o_1_port, ZN => dp_n607);
   dp_U253 : OAI22_X1 port map( A1 => dp_n99, A2 => dp_n415, B1 => dp_n77, B2 
                           => dp_n607, ZN => dp_n713);
   dp_U252 : OAI221_X1 port map( B1 => dp_n579, B2 => regrd_sel_i, C1 => 
                           dp_n578, C2 => dp_n1028, A => dp_n1026, ZN => 
                           dp_rd_fwd_id_o_2_port);
   dp_U251 : INV_X1 port map( A => dp_rd_fwd_id_o_2_port, ZN => dp_n609);
   dp_U250 : OAI22_X1 port map( A1 => dp_n99, A2 => dp_n416, B1 => dp_n80, B2 
                           => dp_n609, ZN => dp_n714);
   dp_U249 : OAI221_X1 port map( B1 => dp_n581, B2 => regrd_sel_i, C1 => 
                           dp_n580, C2 => dp_n1028, A => dp_n1026, ZN => 
                           dp_rd_fwd_id_o_3_port);
   dp_U248 : INV_X1 port map( A => dp_rd_fwd_id_o_3_port, ZN => dp_n611);
   dp_U247 : OAI22_X1 port map( A1 => dp_n99, A2 => dp_n417, B1 => dp_n76, B2 
                           => dp_n611, ZN => dp_n715);
   dp_U246 : OAI221_X1 port map( B1 => dp_n583, B2 => regrd_sel_i, C1 => 
                           dp_n582, C2 => dp_n1028, A => dp_n1026, ZN => 
                           dp_rd_fwd_id_o_4_port);
   dp_U245 : INV_X1 port map( A => dp_rd_fwd_id_o_4_port, ZN => dp_n613);
   dp_U244 : OAI22_X1 port map( A1 => dp_n99, A2 => dp_n418, B1 => dp_n78, B2 
                           => dp_n613, ZN => dp_n716);
   dp_U243 : INV_X1 port map( A => dp_npc_id_o_0_port, ZN => dp_n626);
   dp_U242 : OAI22_X1 port map( A1 => dp_n99, A2 => dp_n260, B1 => dp_n77, B2 
                           => dp_n626, ZN => dp_n717);
   dp_U241 : INV_X1 port map( A => dp_npc_id_o_1_port, ZN => dp_n627);
   dp_U240 : OAI22_X1 port map( A1 => dp_n99, A2 => dp_n261, B1 => dp_n78, B2 
                           => dp_n627, ZN => dp_n718);
   dp_U239 : INV_X1 port map( A => dp_npc_id_o_2_port, ZN => dp_n628);
   dp_U238 : OAI22_X1 port map( A1 => dp_n99, A2 => dp_n262, B1 => dp_n78, B2 
                           => dp_n628, ZN => dp_n719);
   dp_U237 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_8_port, A2 => dp_n51, B1
                           => dp_z_word_8_port, B2 => dp_n47, ZN => dp_n392);
   dp_U236 : OAI221_X1 port map( B1 => dp_n268, B2 => dp_n53, C1 => dp_n72, C2 
                           => dp_n358, A => dp_n392, ZN => dp_n996);
   dp_U235 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_9_port, A2 => dp_n50, B1
                           => dp_z_word_9_port, B2 => dp_n47, ZN => dp_n391);
   dp_U234 : OAI221_X1 port map( B1 => dp_n269, B2 => dp_n53, C1 => dp_n73, C2 
                           => dp_n357, A => dp_n391, ZN => dp_n995);
   dp_U233 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_10_port, A2 => dp_n50, 
                           B1 => dp_z_word_10_port, B2 => dp_n47, ZN => dp_n390
                           );
   dp_U232 : OAI221_X1 port map( B1 => dp_n270, B2 => dp_n53, C1 => dp_n71, C2 
                           => dp_n356, A => dp_n390, ZN => dp_n994);
   dp_U231 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_11_port, A2 => dp_n49, 
                           B1 => dp_z_word_11_port, B2 => dp_n47, ZN => dp_n389
                           );
   dp_U230 : OAI221_X1 port map( B1 => dp_n271, B2 => dp_n53, C1 => dp_n72, C2 
                           => dp_n355, A => dp_n389, ZN => dp_n993);
   dp_U229 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_12_port, A2 => dp_n51, 
                           B1 => dp_z_word_12_port, B2 => dp_n47, ZN => dp_n388
                           );
   dp_U228 : OAI221_X1 port map( B1 => dp_n272, B2 => dp_n53, C1 => dp_n73, C2 
                           => dp_n354, A => dp_n388, ZN => dp_n992);
   dp_U227 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_13_port, A2 => dp_n49, 
                           B1 => dp_z_word_13_port, B2 => dp_n47, ZN => dp_n387
                           );
   dp_U226 : OAI221_X1 port map( B1 => dp_n273, B2 => dp_n53, C1 => dp_n73, C2 
                           => dp_n353, A => dp_n387, ZN => dp_n991);
   dp_U225 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_14_port, A2 => dp_n51, 
                           B1 => dp_z_word_14_port, B2 => dp_n47, ZN => dp_n386
                           );
   dp_U224 : OAI221_X1 port map( B1 => dp_n274, B2 => dp_n53, C1 => dp_n73, C2 
                           => dp_n352, A => dp_n386, ZN => dp_n990);
   dp_U223 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_15_port, A2 => dp_n49, 
                           B1 => dp_z_word_15_port, B2 => dp_n47, ZN => dp_n385
                           );
   dp_U222 : OAI221_X1 port map( B1 => dp_n275, B2 => dp_n53, C1 => dp_n71, C2 
                           => dp_n351, A => dp_n385, ZN => dp_n989);
   dp_U221 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_16_port, A2 => dp_n51, 
                           B1 => dp_z_word_16_port, B2 => dp_n47, ZN => dp_n384
                           );
   dp_U220 : OAI221_X1 port map( B1 => dp_n276, B2 => dp_n53, C1 => dp_n72, C2 
                           => dp_n350, A => dp_n384, ZN => dp_n988);
   dp_U219 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_17_port, A2 => dp_n49, 
                           B1 => dp_z_word_17_port, B2 => dp_n47, ZN => dp_n383
                           );
   dp_U218 : OAI221_X1 port map( B1 => dp_n277, B2 => dp_n53, C1 => dp_n71, C2 
                           => dp_n349, A => dp_n383, ZN => dp_n987);
   dp_U217 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_18_port, A2 => dp_n51, 
                           B1 => dp_z_word_18_port, B2 => dp_n47, ZN => dp_n382
                           );
   dp_U216 : OAI221_X1 port map( B1 => dp_n278, B2 => dp_n53, C1 => dp_n73, C2 
                           => dp_n348, A => dp_n382, ZN => dp_n986);
   dp_U215 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_19_port, A2 => dp_n49, 
                           B1 => dp_z_word_19_port, B2 => dp_n47, ZN => dp_n381
                           );
   dp_U214 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_20_port, A2 => dp_n49, 
                           B1 => dp_z_word_20_port, B2 => dp_n46, ZN => dp_n380
                           );
   dp_U213 : OAI221_X1 port map( B1 => dp_n280, B2 => dp_n52, C1 => dp_n71, C2 
                           => dp_n346, A => dp_n380, ZN => dp_n984);
   dp_U212 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_21_port, A2 => dp_n51, 
                           B1 => dp_z_word_21_port, B2 => dp_n46, ZN => dp_n379
                           );
   dp_U211 : OAI221_X1 port map( B1 => dp_n281, B2 => dp_n52, C1 => dp_n73, C2 
                           => dp_n345, A => dp_n379, ZN => dp_n983);
   dp_U210 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_22_port, A2 => dp_n49, 
                           B1 => dp_z_word_22_port, B2 => dp_n46, ZN => dp_n378
                           );
   dp_U209 : OAI221_X1 port map( B1 => dp_n282, B2 => dp_n52, C1 => dp_n71, C2 
                           => dp_n344, A => dp_n378, ZN => dp_n982);
   dp_U208 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_23_port, A2 => dp_n51, 
                           B1 => dp_z_word_23_port, B2 => dp_n46, ZN => dp_n377
                           );
   dp_U207 : OAI221_X1 port map( B1 => dp_n283, B2 => dp_n52, C1 => dp_n72, C2 
                           => dp_n343, A => dp_n377, ZN => dp_n981);
   dp_U206 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_24_port, A2 => dp_n49, 
                           B1 => dp_z_word_24_port, B2 => dp_n46, ZN => dp_n376
                           );
   dp_U205 : OAI221_X1 port map( B1 => dp_n284, B2 => dp_n52, C1 => dp_n73, C2 
                           => dp_n342, A => dp_n376, ZN => dp_n980);
   dp_U204 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_25_port, A2 => dp_n49, 
                           B1 => dp_z_word_25_port, B2 => dp_n46, ZN => dp_n375
                           );
   dp_U203 : OAI221_X1 port map( B1 => dp_n285, B2 => dp_n52, C1 => dp_n71, C2 
                           => dp_n341, A => dp_n375, ZN => dp_n979);
   dp_U202 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_26_port, A2 => dp_n51, 
                           B1 => dp_z_word_26_port, B2 => dp_n46, ZN => dp_n374
                           );
   dp_U201 : OAI221_X1 port map( B1 => dp_n286, B2 => dp_n52, C1 => dp_n71, C2 
                           => dp_n340, A => dp_n374, ZN => dp_n978);
   dp_U200 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_27_port, A2 => dp_n49, 
                           B1 => dp_z_word_27_port, B2 => dp_n46, ZN => dp_n373
                           );
   dp_U199 : OAI221_X1 port map( B1 => dp_n287, B2 => dp_n52, C1 => dp_n72, C2 
                           => dp_n339, A => dp_n373, ZN => dp_n977);
   dp_U198 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_28_port, A2 => dp_n51, 
                           B1 => dp_z_word_28_port, B2 => dp_n46, ZN => dp_n372
                           );
   dp_U197 : OAI221_X1 port map( B1 => dp_n288, B2 => dp_n52, C1 => dp_n73, C2 
                           => dp_n338, A => dp_n372, ZN => dp_n976);
   dp_U196 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_29_port, A2 => dp_n49, 
                           B1 => dp_z_word_29_port, B2 => dp_n46, ZN => dp_n371
                           );
   dp_U195 : OAI221_X1 port map( B1 => dp_n289, B2 => dp_n52, C1 => dp_n71, C2 
                           => dp_n337, A => dp_n371, ZN => dp_n975);
   dp_U194 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_30_port, A2 => dp_n51, 
                           B1 => dp_z_word_30_port, B2 => dp_n46, ZN => dp_n370
                           );
   dp_U193 : OAI221_X1 port map( B1 => dp_n290, B2 => dp_n52, C1 => dp_n72, C2 
                           => dp_n336, A => dp_n370, ZN => dp_n974);
   dp_U192 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_31_port, A2 => dp_n50, 
                           B1 => dp_z_word_31_port, B2 => dp_n46, ZN => dp_n367
                           );
   dp_U191 : OAI221_X1 port map( B1 => dp_n291, B2 => dp_n52, C1 => dp_n72, C2 
                           => dp_n335, A => dp_n367, ZN => dp_n973);
   dp_U190 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_0_port, A2 => dp_n50, B1
                           => dp_z_word_0_port, B2 => dp_n48, ZN => dp_n401);
   dp_U189 : OAI221_X1 port map( B1 => dp_n260, B2 => dp_n54, C1 => dp_n73, C2 
                           => dp_n400, A => dp_n401, ZN => dp_n1004);
   dp_U188 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_1_port, A2 => dp_n50, B1
                           => dp_z_word_1_port, B2 => dp_n48, ZN => dp_n399);
   dp_U187 : OAI221_X1 port map( B1 => dp_n261, B2 => dp_n54, C1 => dp_n71, C2 
                           => dp_n365, A => dp_n399, ZN => dp_n1003);
   dp_U186 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_2_port, A2 => dp_n50, B1
                           => dp_z_word_2_port, B2 => dp_n48, ZN => dp_n398);
   dp_U185 : OAI221_X1 port map( B1 => dp_n262, B2 => dp_n54, C1 => dp_n72, C2 
                           => dp_n364, A => dp_n398, ZN => dp_n1002);
   dp_U184 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_3_port, A2 => dp_n50, B1
                           => dp_z_word_3_port, B2 => dp_n48, ZN => dp_n397);
   dp_U183 : OAI221_X1 port map( B1 => dp_n263, B2 => dp_n54, C1 => dp_n73, C2 
                           => dp_n363, A => dp_n397, ZN => dp_n1001);
   dp_U182 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_4_port, A2 => dp_n50, B1
                           => dp_z_word_4_port, B2 => dp_n48, ZN => dp_n396);
   dp_U181 : OAI221_X1 port map( B1 => dp_n264, B2 => dp_n54, C1 => dp_n71, C2 
                           => dp_n362, A => dp_n396, ZN => dp_n1000);
   dp_U180 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_5_port, A2 => dp_n50, B1
                           => dp_z_word_5_port, B2 => dp_n48, ZN => dp_n395);
   dp_U179 : OAI221_X1 port map( B1 => dp_n265, B2 => dp_n54, C1 => dp_n72, C2 
                           => dp_n361, A => dp_n395, ZN => dp_n999);
   dp_U178 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_6_port, A2 => dp_n50, B1
                           => dp_z_word_6_port, B2 => dp_n48, ZN => dp_n394);
   dp_U177 : OAI221_X1 port map( B1 => dp_n266, B2 => dp_n54, C1 => dp_n73, C2 
                           => dp_n360, A => dp_n394, ZN => dp_n998);
   dp_U176 : AOI22_X1 port map( A1 => dp_data_mem_ex_o_7_port, A2 => dp_n50, B1
                           => dp_z_word_7_port, B2 => dp_n48, ZN => dp_n393);
   dp_U175 : OAI221_X1 port map( B1 => dp_n267, B2 => dp_n54, C1 => dp_n71, C2 
                           => dp_n359, A => dp_n393, ZN => dp_n997);
   dp_U174 : OAI22_X1 port map( A1 => dp_n66, A2 => dp_n516, B1 => dp_n60, B2 
                           => dp_n293, ZN => dp_n1009);
   dp_U173 : OAI22_X1 port map( A1 => dp_n66, A2 => dp_n518, B1 => dp_n60, B2 
                           => dp_n294, ZN => dp_n1008);
   dp_U172 : OAI22_X1 port map( A1 => dp_n66, A2 => dp_n520, B1 => dp_n60, B2 
                           => dp_n295, ZN => dp_n1007);
   dp_U171 : OAI22_X1 port map( A1 => dp_n66, A2 => dp_n522, B1 => dp_n60, B2 
                           => dp_n296, ZN => dp_n1006);
   dp_U170 : OAI22_X1 port map( A1 => dp_n66, A2 => dp_n524, B1 => dp_n60, B2 
                           => dp_n297, ZN => dp_n1005);
   dp_U169 : BUF_X1 port map( A => dp_n1029, Z => dp_n24);
   dp_U168 : BUF_X1 port map( A => dp_n1029, Z => dp_n23);
   dp_U167 : BUF_X1 port map( A => dp_n122, Z => dp_n121);
   dp_U166 : BUF_X1 port map( A => dp_n122, Z => dp_n119);
   dp_U165 : BUF_X1 port map( A => dp_n122, Z => dp_n118);
   dp_U164 : BUF_X1 port map( A => dp_n122, Z => dp_n117);
   dp_U163 : BUF_X1 port map( A => dp_n122, Z => dp_n116);
   dp_U162 : BUF_X1 port map( A => dp_n122, Z => dp_n115);
   dp_U161 : BUF_X1 port map( A => dp_n122, Z => dp_n120);
   dp_U160 : AND2_X2 port map( A1 => pipe_clear_n_i, A2 => dp_n112, ZN => 
                           dp_n17);
   dp_U159 : NAND2_X1 port map( A1 => pipe_clear_n_i, A2 => dp_n131, ZN => 
                           dp_n132);
   dp_U158 : AND2_X2 port map( A1 => pipe_ex_mem_en_i, A2 => pipe_clear_n_i, ZN
                           => dp_n16);
   dp_U157 : OAI22_X1 port map( A1 => dp_n327, A2 => dp_n63, B1 => dp_n57, B2 
                           => dp_n338, ZN => dp_n945);
   dp_U156 : OAI22_X1 port map( A1 => dp_n328, A2 => dp_n63, B1 => dp_n57, B2 
                           => dp_n337, ZN => dp_n944);
   dp_U155 : OAI22_X1 port map( A1 => dp_n329, A2 => dp_n63, B1 => dp_n57, B2 
                           => dp_n336, ZN => dp_n943);
   dp_U154 : OAI22_X1 port map( A1 => dp_n330, A2 => dp_n63, B1 => dp_n57, B2 
                           => dp_n335, ZN => dp_n942);
   dp_U153 : OAI22_X1 port map( A1 => dp_n299, A2 => dp_n61, B1 => dp_n59, B2 
                           => dp_n364, ZN => dp_n971);
   dp_U152 : OAI22_X1 port map( A1 => dp_n300, A2 => dp_n61, B1 => dp_n59, B2 
                           => dp_n363, ZN => dp_n970);
   dp_U151 : OAI22_X1 port map( A1 => dp_n303, A2 => dp_n61, B1 => dp_n59, B2 
                           => dp_n362, ZN => dp_n969);
   dp_U150 : OAI22_X1 port map( A1 => dp_n304, A2 => dp_n61, B1 => dp_n59, B2 
                           => dp_n361, ZN => dp_n968);
   dp_U149 : OAI22_X1 port map( A1 => dp_n305, A2 => dp_n61, B1 => dp_n59, B2 
                           => dp_n360, ZN => dp_n967);
   dp_U148 : OAI22_X1 port map( A1 => dp_n306, A2 => dp_n61, B1 => dp_n59, B2 
                           => dp_n359, ZN => dp_n966);
   dp_U147 : OAI22_X1 port map( A1 => dp_n307, A2 => dp_n61, B1 => dp_n59, B2 
                           => dp_n358, ZN => dp_n965);
   dp_U146 : OAI22_X1 port map( A1 => dp_n308, A2 => dp_n61, B1 => dp_n59, B2 
                           => dp_n357, ZN => dp_n964);
   dp_U145 : OAI22_X1 port map( A1 => dp_n309, A2 => dp_n63, B1 => dp_n59, B2 
                           => dp_n356, ZN => dp_n963);
   dp_U144 : OAI22_X1 port map( A1 => dp_n310, A2 => dp_n62, B1 => dp_n59, B2 
                           => dp_n355, ZN => dp_n962);
   dp_U143 : OAI22_X1 port map( A1 => dp_n311, A2 => dp_n62, B1 => dp_n59, B2 
                           => dp_n354, ZN => dp_n961);
   dp_U142 : OAI22_X1 port map( A1 => dp_n312, A2 => dp_n62, B1 => dp_n59, B2 
                           => dp_n353, ZN => dp_n960);
   dp_U141 : OAI22_X1 port map( A1 => dp_n313, A2 => dp_n62, B1 => dp_n59, B2 
                           => dp_n352, ZN => dp_n959);
   dp_U140 : OAI22_X1 port map( A1 => dp_n314, A2 => dp_n62, B1 => dp_n58, B2 
                           => dp_n351, ZN => dp_n958);
   dp_U139 : OAI22_X1 port map( A1 => dp_n315, A2 => dp_n62, B1 => dp_n58, B2 
                           => dp_n350, ZN => dp_n957);
   dp_U138 : OAI22_X1 port map( A1 => dp_n316, A2 => dp_n62, B1 => dp_n58, B2 
                           => dp_n349, ZN => dp_n956);
   dp_U137 : OAI22_X1 port map( A1 => dp_n317, A2 => dp_n62, B1 => dp_n58, B2 
                           => dp_n348, ZN => dp_n955);
   dp_U136 : OAI22_X1 port map( A1 => dp_n318, A2 => dp_n62, B1 => dp_n58, B2 
                           => dp_n347, ZN => dp_n954);
   dp_U135 : OAI22_X1 port map( A1 => dp_n319, A2 => dp_n62, B1 => dp_n58, B2 
                           => dp_n346, ZN => dp_n953);
   dp_U134 : OAI22_X1 port map( A1 => dp_n320, A2 => dp_n62, B1 => dp_n58, B2 
                           => dp_n345, ZN => dp_n952);
   dp_U133 : OAI22_X1 port map( A1 => dp_n321, A2 => dp_n62, B1 => dp_n58, B2 
                           => dp_n344, ZN => dp_n951);
   dp_U132 : OAI22_X1 port map( A1 => dp_n322, A2 => dp_n63, B1 => dp_n58, B2 
                           => dp_n343, ZN => dp_n950);
   dp_U131 : OAI22_X1 port map( A1 => dp_n323, A2 => dp_n63, B1 => dp_n58, B2 
                           => dp_n342, ZN => dp_n949);
   dp_U130 : OAI22_X1 port map( A1 => dp_n324, A2 => dp_n63, B1 => dp_n58, B2 
                           => dp_n341, ZN => dp_n948);
   dp_U129 : OAI22_X1 port map( A1 => dp_n325, A2 => dp_n63, B1 => dp_n58, B2 
                           => dp_n340, ZN => dp_n947);
   dp_U128 : OAI22_X1 port map( A1 => dp_n326, A2 => dp_n63, B1 => dp_n58, B2 
                           => dp_n339, ZN => dp_n946);
   dp_U127 : CLKBUF_X1 port map( A => dp_n366, Z => dp_n54);
   dp_U126 : BUF_X1 port map( A => dp_n366, Z => dp_n52);
   dp_U125 : NOR2_X1 port map( A1 => dp_n1027, A2 => dp_n70, ZN => dp_n369);
   dp_U124 : OAI22_X1 port map( A1 => dp_n254, A2 => dp_n61, B1 => dp_n60, B2 
                           => dp_n400, ZN => dp_n1015);
   dp_U123 : OAI22_X1 port map( A1 => dp_n298, A2 => dp_n61, B1 => dp_n60, B2 
                           => dp_n365, ZN => dp_n972);
   dp_U122 : NAND2_X1 port map( A1 => pipe_clear_n_i, A2 => dp_n61, ZN => 
                           dp_n302);
   dp_U121 : BUF_X1 port map( A => dp_n23, Z => dp_n22);
   dp_U120 : BUF_X1 port map( A => dp_n24, Z => dp_n18);
   dp_U119 : BUF_X1 port map( A => dp_n23, Z => dp_n21);
   dp_U118 : BUF_X1 port map( A => dp_n23, Z => dp_n20);
   dp_U117 : OR2_X1 port map( A1 => pipe_if_id_en_i, A2 => dp_n142, ZN => 
                           dp_n131);
   dp_U116 : INV_X1 port map( A => dp_n16, ZN => dp_n70);
   dp_U115 : INV_X1 port map( A => dp_n69, ZN => dp_n103);
   dp_U114 : BUF_X1 port map( A => dp_n369, Z => dp_n48);
   dp_U113 : BUF_X1 port map( A => dp_n369, Z => dp_n47);
   dp_U112 : BUF_X1 port map( A => dp_n369, Z => dp_n46);
   dp_U111 : INV_X1 port map( A => dp_n17, ZN => dp_n71);
   dp_U110 : INV_X1 port map( A => dp_n17, ZN => dp_n72);
   dp_U109 : INV_X1 port map( A => dp_n17, ZN => dp_n73);
   dp_U108 : BUF_X1 port map( A => dp_n68, Z => dp_n106);
   dp_U107 : BUF_X1 port map( A => dp_n75, Z => dp_n85);
   dp_U106 : BUF_X1 port map( A => dp_n74, Z => dp_n77);
   dp_U105 : BUF_X1 port map( A => dp_n74, Z => dp_n78);
   dp_U104 : BUF_X1 port map( A => dp_n74, Z => dp_n79);
   dp_U103 : BUF_X1 port map( A => dp_n74, Z => dp_n80);
   dp_U102 : BUF_X1 port map( A => dp_n74, Z => dp_n76);
   dp_U101 : CLKBUF_X1 port map( A => dp_n301, Z => dp_n66);
   dp_U100 : INV_X1 port map( A => dp_n103, ZN => dp_n100);
   dp_U99 : CLKBUF_X1 port map( A => dp_n301, Z => dp_n63);
   dp_U98 : CLKBUF_X1 port map( A => dp_n301, Z => dp_n62);
   dp_U97 : CLKBUF_X1 port map( A => dp_n301, Z => dp_n64);
   dp_U96 : CLKBUF_X1 port map( A => dp_n301, Z => dp_n65);
   dp_U95 : BUF_X1 port map( A => dp_n105, Z => dp_n107);
   dp_U94 : BUF_X1 port map( A => dp_n105, Z => dp_n108);
   dp_U93 : BUF_X1 port map( A => dp_n88, Z => dp_n91);
   dp_U92 : BUF_X1 port map( A => dp_n89, Z => dp_n98);
   dp_U91 : BUF_X1 port map( A => dp_n89, Z => dp_n97);
   dp_U90 : BUF_X1 port map( A => dp_n89, Z => dp_n96);
   dp_U89 : BUF_X1 port map( A => dp_n89, Z => dp_n95);
   dp_U88 : BUF_X1 port map( A => dp_n88, Z => dp_n94);
   dp_U87 : BUF_X1 port map( A => dp_n88, Z => dp_n93);
   dp_U86 : BUF_X1 port map( A => dp_n88, Z => dp_n92);
   dp_U85 : BUF_X1 port map( A => dp_n105, Z => dp_n109);
   dp_U84 : CLKBUF_X1 port map( A => dp_n68, Z => dp_n105);
   dp_U83 : CLKBUF_X1 port map( A => dp_n131, Z => dp_n89);
   dp_U82 : BUF_X2 port map( A => dp_n301, Z => dp_n61);
   dp_U81 : CLKBUF_X1 port map( A => dp_n106, Z => dp_n111);
   dp_U80 : OAI22_X4 port map( A1 => dp_n115, A2 => dp_n331, B1 => dp_n114, B2 
                           => dp_n254, ZN => dp_wr_data_id_i_0_port);
   dp_U79 : OAI22_X4 port map( A1 => dp_n117, A2 => dp_n332, B1 => dp_n113, B2 
                           => dp_n298, ZN => dp_wr_data_id_i_1_port);
   dp_U78 : OAI22_X4 port map( A1 => dp_n119, A2 => dp_n333, B1 => dp_n113, B2 
                           => dp_n299, ZN => dp_wr_data_id_i_2_port);
   dp_U77 : OAI22_X4 port map( A1 => dp_n120, A2 => dp_n334, B1 => dp_n113, B2 
                           => dp_n300, ZN => dp_wr_data_id_i_3_port);
   dp_U76 : OAI22_X4 port map( A1 => dp_n115, A2 => dp_n408, B1 => dp_n114, B2 
                           => dp_n309, ZN => dp_wr_data_id_i_10_port);
   dp_U75 : OAI22_X4 port map( A1 => dp_n116, A2 => dp_n519, B1 => wb_mux_sel_i
                           , B2 => dp_n316, ZN => dp_wr_data_id_i_17_port);
   dp_U74 : OAI22_X4 port map( A1 => dp_n120, A2 => dp_n402, B1 => dp_n113, B2 
                           => dp_n303, ZN => dp_wr_data_id_i_4_port);
   dp_U73 : OAI22_X4 port map( A1 => dp_n115, A2 => dp_n409, B1 => dp_n114, B2 
                           => dp_n310, ZN => dp_wr_data_id_i_11_port);
   dp_U72 : OAI22_X4 port map( A1 => dp_n116, A2 => dp_n521, B1 => wb_mux_sel_i
                           , B2 => dp_n317, ZN => dp_wr_data_id_i_18_port);
   dp_U71 : OAI22_X4 port map( A1 => dp_n120, A2 => dp_n403, B1 => dp_n113, B2 
                           => dp_n304, ZN => dp_wr_data_id_i_5_port);
   dp_U70 : OAI22_X4 port map( A1 => dp_n115, A2 => dp_n410, B1 => dp_n114, B2 
                           => dp_n311, ZN => dp_wr_data_id_i_12_port);
   dp_U69 : OAI22_X4 port map( A1 => dp_n117, A2 => dp_n523, B1 => dp_n113, B2 
                           => dp_n318, ZN => dp_wr_data_id_i_19_port);
   dp_U68 : OAI22_X4 port map( A1 => dp_n120, A2 => dp_n404, B1 => dp_n113, B2 
                           => dp_n305, ZN => dp_wr_data_id_i_6_port);
   dp_U67 : OAI22_X4 port map( A1 => dp_n115, A2 => dp_n411, B1 => dp_n114, B2 
                           => dp_n312, ZN => dp_wr_data_id_i_13_port);
   dp_U66 : OAI22_X4 port map( A1 => dp_n117, A2 => dp_n525, B1 => dp_n113, B2 
                           => dp_n319, ZN => dp_wr_data_id_i_20_port);
   dp_U65 : INV_X2 port map( A => dp_n121, ZN => dp_n113);
   dp_U64 : OAI22_X4 port map( A1 => dp_n120, A2 => dp_n405, B1 => dp_n113, B2 
                           => dp_n306, ZN => dp_wr_data_id_i_7_port);
   dp_U63 : OAI22_X4 port map( A1 => dp_n121, A2 => dp_n406, B1 => dp_n113, B2 
                           => dp_n307, ZN => dp_wr_data_id_i_8_port);
   dp_U62 : OAI22_X4 port map( A1 => dp_n116, A2 => dp_n412, B1 => dp_n114, B2 
                           => dp_n313, ZN => dp_wr_data_id_i_14_port);
   dp_U61 : OAI22_X4 port map( A1 => dp_n117, A2 => dp_n584, B1 => wb_mux_sel_i
                           , B2 => dp_n320, ZN => dp_wr_data_id_i_21_port);
   dp_U60 : OAI22_X4 port map( A1 => dp_n118, A2 => dp_n586, B1 => wb_mux_sel_i
                           , B2 => dp_n322, ZN => dp_wr_data_id_i_23_port);
   dp_U59 : OAI22_X4 port map( A1 => dp_n121, A2 => dp_n407, B1 => dp_n113, B2 
                           => dp_n308, ZN => dp_wr_data_id_i_9_port);
   dp_U58 : OAI22_X4 port map( A1 => dp_n116, A2 => dp_n413, B1 => dp_n114, B2 
                           => dp_n314, ZN => dp_wr_data_id_i_15_port);
   dp_U57 : OAI22_X4 port map( A1 => dp_n117, A2 => dp_n585, B1 => dp_n113, B2 
                           => dp_n321, ZN => dp_wr_data_id_i_22_port);
   dp_U56 : OAI22_X4 port map( A1 => dp_n116, A2 => dp_n517, B1 => dp_n114, B2 
                           => dp_n315, ZN => dp_wr_data_id_i_16_port);
   dp_U55 : OAI22_X4 port map( A1 => dp_n118, A2 => dp_n587, B1 => wb_mux_sel_i
                           , B2 => dp_n323, ZN => dp_wr_data_id_i_24_port);
   dp_U54 : OAI22_X4 port map( A1 => dp_n119, A2 => dp_n591, B1 => dp_n113, B2 
                           => dp_n327, ZN => dp_wr_data_id_i_28_port);
   dp_U53 : OAI22_X4 port map( A1 => dp_n118, A2 => dp_n588, B1 => wb_mux_sel_i
                           , B2 => dp_n324, ZN => dp_wr_data_id_i_25_port);
   dp_U52 : OAI22_X4 port map( A1 => dp_n119, A2 => dp_n592, B1 => dp_n113, B2 
                           => dp_n328, ZN => dp_wr_data_id_i_29_port);
   dp_U51 : BUF_X2 port map( A => dp_n368, Z => dp_n49);
   dp_U50 : BUF_X2 port map( A => dp_n368, Z => dp_n50);
   dp_U49 : BUF_X2 port map( A => dp_n88, Z => dp_n90);
   dp_U48 : BUF_X2 port map( A => dp_n132, Z => dp_n75);
   dp_U47 : BUF_X2 port map( A => dp_n75, Z => dp_n84);
   dp_U46 : BUF_X2 port map( A => dp_n368, Z => dp_n51);
   dp_U45 : OR2_X1 port map( A1 => pipe_if_id_en_i, A2 => dp_n142, ZN => 
                           dp_n301);
   dp_U44 : INV_X4 port map( A => dp_n16, ZN => dp_n67);
   dp_U43 : BUF_X2 port map( A => dp_n366, Z => dp_n53);
   dp_U42 : INV_X1 port map( A => dp_n67, ZN => dp_n15);
   dp_U41 : NAND3_X1 port map( A1 => dp_n13, A2 => dp_n14, A3 => dp_n381, ZN =>
                           dp_n985);
   dp_U40 : OR2_X1 port map( A1 => dp_n72, A2 => dp_n347, ZN => dp_n14);
   dp_U39 : OR2_X1 port map( A1 => dp_n279, A2 => dp_n53, ZN => dp_n13);
   dp_U38 : BUF_X2 port map( A => dp_n75, Z => dp_n87);
   dp_U37 : BUF_X1 port map( A => dp_n131, Z => dp_n88);
   dp_U36 : INV_X8 port map( A => RST, ZN => dp_n1029);
   dp_U35 : OAI22_X1 port map( A1 => dp_n119, A2 => dp_n1025, B1 => dp_n113, B2
                           => dp_n330, ZN => dp_wr_data_id_i_31_port);
   dp_U34 : INV_X1 port map( A => dp_wr_data_id_i_31_port, ZN => dp_n11);
   dp_U33 : OAI22_X1 port map( A1 => dp_n119, A2 => dp_n593, B1 => dp_n113, B2 
                           => dp_n329, ZN => dp_wr_data_id_i_30_port);
   dp_U32 : INV_X1 port map( A => dp_wr_data_id_i_30_port, ZN => dp_n9);
   dp_U31 : OAI22_X1 port map( A1 => dp_n118, A2 => dp_n590, B1 => dp_n113, B2 
                           => dp_n326, ZN => dp_wr_data_id_i_27_port);
   dp_U30 : INV_X1 port map( A => dp_wr_data_id_i_27_port, ZN => dp_n7);
   dp_U29 : OAI22_X1 port map( A1 => dp_n118, A2 => dp_n589, B1 => dp_n113, B2 
                           => dp_n325, ZN => dp_wr_data_id_i_26_port);
   dp_U28 : INV_X1 port map( A => dp_wr_data_id_i_26_port, ZN => dp_n5);
   dp_U27 : CLKBUF_X1 port map( A => dp_n24, Z => dp_n19);
   dp_U26 : INV_X1 port map( A => dp_n103, ZN => dp_n101);
   dp_U25 : INV_X1 port map( A => dp_n103, ZN => dp_n4);
   dp_U24 : INV_X1 port map( A => dp_n103, ZN => dp_n3);
   dp_U23 : NAND2_X2 port map( A1 => dp_n106, A2 => pipe_clear_n_i, ZN => 
                           dp_n69);
   dp_U22 : INV_X2 port map( A => dp_n69, ZN => dp_n104);
   dp_U21 : BUF_X2 port map( A => dp_n302, Z => dp_n60);
   dp_U20 : BUF_X2 port map( A => dp_n302, Z => dp_n58);
   dp_U19 : BUF_X2 port map( A => dp_n302, Z => dp_n59);
   dp_U18 : BUF_X2 port map( A => dp_n302, Z => dp_n57);
   dp_U17 : BUF_X2 port map( A => dp_n302, Z => dp_n56);
   dp_U16 : BUF_X2 port map( A => dp_n302, Z => dp_n55);
   dp_U15 : BUF_X2 port map( A => dp_n74, Z => dp_n81);
   dp_U14 : BUF_X2 port map( A => dp_n75, Z => dp_n83);
   dp_U13 : BUF_X2 port map( A => dp_n75, Z => dp_n82);
   dp_U12 : BUF_X2 port map( A => dp_n75, Z => dp_n86);
   dp_U11 : BUF_X2 port map( A => dp_n106, Z => dp_n110);
   dp_U10 : INV_X1 port map( A => dp_n11, ZN => dp_n12);
   dp_U9 : INV_X1 port map( A => dp_n9, ZN => dp_n10);
   dp_U8 : INV_X1 port map( A => dp_n7, ZN => dp_n8);
   dp_U7 : INV_X1 port map( A => dp_n5, ZN => dp_n6);
   dp_U6 : BUF_X1 port map( A => dp_n132, Z => dp_n74);
   dp_npc_id_i_reg_16_inst : DFFR_X2 port map( D => dp_n691, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_16_port, QN => dp_n558);
   dp_npc_id_i_reg_17_inst : DFFR_X2 port map( D => dp_n692, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_17_port, QN => dp_n559);
   dp_npc_id_i_reg_18_inst : DFFR_X2 port map( D => dp_n693, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_18_port, QN => dp_n560);
   dp_npc_id_i_reg_19_inst : DFFR_X2 port map( D => dp_n694, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_19_port, QN => dp_n561);
   dp_npc_id_i_reg_20_inst : DFFR_X2 port map( D => dp_n695, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_20_port, QN => dp_n562);
   dp_npc_id_i_reg_21_inst : DFFR_X2 port map( D => dp_n696, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_21_port, QN => dp_n563);
   dp_npc_id_i_reg_22_inst : DFFR_X2 port map( D => dp_n697, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_22_port, QN => dp_n564);
   dp_npc_id_i_reg_23_inst : DFFR_X2 port map( D => dp_n698, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_23_port, QN => dp_n565);
   dp_npc_id_i_reg_24_inst : DFFR_X2 port map( D => dp_n699, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_24_port, QN => dp_n566);
   dp_npc_id_i_reg_26_inst : DFFR_X2 port map( D => dp_n701, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_26_port, QN => dp_n568);
   dp_npc_id_i_reg_27_inst : DFFR_X2 port map( D => dp_n702, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_27_port, QN => dp_n569);
   dp_npc_id_i_reg_25_inst : DFFR_X2 port map( D => dp_n700, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_25_port, QN => dp_n567);
   dp_npc_id_i_reg_28_inst : DFFR_X2 port map( D => dp_n703, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_28_port, QN => dp_n570);
   dp_npc_id_i_reg_29_inst : DFFR_X2 port map( D => dp_n704, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_29_port, QN => dp_n571);
   dp_npc_id_i_reg_30_inst : DFFR_X2 port map( D => dp_n705, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_30_port, QN => dp_n572);
   dp_data_mem_mem_i_reg_20_inst : DFFR_X1 port map( D => dp_n984, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(20), QN => n_1039);
   dp_data_mem_mem_i_reg_21_inst : DFFR_X1 port map( D => dp_n983, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(21), QN => n_1040);
   dp_data_mem_mem_i_reg_22_inst : DFFR_X1 port map( D => dp_n982, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(22), QN => n_1041);
   dp_data_mem_mem_i_reg_23_inst : DFFR_X1 port map( D => dp_n981, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(23), QN => n_1042);
   dp_data_mem_mem_i_reg_24_inst : DFFR_X1 port map( D => dp_n980, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(24), QN => n_1043);
   dp_data_mem_mem_i_reg_25_inst : DFFR_X1 port map( D => dp_n979, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(25), QN => n_1044);
   dp_data_mem_mem_i_reg_26_inst : DFFR_X1 port map( D => dp_n978, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(26), QN => n_1045);
   dp_data_mem_mem_i_reg_27_inst : DFFR_X1 port map( D => dp_n977, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(27), QN => n_1046);
   dp_data_mem_mem_i_reg_28_inst : DFFR_X1 port map( D => dp_n976, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(28), QN => n_1047);
   dp_data_mem_mem_i_reg_29_inst : DFFR_X1 port map( D => dp_n975, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(29), QN => n_1048);
   dp_data_mem_mem_i_reg_30_inst : DFFR_X1 port map( D => dp_n974, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(30), QN => n_1049);
   dp_data_mem_mem_i_reg_31_inst : DFFR_X1 port map( D => dp_n973, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(31), QN => n_1050);
   dp_data_mem_mem_i_reg_8_inst : DFFR_X1 port map( D => dp_n996, CK => CLK, RN
                           => dp_n1029, Q => DRAM_DATA(8), QN => n_1051);
   dp_data_mem_mem_i_reg_9_inst : DFFR_X1 port map( D => dp_n995, CK => CLK, RN
                           => dp_n1029, Q => DRAM_DATA(9), QN => n_1052);
   dp_data_mem_mem_i_reg_10_inst : DFFR_X1 port map( D => dp_n994, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(10), QN => n_1053);
   dp_data_mem_mem_i_reg_11_inst : DFFR_X1 port map( D => dp_n993, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(11), QN => n_1054);
   dp_data_mem_mem_i_reg_12_inst : DFFR_X1 port map( D => dp_n992, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(12), QN => n_1055);
   dp_data_mem_mem_i_reg_13_inst : DFFR_X1 port map( D => dp_n991, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(13), QN => n_1056);
   dp_data_mem_mem_i_reg_14_inst : DFFR_X1 port map( D => dp_n990, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(14), QN => n_1057);
   dp_data_mem_mem_i_reg_15_inst : DFFR_X1 port map( D => dp_n989, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(15), QN => n_1058);
   dp_data_mem_mem_i_reg_16_inst : DFFR_X1 port map( D => dp_n988, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(16), QN => n_1059);
   dp_data_mem_mem_i_reg_17_inst : DFFR_X1 port map( D => dp_n987, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(17), QN => n_1060);
   dp_data_mem_mem_i_reg_18_inst : DFFR_X1 port map( D => dp_n986, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(18), QN => n_1061);
   dp_data_mem_mem_i_reg_0_inst : DFFR_X1 port map( D => dp_n1004, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(0), QN => n_1062);
   dp_data_mem_mem_i_reg_1_inst : DFFR_X1 port map( D => dp_n1003, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(1), QN => n_1063);
   dp_data_mem_mem_i_reg_2_inst : DFFR_X1 port map( D => dp_n1002, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(2), QN => n_1064);
   dp_data_mem_mem_i_reg_3_inst : DFFR_X1 port map( D => dp_n1001, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(3), QN => n_1065);
   dp_data_mem_mem_i_reg_4_inst : DFFR_X1 port map( D => dp_n1000, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(4), QN => n_1066);
   dp_data_mem_mem_i_reg_5_inst : DFFR_X1 port map( D => dp_n999, CK => CLK, RN
                           => dp_n1029, Q => DRAM_DATA(5), QN => n_1067);
   dp_data_mem_mem_i_reg_6_inst : DFFR_X1 port map( D => dp_n998, CK => CLK, RN
                           => dp_n1029, Q => DRAM_DATA(6), QN => n_1068);
   dp_data_mem_mem_i_reg_7_inst : DFFR_X1 port map( D => dp_n997, CK => CLK, RN
                           => dp_n1029, Q => DRAM_DATA(7), QN => n_1069);
   dp_data_mem_wb_i_reg_10_inst : DFFR_X1 port map( D => dp_n963, CK => CLK, RN
                           => dp_n1029, Q => n_1070, QN => dp_n309);
   dp_data_mem_wb_i_reg_11_inst : DFFR_X1 port map( D => dp_n962, CK => CLK, RN
                           => dp_n1029, Q => n_1071, QN => dp_n310);
   dp_data_mem_wb_i_reg_12_inst : DFFR_X1 port map( D => dp_n961, CK => CLK, RN
                           => dp_n1029, Q => n_1072, QN => dp_n311);
   dp_data_mem_wb_i_reg_13_inst : DFFR_X1 port map( D => dp_n960, CK => CLK, RN
                           => dp_n1029, Q => n_1073, QN => dp_n312);
   dp_data_mem_wb_i_reg_14_inst : DFFR_X1 port map( D => dp_n959, CK => CLK, RN
                           => dp_n1029, Q => n_1074, QN => dp_n313);
   dp_data_mem_wb_i_reg_15_inst : DFFR_X1 port map( D => dp_n958, CK => CLK, RN
                           => dp_n1029, Q => n_1075, QN => dp_n314);
   dp_data_mem_wb_i_reg_16_inst : DFFR_X1 port map( D => dp_n957, CK => CLK, RN
                           => dp_n1029, Q => n_1076, QN => dp_n315);
   dp_data_mem_wb_i_reg_17_inst : DFFR_X1 port map( D => dp_n956, CK => CLK, RN
                           => dp_n1029, Q => n_1077, QN => dp_n316);
   dp_data_mem_wb_i_reg_18_inst : DFFR_X1 port map( D => dp_n955, CK => CLK, RN
                           => dp_n1029, Q => n_1078, QN => dp_n317);
   dp_data_mem_wb_i_reg_19_inst : DFFR_X1 port map( D => dp_n954, CK => CLK, RN
                           => dp_n1029, Q => n_1079, QN => dp_n318);
   dp_data_mem_wb_i_reg_20_inst : DFFR_X1 port map( D => dp_n953, CK => CLK, RN
                           => dp_n1029, Q => n_1080, QN => dp_n319);
   dp_data_mem_wb_i_reg_21_inst : DFFR_X1 port map( D => dp_n952, CK => CLK, RN
                           => dp_n1029, Q => n_1081, QN => dp_n320);
   dp_data_mem_wb_i_reg_22_inst : DFFR_X1 port map( D => dp_n951, CK => CLK, RN
                           => dp_n1029, Q => n_1082, QN => dp_n321);
   dp_data_mem_wb_i_reg_23_inst : DFFR_X1 port map( D => dp_n950, CK => CLK, RN
                           => dp_n1029, Q => n_1083, QN => dp_n322);
   dp_data_mem_wb_i_reg_24_inst : DFFR_X1 port map( D => dp_n949, CK => CLK, RN
                           => dp_n1029, Q => n_1084, QN => dp_n323);
   dp_data_mem_wb_i_reg_25_inst : DFFR_X1 port map( D => dp_n948, CK => CLK, RN
                           => dp_n1029, Q => n_1085, QN => dp_n324);
   dp_data_mem_wb_i_reg_26_inst : DFFR_X1 port map( D => dp_n947, CK => CLK, RN
                           => dp_n1029, Q => n_1086, QN => dp_n325);
   dp_data_mem_wb_i_reg_27_inst : DFFR_X1 port map( D => dp_n946, CK => CLK, RN
                           => dp_n1029, Q => n_1087, QN => dp_n326);
   dp_data_mem_mem_i_reg_19_inst : DFFR_X1 port map( D => dp_n985, CK => CLK, 
                           RN => dp_n1029, Q => DRAM_DATA(19), QN => n_1088);
   dp_data_mem_wb_i_reg_2_inst : DFFR_X1 port map( D => dp_n971, CK => CLK, RN 
                           => dp_n1029, Q => n_1089, QN => dp_n299);
   dp_data_mem_wb_i_reg_3_inst : DFFR_X1 port map( D => dp_n970, CK => CLK, RN 
                           => dp_n1029, Q => n_1090, QN => dp_n300);
   dp_data_mem_wb_i_reg_4_inst : DFFR_X1 port map( D => dp_n969, CK => CLK, RN 
                           => dp_n1029, Q => n_1091, QN => dp_n303);
   dp_data_mem_wb_i_reg_5_inst : DFFR_X1 port map( D => dp_n968, CK => CLK, RN 
                           => dp_n1029, Q => n_1092, QN => dp_n304);
   dp_data_mem_wb_i_reg_6_inst : DFFR_X1 port map( D => dp_n967, CK => CLK, RN 
                           => dp_n1029, Q => n_1093, QN => dp_n305);
   dp_data_mem_wb_i_reg_7_inst : DFFR_X1 port map( D => dp_n966, CK => CLK, RN 
                           => dp_n1029, Q => n_1094, QN => dp_n306);
   dp_data_mem_wb_i_reg_8_inst : DFFR_X1 port map( D => dp_n965, CK => CLK, RN 
                           => dp_n1029, Q => n_1095, QN => dp_n307);
   dp_data_mem_wb_i_reg_9_inst : DFFR_X1 port map( D => dp_n964, CK => CLK, RN 
                           => dp_n1029, Q => n_1096, QN => dp_n308);
   dp_alu_out_wb_i_reg_0_inst : DFFR_X1 port map( D => dp_n909, CK => CLK, RN 
                           => dp_n1029, Q => n_1097, QN => dp_n331);
   dp_alu_out_wb_i_reg_1_inst : DFFR_X1 port map( D => dp_n908, CK => CLK, RN 
                           => dp_n1029, Q => n_1098, QN => dp_n332);
   dp_alu_out_wb_i_reg_2_inst : DFFR_X1 port map( D => dp_n907, CK => CLK, RN 
                           => dp_n1029, Q => n_1099, QN => dp_n333);
   dp_alu_out_wb_i_reg_3_inst : DFFR_X1 port map( D => dp_n906, CK => CLK, RN 
                           => dp_n1029, Q => n_1100, QN => dp_n334);
   dp_alu_out_wb_i_reg_4_inst : DFFR_X1 port map( D => dp_n905, CK => CLK, RN 
                           => dp_n1029, Q => n_1101, QN => dp_n402);
   dp_alu_out_wb_i_reg_5_inst : DFFR_X1 port map( D => dp_n904, CK => CLK, RN 
                           => dp_n1029, Q => n_1102, QN => dp_n403);
   dp_alu_out_wb_i_reg_6_inst : DFFR_X1 port map( D => dp_n903, CK => CLK, RN 
                           => dp_n1029, Q => n_1103, QN => dp_n404);
   dp_alu_out_wb_i_reg_7_inst : DFFR_X1 port map( D => dp_n902, CK => CLK, RN 
                           => dp_n1029, Q => n_1104, QN => dp_n405);
   dp_alu_out_wb_i_reg_8_inst : DFFR_X1 port map( D => dp_n901, CK => CLK, RN 
                           => dp_n1029, Q => n_1105, QN => dp_n406);
   dp_alu_out_wb_i_reg_9_inst : DFFR_X1 port map( D => dp_n900, CK => CLK, RN 
                           => dp_n1029, Q => n_1106, QN => dp_n407);
   dp_alu_out_wb_i_reg_10_inst : DFFR_X1 port map( D => dp_n899, CK => CLK, RN 
                           => dp_n1029, Q => n_1107, QN => dp_n408);
   dp_alu_out_wb_i_reg_11_inst : DFFR_X1 port map( D => dp_n898, CK => CLK, RN 
                           => dp_n1029, Q => n_1108, QN => dp_n409);
   dp_alu_out_wb_i_reg_12_inst : DFFR_X1 port map( D => dp_n897, CK => CLK, RN 
                           => dp_n1029, Q => n_1109, QN => dp_n410);
   dp_alu_out_wb_i_reg_13_inst : DFFR_X1 port map( D => dp_n896, CK => CLK, RN 
                           => dp_n1029, Q => n_1110, QN => dp_n411);
   dp_alu_out_wb_i_reg_14_inst : DFFR_X1 port map( D => dp_n895, CK => CLK, RN 
                           => dp_n1029, Q => n_1111, QN => dp_n412);
   dp_alu_out_wb_i_reg_15_inst : DFFR_X1 port map( D => dp_n894, CK => CLK, RN 
                           => dp_n1029, Q => n_1112, QN => dp_n413);
   dp_alu_out_wb_i_reg_16_inst : DFFR_X1 port map( D => dp_n893, CK => CLK, RN 
                           => dp_n1029, Q => n_1113, QN => dp_n517);
   dp_alu_out_wb_i_reg_17_inst : DFFR_X1 port map( D => dp_n892, CK => CLK, RN 
                           => dp_n1029, Q => n_1114, QN => dp_n519);
   dp_alu_out_wb_i_reg_18_inst : DFFR_X1 port map( D => dp_n891, CK => CLK, RN 
                           => dp_n1029, Q => n_1115, QN => dp_n521);
   dp_alu_out_wb_i_reg_19_inst : DFFR_X1 port map( D => dp_n890, CK => CLK, RN 
                           => dp_n1029, Q => n_1116, QN => dp_n523);
   dp_alu_out_wb_i_reg_20_inst : DFFR_X1 port map( D => dp_n889, CK => CLK, RN 
                           => dp_n1029, Q => n_1117, QN => dp_n525);
   dp_alu_out_wb_i_reg_21_inst : DFFR_X1 port map( D => dp_n888, CK => CLK, RN 
                           => dp_n1029, Q => n_1118, QN => dp_n584);
   dp_alu_out_wb_i_reg_22_inst : DFFR_X1 port map( D => dp_n887, CK => CLK, RN 
                           => dp_n1029, Q => n_1119, QN => dp_n585);
   dp_alu_out_wb_i_reg_23_inst : DFFR_X1 port map( D => dp_n886, CK => CLK, RN 
                           => dp_n1029, Q => n_1120, QN => dp_n586);
   dp_alu_out_wb_i_reg_24_inst : DFFR_X1 port map( D => dp_n885, CK => CLK, RN 
                           => dp_n1029, Q => n_1121, QN => dp_n587);
   dp_alu_out_wb_i_reg_25_inst : DFFR_X1 port map( D => dp_n884, CK => CLK, RN 
                           => dp_n1029, Q => n_1122, QN => dp_n588);
   dp_alu_out_wb_i_reg_26_inst : DFFR_X1 port map( D => dp_n883, CK => CLK, RN 
                           => dp_n1029, Q => n_1123, QN => dp_n589);
   dp_alu_out_wb_i_reg_27_inst : DFFR_X1 port map( D => dp_n882, CK => CLK, RN 
                           => dp_n1029, Q => n_1124, QN => dp_n590);
   dp_alu_out_wb_i_reg_28_inst : DFFR_X1 port map( D => dp_n881, CK => CLK, RN 
                           => dp_n1029, Q => n_1125, QN => dp_n591);
   dp_alu_out_wb_i_reg_29_inst : DFFR_X1 port map( D => dp_n880, CK => CLK, RN 
                           => dp_n1029, Q => n_1126, QN => dp_n592);
   dp_alu_out_wb_i_reg_30_inst : DFFR_X1 port map( D => dp_n879, CK => CLK, RN 
                           => dp_n1029, Q => n_1127, QN => dp_n593);
   dp_alu_out_wb_i_reg_31_inst : DFFR_X1 port map( D => dp_n878, CK => CLK, RN 
                           => dp_n1029, Q => n_1128, QN => dp_n1025);
   dp_data_mem_wb_i_reg_28_inst : DFFR_X1 port map( D => dp_n945, CK => CLK, RN
                           => dp_n1029, Q => n_1129, QN => dp_n327);
   dp_data_mem_wb_i_reg_29_inst : DFFR_X1 port map( D => dp_n944, CK => CLK, RN
                           => dp_n1029, Q => n_1130, QN => dp_n328);
   dp_data_mem_wb_i_reg_30_inst : DFFR_X1 port map( D => dp_n943, CK => CLK, RN
                           => dp_n1029, Q => n_1131, QN => dp_n329);
   dp_data_mem_wb_i_reg_31_inst : DFFR_X1 port map( D => dp_n942, CK => CLK, RN
                           => dp_n1029, Q => n_1132, QN => dp_n330);
   dp_data_mem_wb_i_reg_0_inst : DFFR_X1 port map( D => dp_n1015, CK => CLK, RN
                           => dp_n1029, Q => n_1133, QN => dp_n254);
   dp_data_mem_wb_i_reg_1_inst : DFFR_X1 port map( D => dp_n972, CK => CLK, RN 
                           => dp_n1029, Q => n_1134, QN => dp_n298);
   dp_npc_ex_i_reg_3_inst : DFFR_X1 port map( D => dp_n720, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_3_port, QN => dp_n263);
   dp_npc_ex_i_reg_4_inst : DFFR_X1 port map( D => dp_n721, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_4_port, QN => dp_n264);
   dp_npc_ex_i_reg_6_inst : DFFR_X1 port map( D => dp_n723, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_6_port, QN => dp_n266);
   dp_npc_ex_i_reg_11_inst : DFFR_X1 port map( D => dp_n728, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_11_port, QN => dp_n271);
   dp_npc_ex_i_reg_18_inst : DFFR_X1 port map( D => dp_n735, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_18_port, QN => dp_n278);
   dp_npc_ex_i_reg_19_inst : DFFR_X1 port map( D => dp_n736, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_19_port, QN => dp_n279);
   dp_npc_ex_i_reg_20_inst : DFFR_X1 port map( D => dp_n737, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_20_port, QN => dp_n280);
   dp_npc_ex_i_reg_24_inst : DFFR_X1 port map( D => dp_n741, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_24_port, QN => dp_n284);
   dp_npc_ex_i_reg_26_inst : DFFR_X1 port map( D => dp_n743, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_26_port, QN => dp_n286);
   dp_npc_ex_i_reg_5_inst : DFFR_X1 port map( D => dp_n722, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_5_port, QN => dp_n265);
   dp_npc_ex_i_reg_7_inst : DFFR_X1 port map( D => dp_n724, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_7_port, QN => dp_n267);
   dp_npc_ex_i_reg_8_inst : DFFR_X1 port map( D => dp_n725, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_8_port, QN => dp_n268);
   dp_npc_ex_i_reg_9_inst : DFFR_X1 port map( D => dp_n726, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_9_port, QN => dp_n269);
   dp_npc_ex_i_reg_10_inst : DFFR_X1 port map( D => dp_n727, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_10_port, QN => dp_n270);
   dp_npc_ex_i_reg_12_inst : DFFR_X1 port map( D => dp_n729, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_12_port, QN => dp_n272);
   dp_npc_ex_i_reg_13_inst : DFFR_X1 port map( D => dp_n730, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_13_port, QN => dp_n273);
   dp_npc_ex_i_reg_14_inst : DFFR_X1 port map( D => dp_n731, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_14_port, QN => dp_n274);
   dp_npc_ex_i_reg_15_inst : DFFR_X1 port map( D => dp_n732, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_15_port, QN => dp_n275);
   dp_npc_ex_i_reg_16_inst : DFFR_X1 port map( D => dp_n733, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_16_port, QN => dp_n276);
   dp_npc_ex_i_reg_17_inst : DFFR_X1 port map( D => dp_n734, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_17_port, QN => dp_n277);
   dp_npc_ex_i_reg_21_inst : DFFR_X1 port map( D => dp_n738, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_21_port, QN => dp_n281);
   dp_npc_ex_i_reg_22_inst : DFFR_X1 port map( D => dp_n739, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_22_port, QN => dp_n282);
   dp_npc_ex_i_reg_23_inst : DFFR_X1 port map( D => dp_n740, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_23_port, QN => dp_n283);
   dp_npc_ex_i_reg_25_inst : DFFR_X1 port map( D => dp_n742, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_25_port, QN => dp_n285);
   dp_npc_ex_i_reg_27_inst : DFFR_X1 port map( D => dp_n744, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_27_port, QN => dp_n287);
   dp_npc_ex_i_reg_28_inst : DFFR_X1 port map( D => dp_n745, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_28_port, QN => dp_n288);
   dp_npc_ex_i_reg_29_inst : DFFR_X1 port map( D => dp_n746, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_29_port, QN => dp_n289);
   dp_npc_ex_i_reg_30_inst : DFFR_X1 port map( D => dp_n747, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_30_port, QN => dp_n290);
   dp_npc_ex_i_reg_31_inst : DFFR_X1 port map( D => dp_n748, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_31_port, QN => dp_n291);
   dp_npc_ex_i_reg_0_inst : DFFR_X1 port map( D => dp_n717, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_0_port, QN => dp_n260);
   dp_npc_ex_i_reg_1_inst : DFFR_X1 port map( D => dp_n718, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_1_port, QN => dp_n261);
   dp_npc_ex_i_reg_2_inst : DFFR_X1 port map( D => dp_n719, CK => CLK, RN => 
                           dp_n1029, Q => dp_npc_ex_i_2_port, QN => dp_n262);
   dp_rd_fwd_mem_i_reg_0_inst : DFFR_X1 port map( D => dp_n1014, CK => CLK, RN 
                           => dp_n1029, Q => n_1135, QN => dp_n293);
   dp_rd_fwd_mem_i_reg_1_inst : DFFR_X1 port map( D => dp_n1013, CK => CLK, RN 
                           => dp_n1029, Q => n_1136, QN => dp_n294);
   dp_rd_fwd_mem_i_reg_2_inst : DFFR_X1 port map( D => dp_n1012, CK => CLK, RN 
                           => dp_n1029, Q => n_1137, QN => dp_n295);
   dp_rd_fwd_mem_i_reg_4_inst : DFFR_X1 port map( D => dp_n1010, CK => CLK, RN 
                           => dp_n1029, Q => n_1138, QN => dp_n297);
   dp_rd_fwd_mem_i_reg_3_inst : DFFR_X1 port map( D => dp_n1011, CK => CLK, RN 
                           => dp_n1029, Q => n_1139, QN => dp_n296);
   dp_z_word_tri_31_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_31_port);
   dp_z_word_tri_30_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_30_port);
   dp_z_word_tri_29_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_29_port);
   dp_z_word_tri_28_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_28_port);
   dp_z_word_tri_27_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_27_port);
   dp_z_word_tri_26_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_26_port);
   dp_z_word_tri_25_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_25_port);
   dp_z_word_tri_24_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_24_port);
   dp_z_word_tri_23_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_23_port);
   dp_z_word_tri_22_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_22_port);
   dp_z_word_tri_21_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_21_port);
   dp_z_word_tri_20_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_20_port);
   dp_z_word_tri_19_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_19_port);
   dp_z_word_tri_18_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_18_port);
   dp_z_word_tri_17_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_17_port);
   dp_z_word_tri_16_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_16_port);
   dp_z_word_tri_15_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_15_port);
   dp_z_word_tri_14_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_14_port);
   dp_z_word_tri_13_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_13_port);
   dp_z_word_tri_12_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_12_port);
   dp_z_word_tri_11_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_11_port);
   dp_z_word_tri_10_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_10_port);
   dp_z_word_tri_9_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_9_port);
   dp_z_word_tri_8_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_8_port);
   dp_z_word_tri_7_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_7_port);
   dp_z_word_tri_6_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_6_port);
   dp_z_word_tri_5_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_5_port);
   dp_z_word_tri_4_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_4_port);
   dp_z_word_tri_3_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_3_port);
   dp_z_word_tri_2_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_2_port);
   dp_z_word_tri_1_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_1_port);
   dp_z_word_tri_0_inst : TBUF_X1 port map( A => dp_n1, EN => dp_n2, Z => 
                           dp_z_word_0_port);
   dp_U752 : NOR3_X2 port map( A1 => mem_in_en_i, A2 => npc_wb_en_i, A3 => 
                           dp_n70, ZN => dp_n368);
   dp_U753 : NAND3_X1 port map( A1 => dp_n16, A2 => dp_n1027, A3 => npc_wb_en_i
                           , ZN => dp_n366);
   dp_n1 <= '0';
   dp_n2 <= '1';
   dp_npc_id_i_reg_31_inst : DFFR_X1 port map( D => dp_n706, CK => CLK, RN => 
                           dp_n25, Q => dp_npc_id_o_31_port, QN => dp_n573);
   dp_npc_id_i_reg_15_inst : DFFR_X1 port map( D => dp_n690, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_15_port, QN => dp_n557);
   dp_npc_id_i_reg_14_inst : DFFR_X1 port map( D => dp_n689, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_14_port, QN => dp_n556);
   dp_npc_id_i_reg_13_inst : DFFR_X1 port map( D => dp_n688, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_13_port, QN => dp_n555);
   dp_npc_id_i_reg_12_inst : DFFR_X1 port map( D => dp_n687, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_12_port, QN => dp_n554);
   dp_npc_id_i_reg_11_inst : DFFR_X1 port map( D => dp_n686, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_11_port, QN => dp_n553);
   dp_npc_id_i_reg_10_inst : DFFR_X1 port map( D => dp_n685, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_10_port, QN => dp_n552);
   dp_npc_id_i_reg_9_inst : DFFR_X1 port map( D => dp_n684, CK => CLK, RN => 
                           dp_n26, Q => dp_npc_id_o_9_port, QN => dp_n551);
   dp_npc_id_i_reg_8_inst : DFFR_X1 port map( D => dp_n683, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_8_port, QN => dp_n550);
   dp_npc_id_i_reg_7_inst : DFFR_X1 port map( D => dp_n682, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_7_port, QN => dp_n549);
   dp_npc_id_i_reg_6_inst : DFFR_X1 port map( D => dp_n681, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_6_port, QN => dp_n548);
   dp_npc_id_i_reg_5_inst : DFFR_X1 port map( D => dp_n680, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_5_port, QN => dp_n547);
   dp_npc_id_i_reg_4_inst : DFFR_X1 port map( D => dp_n679, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_4_port, QN => dp_n546);
   dp_npc_id_i_reg_3_inst : DFFR_X1 port map( D => dp_n678, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_3_port, QN => dp_n545);
   dp_npc_id_i_reg_2_inst : DFFR_X1 port map( D => dp_n677, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_2_port, QN => dp_n544);
   dp_npc_id_i_reg_1_inst : DFFR_X1 port map( D => dp_n676, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_1_port, QN => dp_n543);
   dp_npc_id_i_reg_0_inst : DFFR_X1 port map( D => dp_n675, CK => CLK, RN => 
                           dp_n27, Q => dp_npc_id_o_0_port, QN => dp_n542);
   dp_ir_reg_25_inst : DFFR_X1 port map( D => dp_n674, CK => CLK, RN => dp_n27,
                           Q => dp_ir_25_port, QN => dp_n541);
   dp_ir_reg_24_inst : DFFR_X1 port map( D => dp_n673, CK => CLK, RN => dp_n27,
                           Q => dp_ir_24_port, QN => dp_n540);
   dp_ir_reg_23_inst : DFFR_X1 port map( D => dp_n672, CK => CLK, RN => dp_n27,
                           Q => dp_ir_23_port, QN => dp_n539);
   dp_ir_reg_22_inst : DFFR_X1 port map( D => dp_n671, CK => CLK, RN => dp_n28,
                           Q => dp_ir_22_port, QN => dp_n538);
   dp_ir_reg_21_inst : DFFR_X1 port map( D => dp_n670, CK => CLK, RN => dp_n28,
                           Q => dp_ir_21_port, QN => dp_n537);
   dp_ir_reg_20_inst : DFFR_X1 port map( D => dp_n669, CK => CLK, RN => dp_n28,
                           Q => dp_ir_20_port, QN => dp_n582);
   dp_ir_reg_19_inst : DFFR_X1 port map( D => dp_n668, CK => CLK, RN => dp_n28,
                           Q => dp_ir_19_port, QN => dp_n580);
   dp_ir_reg_18_inst : DFFR_X1 port map( D => dp_n667, CK => CLK, RN => dp_n28,
                           Q => dp_ir_18_port, QN => dp_n578);
   dp_ir_reg_17_inst : DFFR_X1 port map( D => dp_n666, CK => CLK, RN => dp_n28,
                           Q => dp_ir_17_port, QN => dp_n576);
   dp_ir_reg_16_inst : DFFR_X1 port map( D => dp_n665, CK => CLK, RN => dp_n28,
                           Q => dp_ir_16_port, QN => dp_n574);
   dp_ir_reg_15_inst : DFFR_X1 port map( D => dp_n664, CK => CLK, RN => dp_n28,
                           Q => dp_ir_15_port, QN => dp_n583);
   dp_ir_reg_14_inst : DFFR_X1 port map( D => dp_n663, CK => CLK, RN => dp_n28,
                           Q => dp_ir_14_port, QN => dp_n581);
   dp_ir_reg_13_inst : DFFR_X1 port map( D => dp_n662, CK => CLK, RN => dp_n28,
                           Q => dp_ir_13_port, QN => dp_n579);
   dp_ir_reg_12_inst : DFFR_X1 port map( D => dp_n661, CK => CLK, RN => dp_n28,
                           Q => dp_ir_12_port, QN => dp_n577);
   dp_ir_reg_11_inst : DFFR_X1 port map( D => dp_n660, CK => CLK, RN => dp_n28,
                           Q => dp_ir_11_port, QN => dp_n575);
   dp_ir_reg_10_inst : DFFR_X1 port map( D => dp_n659, CK => CLK, RN => dp_n29,
                           Q => dp_ir_10_port, QN => dp_n536);
   dp_ir_reg_9_inst : DFFR_X1 port map( D => dp_n658, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_9_port, QN => dp_n535);
   dp_ir_reg_8_inst : DFFR_X1 port map( D => dp_n657, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_8_port, QN => dp_n534);
   dp_ir_reg_7_inst : DFFR_X1 port map( D => dp_n656, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_7_port, QN => dp_n533);
   dp_ir_reg_6_inst : DFFR_X1 port map( D => dp_n655, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_6_port, QN => dp_n532);
   dp_ir_reg_5_inst : DFFR_X1 port map( D => dp_n654, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_5_port, QN => dp_n531);
   dp_ir_reg_4_inst : DFFR_X1 port map( D => dp_n653, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_4_port, QN => dp_n530);
   dp_ir_reg_3_inst : DFFR_X1 port map( D => dp_n652, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_3_port, QN => dp_n529);
   dp_ir_reg_2_inst : DFFR_X1 port map( D => dp_n651, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_2_port, QN => dp_n528);
   dp_ir_reg_1_inst : DFFR_X1 port map( D => dp_n650, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_1_port, QN => dp_n527);
   dp_ir_reg_0_inst : DFFR_X1 port map( D => dp_n649, CK => CLK, RN => dp_n29, 
                           Q => dp_ir_0_port, QN => dp_n526);
   dp_alu_out_mem_i_reg_31_inst : DFFR_X1 port map( D => dp_n910, CK => CLK, RN
                           => dp_n29, Q => DRAM_ADDRESS_31_port, QN => dp_n846)
                           ;
   dp_alu_out_mem_i_reg_30_inst : DFFR_X1 port map( D => dp_n911, CK => CLK, RN
                           => dp_n30, Q => DRAM_ADDRESS_30_port, QN => dp_n847)
                           ;
   dp_alu_out_mem_i_reg_29_inst : DFFR_X1 port map( D => dp_n912, CK => CLK, RN
                           => dp_n30, Q => DRAM_ADDRESS_29_port, QN => dp_n848)
                           ;
   dp_alu_out_mem_i_reg_28_inst : DFFR_X1 port map( D => dp_n913, CK => CLK, RN
                           => dp_n30, Q => DRAM_ADDRESS_28_port, QN => dp_n849)
                           ;
   dp_alu_out_mem_i_reg_27_inst : DFFR_X1 port map( D => dp_n914, CK => CLK, RN
                           => dp_n30, Q => DRAM_ADDRESS_27_port, QN => dp_n850)
                           ;
   dp_alu_out_mem_i_reg_26_inst : DFFR_X1 port map( D => dp_n915, CK => CLK, RN
                           => dp_n30, Q => DRAM_ADDRESS_26_port, QN => dp_n851)
                           ;
   dp_alu_out_mem_i_reg_25_inst : DFFR_X1 port map( D => dp_n916, CK => CLK, RN
                           => dp_n30, Q => DRAM_ADDRESS_25_port, QN => dp_n852)
                           ;
   dp_alu_out_mem_i_reg_24_inst : DFFR_X1 port map( D => dp_n917, CK => CLK, RN
                           => dp_n31, Q => DRAM_ADDRESS_24_port, QN => dp_n853)
                           ;
   dp_alu_out_mem_i_reg_23_inst : DFFR_X1 port map( D => dp_n918, CK => CLK, RN
                           => dp_n31, Q => DRAM_ADDRESS_23_port, QN => dp_n854)
                           ;
   dp_alu_out_mem_i_reg_22_inst : DFFR_X1 port map( D => dp_n919, CK => CLK, RN
                           => dp_n31, Q => DRAM_ADDRESS_22_port, QN => dp_n855)
                           ;
   dp_alu_out_mem_i_reg_21_inst : DFFR_X1 port map( D => dp_n920, CK => CLK, RN
                           => dp_n31, Q => DRAM_ADDRESS_21_port, QN => dp_n856)
                           ;
   dp_alu_out_mem_i_reg_20_inst : DFFR_X1 port map( D => dp_n921, CK => CLK, RN
                           => dp_n31, Q => DRAM_ADDRESS_20_port, QN => dp_n857)
                           ;
   dp_alu_out_mem_i_reg_19_inst : DFFR_X1 port map( D => dp_n922, CK => CLK, RN
                           => dp_n31, Q => DRAM_ADDRESS_19_port, QN => dp_n858)
                           ;
   dp_alu_out_mem_i_reg_18_inst : DFFR_X1 port map( D => dp_n923, CK => CLK, RN
                           => dp_n32, Q => DRAM_ADDRESS_18_port, QN => dp_n859)
                           ;
   dp_alu_out_mem_i_reg_17_inst : DFFR_X1 port map( D => dp_n924, CK => CLK, RN
                           => dp_n32, Q => DRAM_ADDRESS_17_port, QN => dp_n860)
                           ;
   dp_alu_out_mem_i_reg_16_inst : DFFR_X1 port map( D => dp_n925, CK => CLK, RN
                           => dp_n32, Q => DRAM_ADDRESS_16_port, QN => dp_n861)
                           ;
   dp_alu_out_mem_i_reg_15_inst : DFFR_X1 port map( D => dp_n926, CK => CLK, RN
                           => dp_n32, Q => DRAM_ADDRESS_15_port, QN => dp_n862)
                           ;
   dp_alu_out_mem_i_reg_14_inst : DFFR_X1 port map( D => dp_n927, CK => CLK, RN
                           => dp_n32, Q => DRAM_ADDRESS_14_port, QN => dp_n863)
                           ;
   dp_alu_out_mem_i_reg_13_inst : DFFR_X1 port map( D => dp_n928, CK => CLK, RN
                           => dp_n32, Q => DRAM_ADDRESS_13_port, QN => dp_n864)
                           ;
   dp_alu_out_mem_i_reg_12_inst : DFFR_X1 port map( D => dp_n929, CK => CLK, RN
                           => dp_n33, Q => DRAM_ADDRESS_12_port, QN => dp_n865)
                           ;
   dp_alu_out_mem_i_reg_11_inst : DFFR_X1 port map( D => dp_n930, CK => CLK, RN
                           => dp_n33, Q => DRAM_ADDRESS_11_port, QN => dp_n866)
                           ;
   dp_alu_out_mem_i_reg_10_inst : DFFR_X1 port map( D => dp_n931, CK => CLK, RN
                           => dp_n33, Q => DRAM_ADDRESS_10_port, QN => dp_n867)
                           ;
   dp_alu_out_mem_i_reg_9_inst : DFFR_X1 port map( D => dp_n932, CK => CLK, RN 
                           => dp_n33, Q => DRAM_ADDRESS_9_port, QN => dp_n868);
   dp_alu_out_mem_i_reg_8_inst : DFFR_X1 port map( D => dp_n933, CK => CLK, RN 
                           => dp_n33, Q => DRAM_ADDRESS_8_port, QN => dp_n869);
   dp_alu_out_mem_i_reg_7_inst : DFFR_X1 port map( D => dp_n934, CK => CLK, RN 
                           => dp_n33, Q => DRAM_ADDRESS_7_port, QN => dp_n870);
   dp_alu_out_mem_i_reg_6_inst : DFFR_X1 port map( D => dp_n935, CK => CLK, RN 
                           => dp_n34, Q => DRAM_ADDRESS_6_port, QN => dp_n871);
   dp_alu_out_mem_i_reg_5_inst : DFFR_X1 port map( D => dp_n936, CK => CLK, RN 
                           => dp_n34, Q => DRAM_ADDRESS_5_port, QN => dp_n872);
   dp_alu_out_mem_i_reg_4_inst : DFFR_X1 port map( D => dp_n937, CK => CLK, RN 
                           => dp_n34, Q => DRAM_ADDRESS_4_port, QN => dp_n873);
   dp_alu_out_mem_i_reg_3_inst : DFFR_X1 port map( D => dp_n938, CK => CLK, RN 
                           => dp_n34, Q => DRAM_ADDRESS_3_port, QN => dp_n874);
   dp_alu_out_mem_i_reg_2_inst : DFFR_X1 port map( D => dp_n939, CK => CLK, RN 
                           => dp_n34, Q => DRAM_ADDRESS_2_port, QN => dp_n875);
   dp_alu_out_mem_i_reg_1_inst : DFFR_X1 port map( D => dp_n940, CK => CLK, RN 
                           => dp_n34, Q => DRAM_ADDRESS_1_port, QN => dp_n876);
   dp_alu_out_mem_i_reg_0_inst : DFFR_X1 port map( D => dp_n941, CK => CLK, RN 
                           => dp_n24, Q => DRAM_ADDRESS_0_port, QN => dp_n877);
   dp_rd_fwd_wb_i_reg_4_inst : DFFR_X1 port map( D => dp_n1005, CK => CLK, RN 
                           => dp_n35, Q => dp_rd_fwd_wb_i_4_port, QN => dp_n524
                           );
   dp_rd_fwd_wb_i_reg_3_inst : DFFR_X1 port map( D => dp_n1006, CK => CLK, RN 
                           => dp_n35, Q => dp_rd_fwd_wb_i_3_port, QN => dp_n522
                           );
   dp_rd_fwd_wb_i_reg_2_inst : DFFR_X1 port map( D => dp_n1007, CK => CLK, RN 
                           => dp_n35, Q => dp_rd_fwd_wb_i_2_port, QN => dp_n520
                           );
   dp_rd_fwd_wb_i_reg_1_inst : DFFR_X1 port map( D => dp_n1008, CK => CLK, RN 
                           => dp_n35, Q => dp_rd_fwd_wb_i_1_port, QN => dp_n518
                           );
   dp_rd_fwd_wb_i_reg_0_inst : DFFR_X1 port map( D => dp_n1009, CK => CLK, RN 
                           => dp_n36, Q => dp_rd_fwd_wb_i_0_port, QN => dp_n516
                           );
   dp_branch_t_mem_i_reg : DFFR_X1 port map( D => dp_n845, CK => CLK, RN => 
                           dp_n36, Q => is_zero_i, QN => dp_n515);
   dp_rf_out1_ex_i_reg_31_inst : DFFR_X1 port map( D => dp_n844, CK => CLK, RN 
                           => dp_n36, Q => dp_rf_out1_ex_i_31_port, QN => 
                           dp_n514);
   dp_rf_out1_ex_i_reg_30_inst : DFFR_X1 port map( D => dp_n843, CK => CLK, RN 
                           => dp_n36, Q => dp_rf_out1_ex_i_30_port, QN => 
                           dp_n513);
   dp_rf_out1_ex_i_reg_29_inst : DFFR_X1 port map( D => dp_n842, CK => CLK, RN 
                           => dp_n36, Q => dp_rf_out1_ex_i_29_port, QN => 
                           dp_n512);
   dp_rf_out1_ex_i_reg_28_inst : DFFR_X1 port map( D => dp_n841, CK => CLK, RN 
                           => dp_n36, Q => dp_rf_out1_ex_i_28_port, QN => 
                           dp_n511);
   dp_rf_out1_ex_i_reg_27_inst : DFFR_X1 port map( D => dp_n840, CK => CLK, RN 
                           => dp_n36, Q => dp_rf_out1_ex_i_27_port, QN => 
                           dp_n510);
   dp_rf_out1_ex_i_reg_26_inst : DFFR_X1 port map( D => dp_n839, CK => CLK, RN 
                           => dp_n36, Q => dp_rf_out1_ex_i_26_port, QN => 
                           dp_n509);
   dp_rf_out1_ex_i_reg_25_inst : DFFR_X1 port map( D => dp_n838, CK => CLK, RN 
                           => dp_n36, Q => dp_rf_out1_ex_i_25_port, QN => 
                           dp_n508);
   dp_rf_out1_ex_i_reg_24_inst : DFFR_X1 port map( D => dp_n837, CK => CLK, RN 
                           => dp_n36, Q => dp_rf_out1_ex_i_24_port, QN => 
                           dp_n507);
   dp_rf_out1_ex_i_reg_23_inst : DFFR_X1 port map( D => dp_n836, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_23_port, QN => 
                           dp_n506);
   dp_rf_out1_ex_i_reg_22_inst : DFFR_X1 port map( D => dp_n835, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_22_port, QN => 
                           dp_n505);
   dp_rf_out1_ex_i_reg_21_inst : DFFR_X1 port map( D => dp_n834, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_21_port, QN => 
                           dp_n504);
   dp_rf_out1_ex_i_reg_20_inst : DFFR_X1 port map( D => dp_n833, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_20_port, QN => 
                           dp_n503);
   dp_rf_out1_ex_i_reg_19_inst : DFFR_X1 port map( D => dp_n832, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_19_port, QN => 
                           dp_n502);
   dp_rf_out1_ex_i_reg_18_inst : DFFR_X1 port map( D => dp_n831, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_18_port, QN => 
                           dp_n501);
   dp_rf_out1_ex_i_reg_17_inst : DFFR_X1 port map( D => dp_n830, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_17_port, QN => 
                           dp_n500);
   dp_rf_out1_ex_i_reg_16_inst : DFFR_X1 port map( D => dp_n829, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_16_port, QN => 
                           dp_n499);
   dp_rf_out1_ex_i_reg_15_inst : DFFR_X1 port map( D => dp_n828, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_15_port, QN => 
                           dp_n498);
   dp_rf_out1_ex_i_reg_14_inst : DFFR_X1 port map( D => dp_n827, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_14_port, QN => 
                           dp_n497);
   dp_rf_out1_ex_i_reg_13_inst : DFFR_X1 port map( D => dp_n826, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_13_port, QN => 
                           dp_n496);
   dp_rf_out1_ex_i_reg_12_inst : DFFR_X1 port map( D => dp_n825, CK => CLK, RN 
                           => dp_n37, Q => dp_rf_out1_ex_i_12_port, QN => 
                           dp_n495);
   dp_rf_out1_ex_i_reg_11_inst : DFFR_X1 port map( D => dp_n824, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_11_port, QN => 
                           dp_n494);
   dp_rf_out1_ex_i_reg_10_inst : DFFR_X1 port map( D => dp_n823, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_10_port, QN => 
                           dp_n493);
   dp_rf_out1_ex_i_reg_9_inst : DFFR_X1 port map( D => dp_n822, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_9_port, QN => 
                           dp_n492);
   dp_rf_out1_ex_i_reg_8_inst : DFFR_X1 port map( D => dp_n821, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_8_port, QN => 
                           dp_n491);
   dp_rf_out1_ex_i_reg_7_inst : DFFR_X1 port map( D => dp_n820, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_7_port, QN => 
                           dp_n490);
   dp_rf_out1_ex_i_reg_6_inst : DFFR_X1 port map( D => dp_n819, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_6_port, QN => 
                           dp_n489);
   dp_rf_out1_ex_i_reg_5_inst : DFFR_X1 port map( D => dp_n818, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_5_port, QN => 
                           dp_n488);
   dp_rf_out1_ex_i_reg_4_inst : DFFR_X1 port map( D => dp_n817, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_4_port, QN => 
                           dp_n487);
   dp_rf_out1_ex_i_reg_3_inst : DFFR_X1 port map( D => dp_n816, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_3_port, QN => 
                           dp_n486);
   dp_rf_out1_ex_i_reg_2_inst : DFFR_X1 port map( D => dp_n815, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_2_port, QN => 
                           dp_n485);
   dp_rf_out1_ex_i_reg_1_inst : DFFR_X1 port map( D => dp_n814, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_1_port, QN => 
                           dp_n484);
   dp_rf_out1_ex_i_reg_0_inst : DFFR_X1 port map( D => dp_n813, CK => CLK, RN 
                           => dp_n38, Q => dp_rf_out1_ex_i_0_port, QN => 
                           dp_n483);
   dp_rf_out2_ex_i_reg_31_inst : DFFR_X1 port map( D => dp_n812, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_31_port, QN => 
                           dp_n482);
   dp_rf_out2_ex_i_reg_30_inst : DFFR_X1 port map( D => dp_n811, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_30_port, QN => 
                           dp_n481);
   dp_rf_out2_ex_i_reg_29_inst : DFFR_X1 port map( D => dp_n810, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_29_port, QN => 
                           dp_n480);
   dp_rf_out2_ex_i_reg_28_inst : DFFR_X1 port map( D => dp_n809, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_28_port, QN => 
                           dp_n479);
   dp_rf_out2_ex_i_reg_27_inst : DFFR_X1 port map( D => dp_n808, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_27_port, QN => 
                           dp_n478);
   dp_rf_out2_ex_i_reg_26_inst : DFFR_X1 port map( D => dp_n807, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_26_port, QN => 
                           dp_n477);
   dp_rf_out2_ex_i_reg_25_inst : DFFR_X1 port map( D => dp_n806, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_25_port, QN => 
                           dp_n476);
   dp_rf_out2_ex_i_reg_24_inst : DFFR_X1 port map( D => dp_n805, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_24_port, QN => 
                           dp_n475);
   dp_rf_out2_ex_i_reg_23_inst : DFFR_X1 port map( D => dp_n804, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_23_port, QN => 
                           dp_n474);
   dp_rf_out2_ex_i_reg_22_inst : DFFR_X1 port map( D => dp_n803, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_22_port, QN => 
                           dp_n473);
   dp_rf_out2_ex_i_reg_21_inst : DFFR_X1 port map( D => dp_n802, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_21_port, QN => 
                           dp_n472);
   dp_rf_out2_ex_i_reg_20_inst : DFFR_X1 port map( D => dp_n801, CK => CLK, RN 
                           => dp_n39, Q => dp_data_mem_ex_o_20_port, QN => 
                           dp_n471);
   dp_rf_out2_ex_i_reg_19_inst : DFFR_X1 port map( D => dp_n800, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_19_port, QN => 
                           dp_n470);
   dp_rf_out2_ex_i_reg_18_inst : DFFR_X1 port map( D => dp_n799, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_18_port, QN => 
                           dp_n469);
   dp_rf_out2_ex_i_reg_17_inst : DFFR_X1 port map( D => dp_n798, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_17_port, QN => 
                           dp_n468);
   dp_rf_out2_ex_i_reg_16_inst : DFFR_X1 port map( D => dp_n797, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_16_port, QN => 
                           dp_n467);
   dp_rf_out2_ex_i_reg_15_inst : DFFR_X1 port map( D => dp_n796, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_15_port, QN => 
                           dp_n466);
   dp_rf_out2_ex_i_reg_14_inst : DFFR_X1 port map( D => dp_n795, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_14_port, QN => 
                           dp_n465);
   dp_rf_out2_ex_i_reg_13_inst : DFFR_X1 port map( D => dp_n794, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_13_port, QN => 
                           dp_n464);
   dp_rf_out2_ex_i_reg_12_inst : DFFR_X1 port map( D => dp_n793, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_12_port, QN => 
                           dp_n463);
   dp_rf_out2_ex_i_reg_11_inst : DFFR_X1 port map( D => dp_n792, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_11_port, QN => 
                           dp_n462);
   dp_rf_out2_ex_i_reg_10_inst : DFFR_X1 port map( D => dp_n791, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_10_port, QN => 
                           dp_n461);
   dp_rf_out2_ex_i_reg_9_inst : DFFR_X1 port map( D => dp_n790, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_9_port, QN => 
                           dp_n460);
   dp_rf_out2_ex_i_reg_8_inst : DFFR_X1 port map( D => dp_n789, CK => CLK, RN 
                           => dp_n40, Q => dp_data_mem_ex_o_8_port, QN => 
                           dp_n459);
   dp_rf_out2_ex_i_reg_7_inst : DFFR_X1 port map( D => dp_n788, CK => CLK, RN 
                           => dp_n41, Q => dp_data_mem_ex_o_7_port, QN => 
                           dp_n458);
   dp_rf_out2_ex_i_reg_6_inst : DFFR_X1 port map( D => dp_n787, CK => CLK, RN 
                           => dp_n41, Q => dp_data_mem_ex_o_6_port, QN => 
                           dp_n457);
   dp_rf_out2_ex_i_reg_5_inst : DFFR_X1 port map( D => dp_n786, CK => CLK, RN 
                           => dp_n41, Q => dp_data_mem_ex_o_5_port, QN => 
                           dp_n456);
   dp_rf_out2_ex_i_reg_4_inst : DFFR_X1 port map( D => dp_n785, CK => CLK, RN 
                           => dp_n41, Q => dp_data_mem_ex_o_4_port, QN => 
                           dp_n455);
   dp_rf_out2_ex_i_reg_3_inst : DFFR_X1 port map( D => dp_n784, CK => CLK, RN 
                           => dp_n41, Q => dp_data_mem_ex_o_3_port, QN => 
                           dp_n454);
   dp_rf_out2_ex_i_reg_2_inst : DFFR_X1 port map( D => dp_n783, CK => CLK, RN 
                           => dp_n41, Q => dp_data_mem_ex_o_2_port, QN => 
                           dp_n453);
   dp_rf_out2_ex_i_reg_1_inst : DFFR_X1 port map( D => dp_n782, CK => CLK, RN 
                           => dp_n41, Q => dp_data_mem_ex_o_1_port, QN => 
                           dp_n452);
   dp_rf_out2_ex_i_reg_0_inst : DFFR_X1 port map( D => dp_n781, CK => CLK, RN 
                           => dp_n41, Q => dp_data_mem_ex_o_0_port, QN => 
                           dp_n451);
   dp_imm_ex_i_reg_31_inst : DFFR_X1 port map( D => dp_n780, CK => CLK, RN => 
                           dp_n41, Q => dp_imm_ex_i_31_port, QN => dp_n450);
   dp_imm_ex_i_reg_30_inst : DFFR_X1 port map( D => dp_n779, CK => CLK, RN => 
                           dp_n41, Q => dp_imm_ex_i_30_port, QN => dp_n449);
   dp_imm_ex_i_reg_29_inst : DFFR_X1 port map( D => dp_n778, CK => CLK, RN => 
                           dp_n41, Q => dp_imm_ex_i_29_port, QN => dp_n448);
   dp_imm_ex_i_reg_28_inst : DFFR_X1 port map( D => dp_n777, CK => CLK, RN => 
                           dp_n41, Q => dp_imm_ex_i_28_port, QN => dp_n447);
   dp_imm_ex_i_reg_27_inst : DFFR_X1 port map( D => dp_n776, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_27_port, QN => dp_n446);
   dp_imm_ex_i_reg_26_inst : DFFR_X1 port map( D => dp_n775, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_26_port, QN => dp_n445);
   dp_imm_ex_i_reg_25_inst : DFFR_X1 port map( D => dp_n774, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_25_port, QN => dp_n444);
   dp_imm_ex_i_reg_24_inst : DFFR_X1 port map( D => dp_n773, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_24_port, QN => dp_n443);
   dp_imm_ex_i_reg_23_inst : DFFR_X1 port map( D => dp_n772, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_23_port, QN => dp_n442);
   dp_imm_ex_i_reg_22_inst : DFFR_X1 port map( D => dp_n771, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_22_port, QN => dp_n441);
   dp_imm_ex_i_reg_21_inst : DFFR_X1 port map( D => dp_n770, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_21_port, QN => dp_n440);
   dp_imm_ex_i_reg_20_inst : DFFR_X1 port map( D => dp_n769, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_20_port, QN => dp_n439);
   dp_imm_ex_i_reg_19_inst : DFFR_X1 port map( D => dp_n768, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_19_port, QN => dp_n438);
   dp_imm_ex_i_reg_18_inst : DFFR_X1 port map( D => dp_n767, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_18_port, QN => dp_n437);
   dp_imm_ex_i_reg_17_inst : DFFR_X1 port map( D => dp_n766, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_17_port, QN => dp_n436);
   dp_imm_ex_i_reg_16_inst : DFFR_X1 port map( D => dp_n765, CK => CLK, RN => 
                           dp_n42, Q => dp_imm_ex_i_16_port, QN => dp_n435);
   dp_imm_ex_i_reg_15_inst : DFFR_X1 port map( D => dp_n764, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_15_port, QN => dp_n434);
   dp_imm_ex_i_reg_14_inst : DFFR_X1 port map( D => dp_n763, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_14_port, QN => dp_n433);
   dp_imm_ex_i_reg_13_inst : DFFR_X1 port map( D => dp_n762, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_13_port, QN => dp_n432);
   dp_imm_ex_i_reg_12_inst : DFFR_X1 port map( D => dp_n761, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_12_port, QN => dp_n431);
   dp_imm_ex_i_reg_11_inst : DFFR_X1 port map( D => dp_n760, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_11_port, QN => dp_n430);
   dp_imm_ex_i_reg_10_inst : DFFR_X1 port map( D => dp_n759, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_10_port, QN => dp_n429);
   dp_imm_ex_i_reg_9_inst : DFFR_X1 port map( D => dp_n758, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_9_port, QN => dp_n428);
   dp_imm_ex_i_reg_8_inst : DFFR_X1 port map( D => dp_n757, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_8_port, QN => dp_n427);
   dp_imm_ex_i_reg_7_inst : DFFR_X1 port map( D => dp_n756, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_7_port, QN => dp_n426);
   dp_imm_ex_i_reg_6_inst : DFFR_X1 port map( D => dp_n755, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_6_port, QN => dp_n425);
   dp_imm_ex_i_reg_5_inst : DFFR_X1 port map( D => dp_n754, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_5_port, QN => dp_n424);
   dp_imm_ex_i_reg_4_inst : DFFR_X1 port map( D => dp_n753, CK => CLK, RN => 
                           dp_n43, Q => dp_imm_ex_i_4_port, QN => dp_n423);
   dp_imm_ex_i_reg_3_inst : DFFR_X1 port map( D => dp_n752, CK => CLK, RN => 
                           dp_n44, Q => dp_imm_ex_i_3_port, QN => dp_n422);
   dp_imm_ex_i_reg_2_inst : DFFR_X1 port map( D => dp_n751, CK => CLK, RN => 
                           dp_n44, Q => dp_imm_ex_i_2_port, QN => dp_n421);
   dp_imm_ex_i_reg_1_inst : DFFR_X1 port map( D => dp_n750, CK => CLK, RN => 
                           dp_n44, Q => dp_imm_ex_i_1_port, QN => dp_n420);
   dp_imm_ex_i_reg_0_inst : DFFR_X1 port map( D => dp_n749, CK => CLK, RN => 
                           dp_n44, Q => dp_imm_ex_i_0_port, QN => dp_n419);
   dp_rd_fwd_ex_i_reg_4_inst : DFFR_X1 port map( D => dp_n716, CK => CLK, RN =>
                           dp_n45, Q => dp_rd_fwd_ex_o_4_port, QN => dp_n418);
   dp_rd_fwd_ex_i_reg_3_inst : DFFR_X1 port map( D => dp_n715, CK => CLK, RN =>
                           dp_n45, Q => dp_rd_fwd_ex_o_3_port, QN => dp_n417);
   dp_rd_fwd_ex_i_reg_2_inst : DFFR_X1 port map( D => dp_n714, CK => CLK, RN =>
                           dp_n45, Q => dp_rd_fwd_ex_o_2_port, QN => dp_n416);
   dp_rd_fwd_ex_i_reg_1_inst : DFFR_X1 port map( D => dp_n713, CK => CLK, RN =>
                           dp_n45, Q => dp_rd_fwd_ex_o_1_port, QN => dp_n415);
   dp_rd_fwd_ex_i_reg_0_inst : DFFR_X1 port map( D => dp_n712, CK => CLK, RN =>
                           dp_n45, Q => dp_rd_fwd_ex_o_0_port, QN => dp_n414);
   dp_if_stage_U59 : INV_X1 port map( A => RST, ZN => dp_if_stage_n41);
   dp_if_stage_U58 : MUX2_X1 port map( A => IRAM_ADDRESS_16_port, B => 
                           dp_npc_if_o_16_port, S => dp_if_stage_n39, Z => 
                           dp_if_stage_n16);
   dp_if_stage_U57 : MUX2_X1 port map( A => IRAM_ADDRESS_17_port, B => 
                           dp_npc_if_o_17_port, S => dp_if_stage_n39, Z => 
                           dp_if_stage_n15);
   dp_if_stage_U56 : MUX2_X1 port map( A => IRAM_ADDRESS_18_port, B => 
                           dp_npc_if_o_18_port, S => dp_if_stage_n39, Z => 
                           dp_if_stage_n14);
   dp_if_stage_U55 : MUX2_X1 port map( A => IRAM_ADDRESS_19_port, B => 
                           dp_npc_if_o_19_port, S => dp_if_stage_n39, Z => 
                           dp_if_stage_n13);
   dp_if_stage_U54 : MUX2_X1 port map( A => IRAM_ADDRESS_20_port, B => 
                           dp_npc_if_o_20_port, S => dp_if_stage_n39, Z => 
                           dp_if_stage_n12);
   dp_if_stage_U53 : MUX2_X1 port map( A => IRAM_ADDRESS_21_port, B => 
                           dp_npc_if_o_21_port, S => dp_if_stage_n39, Z => 
                           dp_if_stage_n11);
   dp_if_stage_U52 : MUX2_X1 port map( A => IRAM_ADDRESS_22_port, B => 
                           dp_npc_if_o_22_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n10);
   dp_if_stage_U51 : MUX2_X1 port map( A => IRAM_ADDRESS_23_port, B => 
                           dp_npc_if_o_23_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n9);
   dp_if_stage_U50 : MUX2_X1 port map( A => IRAM_ADDRESS_24_port, B => 
                           dp_npc_if_o_24_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n8);
   dp_if_stage_U49 : MUX2_X1 port map( A => IRAM_ADDRESS_25_port, B => 
                           dp_npc_if_o_25_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n7);
   dp_if_stage_U48 : MUX2_X1 port map( A => IRAM_ADDRESS_26_port, B => 
                           dp_npc_if_o_26_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n6);
   dp_if_stage_U47 : MUX2_X1 port map( A => IRAM_ADDRESS_27_port, B => 
                           dp_npc_if_o_27_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n5);
   dp_if_stage_U46 : MUX2_X1 port map( A => IRAM_ADDRESS_28_port, B => 
                           dp_npc_if_o_28_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n4);
   dp_if_stage_U45 : MUX2_X1 port map( A => IRAM_ADDRESS_29_port, B => 
                           dp_npc_if_o_29_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n3);
   dp_if_stage_U44 : MUX2_X1 port map( A => IRAM_ADDRESS_30_port, B => 
                           dp_npc_if_o_30_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n2);
   dp_if_stage_U43 : MUX2_X1 port map( A => IRAM_ADDRESS_31_port, B => 
                           dp_npc_if_o_31_port, S => dp_if_stage_n40, Z => 
                           dp_if_stage_n1);
   dp_if_stage_U42 : NAND2_X1 port map( A1 => dp_npc_if_o_0_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n32);
   dp_if_stage_U41 : OAI21_X1 port map( B1 => dp_if_stage_n64, B2 => 
                           dp_if_stage_n39, A => dp_if_stage_n32, ZN => 
                           dp_if_stage_n97);
   dp_if_stage_U40 : NAND2_X1 port map( A1 => dp_npc_if_o_1_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n31);
   dp_if_stage_U39 : OAI21_X1 port map( B1 => dp_if_stage_n63, B2 => 
                           dp_if_stage_n39, A => dp_if_stage_n31, ZN => 
                           dp_if_stage_n95);
   dp_if_stage_U38 : NAND2_X1 port map( A1 => dp_npc_if_o_2_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n30);
   dp_if_stage_U37 : OAI21_X1 port map( B1 => dp_if_stage_n62, B2 => 
                           dp_if_stage_n39, A => dp_if_stage_n30, ZN => 
                           dp_if_stage_n94);
   dp_if_stage_U36 : NAND2_X1 port map( A1 => dp_npc_if_o_3_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n29);
   dp_if_stage_U35 : OAI21_X1 port map( B1 => dp_if_stage_n61, B2 => 
                           dp_if_stage_n39, A => dp_if_stage_n29, ZN => 
                           dp_if_stage_n93);
   dp_if_stage_U34 : NAND2_X1 port map( A1 => dp_npc_if_o_4_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n28);
   dp_if_stage_U33 : OAI21_X1 port map( B1 => dp_if_stage_n60, B2 => 
                           dp_if_stage_n39, A => dp_if_stage_n28, ZN => 
                           dp_if_stage_n92);
   dp_if_stage_U32 : NAND2_X1 port map( A1 => dp_npc_if_o_5_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n27);
   dp_if_stage_U31 : OAI21_X1 port map( B1 => dp_if_stage_n59, B2 => 
                           dp_if_stage_n39, A => dp_if_stage_n27, ZN => 
                           dp_if_stage_n91);
   dp_if_stage_U30 : NAND2_X1 port map( A1 => dp_npc_if_o_6_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n26);
   dp_if_stage_U29 : OAI21_X1 port map( B1 => dp_if_stage_n58, B2 => 
                           dp_if_stage_n39, A => dp_if_stage_n26, ZN => 
                           dp_if_stage_n90);
   dp_if_stage_U28 : NAND2_X1 port map( A1 => dp_npc_if_o_7_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n25);
   dp_if_stage_U27 : OAI21_X1 port map( B1 => dp_if_stage_n57, B2 => 
                           dp_if_stage_n39, A => dp_if_stage_n25, ZN => 
                           dp_if_stage_n89);
   dp_if_stage_U26 : NAND2_X1 port map( A1 => dp_npc_if_o_8_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n24);
   dp_if_stage_U25 : OAI21_X1 port map( B1 => dp_if_stage_n56, B2 => 
                           dp_if_stage_n38, A => dp_if_stage_n24, ZN => 
                           dp_if_stage_n88);
   dp_if_stage_U24 : NAND2_X1 port map( A1 => dp_npc_if_o_9_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n23);
   dp_if_stage_U23 : OAI21_X1 port map( B1 => dp_if_stage_n55, B2 => 
                           dp_if_stage_n38, A => dp_if_stage_n23, ZN => 
                           dp_if_stage_n87);
   dp_if_stage_U22 : NAND2_X1 port map( A1 => dp_npc_if_o_10_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n22);
   dp_if_stage_U21 : OAI21_X1 port map( B1 => dp_if_stage_n54, B2 => 
                           dp_if_stage_n38, A => dp_if_stage_n22, ZN => 
                           dp_if_stage_n86);
   dp_if_stage_U20 : NAND2_X1 port map( A1 => dp_npc_if_o_11_port, A2 => 
                           dp_if_stage_n37, ZN => dp_if_stage_n21);
   dp_if_stage_U19 : OAI21_X1 port map( B1 => dp_if_stage_n53, B2 => 
                           dp_if_stage_n38, A => dp_if_stage_n21, ZN => 
                           dp_if_stage_n85);
   dp_if_stage_U18 : NAND2_X1 port map( A1 => dp_npc_if_o_12_port, A2 => 
                           dp_if_stage_n38, ZN => dp_if_stage_n20);
   dp_if_stage_U17 : OAI21_X1 port map( B1 => dp_if_stage_n52, B2 => 
                           dp_if_stage_n38, A => dp_if_stage_n20, ZN => 
                           dp_if_stage_n84);
   dp_if_stage_U16 : NAND2_X1 port map( A1 => dp_npc_if_o_13_port, A2 => 
                           dp_if_stage_n38, ZN => dp_if_stage_n19);
   dp_if_stage_U15 : OAI21_X1 port map( B1 => dp_if_stage_n51, B2 => 
                           dp_if_stage_n38, A => dp_if_stage_n19, ZN => 
                           dp_if_stage_n83);
   dp_if_stage_U14 : NAND2_X1 port map( A1 => dp_npc_if_o_14_port, A2 => 
                           dp_if_stage_n38, ZN => dp_if_stage_n18);
   dp_if_stage_U13 : OAI21_X1 port map( B1 => dp_if_stage_n50, B2 => 
                           dp_if_stage_n38, A => dp_if_stage_n18, ZN => 
                           dp_if_stage_n82);
   dp_if_stage_U12 : NAND2_X1 port map( A1 => dp_npc_if_o_15_port, A2 => 
                           dp_if_stage_n38, ZN => dp_if_stage_n17);
   dp_if_stage_U11 : OAI21_X1 port map( B1 => dp_if_stage_n49, B2 => 
                           dp_if_stage_n38, A => dp_if_stage_n17, ZN => 
                           dp_if_stage_n81);
   dp_if_stage_U10 : BUF_X1 port map( A => dp_if_stage_n41, Z => 
                           dp_if_stage_n33);
   dp_if_stage_U9 : BUF_X1 port map( A => dp_if_stage_n41, Z => dp_if_stage_n34
                           );
   dp_if_stage_U8 : BUF_X1 port map( A => dp_if_stage_n36, Z => dp_if_stage_n40
                           );
   dp_if_stage_U7 : BUF_X1 port map( A => dp_if_stage_n36, Z => dp_if_stage_n39
                           );
   dp_if_stage_U6 : BUF_X1 port map( A => dp_if_stage_n35, Z => dp_if_stage_n38
                           );
   dp_if_stage_U5 : BUF_X1 port map( A => dp_if_stage_n35, Z => dp_if_stage_n37
                           );
   dp_if_stage_U4 : CLKBUF_X1 port map( A => pipe_ex_mem_en_i, Z => 
                           dp_if_stage_n35);
   dp_if_stage_U3 : CLKBUF_X1 port map( A => pipe_ex_mem_en_i, Z => 
                           dp_if_stage_n36);
   dp_if_stage_PC_i_reg_16_inst : DFFR_X1 port map( D => dp_if_stage_n16, CK =>
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_16_port, QN => n_1140);
   dp_if_stage_PC_i_reg_17_inst : DFFR_X1 port map( D => dp_if_stage_n15, CK =>
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_17_port, QN => n_1141);
   dp_if_stage_PC_i_reg_18_inst : DFFR_X1 port map( D => dp_if_stage_n14, CK =>
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_18_port, QN => n_1142);
   dp_if_stage_PC_i_reg_19_inst : DFFR_X1 port map( D => dp_if_stage_n13, CK =>
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_19_port, QN => n_1143);
   dp_if_stage_PC_i_reg_20_inst : DFFR_X1 port map( D => dp_if_stage_n12, CK =>
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_20_port, QN => n_1144);
   dp_if_stage_PC_i_reg_21_inst : DFFR_X1 port map( D => dp_if_stage_n11, CK =>
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_21_port, QN => n_1145);
   dp_if_stage_PC_i_reg_22_inst : DFFR_X1 port map( D => dp_if_stage_n10, CK =>
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_22_port, QN => n_1146);
   dp_if_stage_PC_i_reg_23_inst : DFFR_X1 port map( D => dp_if_stage_n9, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_23_port, QN => n_1147);
   dp_if_stage_PC_i_reg_24_inst : DFFR_X1 port map( D => dp_if_stage_n8, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_24_port, QN => n_1148);
   dp_if_stage_PC_i_reg_25_inst : DFFR_X1 port map( D => dp_if_stage_n7, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_25_port, QN => n_1149);
   dp_if_stage_PC_i_reg_26_inst : DFFR_X1 port map( D => dp_if_stage_n6, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_26_port, QN => n_1150);
   dp_if_stage_PC_i_reg_27_inst : DFFR_X1 port map( D => dp_if_stage_n5, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_27_port, QN => n_1151);
   dp_if_stage_PC_i_reg_28_inst : DFFR_X1 port map( D => dp_if_stage_n4, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_28_port, QN => n_1152);
   dp_if_stage_PC_i_reg_29_inst : DFFR_X1 port map( D => dp_if_stage_n3, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_29_port, QN => n_1153);
   dp_if_stage_PC_i_reg_30_inst : DFFR_X1 port map( D => dp_if_stage_n2, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_30_port, QN => n_1154);
   dp_if_stage_PC_i_reg_31_inst : DFFR_X1 port map( D => dp_if_stage_n1, CK => 
                           CLK, RN => dp_if_stage_n41, Q => 
                           IRAM_ADDRESS_31_port, QN => n_1155);
   dp_if_stage_n98 <= '0';
   dp_if_stage_PC_i_reg_15_inst : DFFR_X1 port map( D => dp_if_stage_n81, CK =>
                           CLK, RN => dp_if_stage_n34, Q => 
                           IRAM_ADDRESS_15_port, QN => dp_if_stage_n49);
   dp_if_stage_PC_i_reg_14_inst : DFFR_X1 port map( D => dp_if_stage_n82, CK =>
                           CLK, RN => dp_if_stage_n34, Q => 
                           IRAM_ADDRESS_14_port, QN => dp_if_stage_n50);
   dp_if_stage_PC_i_reg_13_inst : DFFR_X1 port map( D => dp_if_stage_n83, CK =>
                           CLK, RN => dp_if_stage_n34, Q => 
                           IRAM_ADDRESS_13_port, QN => dp_if_stage_n51);
   dp_if_stage_PC_i_reg_12_inst : DFFR_X1 port map( D => dp_if_stage_n84, CK =>
                           CLK, RN => dp_if_stage_n34, Q => 
                           IRAM_ADDRESS_12_port, QN => dp_if_stage_n52);
   dp_if_stage_PC_i_reg_11_inst : DFFR_X1 port map( D => dp_if_stage_n85, CK =>
                           CLK, RN => dp_if_stage_n33, Q => 
                           IRAM_ADDRESS_11_port, QN => dp_if_stage_n53);
   dp_if_stage_PC_i_reg_10_inst : DFFR_X1 port map( D => dp_if_stage_n86, CK =>
                           CLK, RN => dp_if_stage_n33, Q => 
                           IRAM_ADDRESS_10_port, QN => dp_if_stage_n54);
   dp_if_stage_PC_i_reg_9_inst : DFFR_X1 port map( D => dp_if_stage_n87, CK => 
                           CLK, RN => dp_if_stage_n33, Q => IRAM_ADDRESS_9_port
                           , QN => dp_if_stage_n55);
   dp_if_stage_PC_i_reg_8_inst : DFFR_X1 port map( D => dp_if_stage_n88, CK => 
                           CLK, RN => dp_if_stage_n33, Q => IRAM_ADDRESS_8_port
                           , QN => dp_if_stage_n56);
   dp_if_stage_PC_i_reg_7_inst : DFFR_X1 port map( D => dp_if_stage_n89, CK => 
                           CLK, RN => dp_if_stage_n33, Q => IRAM_ADDRESS_7_port
                           , QN => dp_if_stage_n57);
   dp_if_stage_PC_i_reg_6_inst : DFFR_X1 port map( D => dp_if_stage_n90, CK => 
                           CLK, RN => dp_if_stage_n33, Q => IRAM_ADDRESS_6_port
                           , QN => dp_if_stage_n58);
   dp_if_stage_PC_i_reg_5_inst : DFFR_X1 port map( D => dp_if_stage_n91, CK => 
                           CLK, RN => dp_if_stage_n33, Q => IRAM_ADDRESS_5_port
                           , QN => dp_if_stage_n59);
   dp_if_stage_PC_i_reg_4_inst : DFFR_X1 port map( D => dp_if_stage_n92, CK => 
                           CLK, RN => dp_if_stage_n33, Q => IRAM_ADDRESS_4_port
                           , QN => dp_if_stage_n60);
   dp_if_stage_PC_i_reg_3_inst : DFFR_X1 port map( D => dp_if_stage_n93, CK => 
                           CLK, RN => dp_if_stage_n33, Q => IRAM_ADDRESS_3_port
                           , QN => dp_if_stage_n61);
   dp_if_stage_PC_i_reg_2_inst : DFFR_X1 port map( D => dp_if_stage_n94, CK => 
                           CLK, RN => dp_if_stage_n33, Q => IRAM_ADDRESS_2_port
                           , QN => dp_if_stage_n62);
   dp_if_stage_PC_i_reg_1_inst : DFFR_X1 port map( D => dp_if_stage_n95, CK => 
                           CLK, RN => dp_if_stage_n33, Q => 
                           dp_if_stage_NPC_4_i_1_port, QN => dp_if_stage_n63);
   dp_if_stage_PC_i_reg_0_inst : DFFR_X1 port map( D => dp_if_stage_n97, CK => 
                           CLK, RN => dp_if_stage_n33, Q => 
                           dp_if_stage_NPC_4_i_0_port, QN => dp_if_stage_n64);
   dp_if_stage_Logic0_port <= '0';
   dp_if_stage_Logic1_port <= '1';
   dp_if_stage_mux_U55 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_31_port, B 
                           => DRAM_ADDRESS_31_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_31_port);
   dp_if_stage_mux_U54 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_30_port, B 
                           => DRAM_ADDRESS_30_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_30_port);
   dp_if_stage_mux_U53 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_29_port, B 
                           => DRAM_ADDRESS_29_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_29_port);
   dp_if_stage_mux_U52 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_28_port, B 
                           => DRAM_ADDRESS_28_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_28_port);
   dp_if_stage_mux_U51 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_27_port, B 
                           => DRAM_ADDRESS_27_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_27_port);
   dp_if_stage_mux_U50 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_26_port, B 
                           => DRAM_ADDRESS_26_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_26_port);
   dp_if_stage_mux_U49 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_25_port, B 
                           => DRAM_ADDRESS_25_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_25_port);
   dp_if_stage_mux_U48 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_24_port, B 
                           => DRAM_ADDRESS_24_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_24_port);
   dp_if_stage_mux_U47 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_23_port, B 
                           => DRAM_ADDRESS_23_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_23_port);
   dp_if_stage_mux_U46 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_22_port, B 
                           => DRAM_ADDRESS_22_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_22_port);
   dp_if_stage_mux_U45 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_21_port, B 
                           => DRAM_ADDRESS_21_port, S => jump_en_i, Z => 
                           dp_npc_if_o_21_port);
   dp_if_stage_mux_U44 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_20_port, B 
                           => DRAM_ADDRESS_20_port, S => jump_en_i, Z => 
                           dp_npc_if_o_20_port);
   dp_if_stage_mux_U43 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_19_port, B 
                           => DRAM_ADDRESS_19_port, S => jump_en_i, Z => 
                           dp_npc_if_o_19_port);
   dp_if_stage_mux_U42 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_18_port, B 
                           => DRAM_ADDRESS_18_port, S => jump_en_i, Z => 
                           dp_npc_if_o_18_port);
   dp_if_stage_mux_U41 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_17_port, B 
                           => DRAM_ADDRESS_17_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_17_port);
   dp_if_stage_mux_U40 : MUX2_X1 port map( A => dp_if_stage_NPC_4_i_16_port, B 
                           => DRAM_ADDRESS_16_port, S => dp_if_stage_mux_n1, Z 
                           => dp_npc_if_o_16_port);
   dp_if_stage_mux_U39 : INV_X1 port map( A => jump_en_i, ZN => 
                           dp_if_stage_mux_n7);
   dp_if_stage_mux_U38 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_1_port, 
                           A2 => dp_if_stage_mux_n3, B1 => DRAM_ADDRESS_1_port,
                           B2 => jump_en_i, ZN => dp_if_stage_mux_n54);
   dp_if_stage_mux_U37 : INV_X1 port map( A => dp_if_stage_mux_n54, ZN => 
                           dp_npc_if_o_1_port);
   dp_if_stage_mux_U36 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_2_port, 
                           A2 => dp_if_stage_mux_n4, B1 => DRAM_ADDRESS_2_port,
                           B2 => jump_en_i, ZN => dp_if_stage_mux_n43);
   dp_if_stage_mux_U35 : INV_X1 port map( A => dp_if_stage_mux_n43, ZN => 
                           dp_npc_if_o_2_port);
   dp_if_stage_mux_U34 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_3_port, 
                           A2 => dp_if_stage_mux_n4, B1 => DRAM_ADDRESS_3_port,
                           B2 => dp_if_stage_mux_n1, ZN => dp_if_stage_mux_n40)
                           ;
   dp_if_stage_mux_U33 : INV_X1 port map( A => dp_if_stage_mux_n40, ZN => 
                           dp_npc_if_o_3_port);
   dp_if_stage_mux_U32 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_4_port, 
                           A2 => dp_if_stage_mux_n4, B1 => DRAM_ADDRESS_4_port,
                           B2 => dp_if_stage_mux_n1, ZN => dp_if_stage_mux_n39)
                           ;
   dp_if_stage_mux_U31 : INV_X1 port map( A => dp_if_stage_mux_n39, ZN => 
                           dp_npc_if_o_4_port);
   dp_if_stage_mux_U30 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_5_port, 
                           A2 => dp_if_stage_mux_n4, B1 => DRAM_ADDRESS_5_port,
                           B2 => dp_if_stage_mux_n1, ZN => dp_if_stage_mux_n38)
                           ;
   dp_if_stage_mux_U29 : INV_X1 port map( A => dp_if_stage_mux_n38, ZN => 
                           dp_npc_if_o_5_port);
   dp_if_stage_mux_U28 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_6_port, 
                           A2 => dp_if_stage_mux_n5, B1 => DRAM_ADDRESS_6_port,
                           B2 => dp_if_stage_mux_n1, ZN => dp_if_stage_mux_n37)
                           ;
   dp_if_stage_mux_U27 : INV_X1 port map( A => dp_if_stage_mux_n37, ZN => 
                           dp_npc_if_o_6_port);
   dp_if_stage_mux_U26 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_8_port, 
                           A2 => dp_if_stage_mux_n5, B1 => DRAM_ADDRESS_8_port,
                           B2 => jump_en_i, ZN => dp_if_stage_mux_n35);
   dp_if_stage_mux_U25 : INV_X1 port map( A => dp_if_stage_mux_n35, ZN => 
                           dp_npc_if_o_8_port);
   dp_if_stage_mux_U24 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_12_port, 
                           A2 => dp_if_stage_mux_n2, B1 => DRAM_ADDRESS_12_port
                           , B2 => jump_en_i, ZN => dp_if_stage_mux_n62);
   dp_if_stage_mux_U23 : INV_X1 port map( A => dp_if_stage_mux_n62, ZN => 
                           dp_npc_if_o_12_port);
   dp_if_stage_mux_U22 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_13_port, 
                           A2 => dp_if_stage_mux_n3, B1 => DRAM_ADDRESS_13_port
                           , B2 => jump_en_i, ZN => dp_if_stage_mux_n61);
   dp_if_stage_mux_U21 : INV_X1 port map( A => dp_if_stage_mux_n61, ZN => 
                           dp_npc_if_o_13_port);
   dp_if_stage_mux_U20 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_14_port, 
                           A2 => dp_if_stage_mux_n3, B1 => DRAM_ADDRESS_14_port
                           , B2 => jump_en_i, ZN => dp_if_stage_mux_n60);
   dp_if_stage_mux_U19 : INV_X1 port map( A => dp_if_stage_mux_n60, ZN => 
                           dp_npc_if_o_14_port);
   dp_if_stage_mux_U18 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_15_port, 
                           A2 => dp_if_stage_mux_n3, B1 => DRAM_ADDRESS_15_port
                           , B2 => jump_en_i, ZN => dp_if_stage_mux_n59);
   dp_if_stage_mux_U17 : INV_X1 port map( A => dp_if_stage_mux_n59, ZN => 
                           dp_npc_if_o_15_port);
   dp_if_stage_mux_U16 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_0_port, 
                           A2 => dp_if_stage_mux_n2, B1 => DRAM_ADDRESS_0_port,
                           B2 => dp_if_stage_mux_n1, ZN => dp_if_stage_mux_n65)
                           ;
   dp_if_stage_mux_U15 : INV_X1 port map( A => dp_if_stage_mux_n65, ZN => 
                           dp_npc_if_o_0_port);
   dp_if_stage_mux_U14 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_10_port, 
                           A2 => dp_if_stage_mux_n2, B1 => DRAM_ADDRESS_10_port
                           , B2 => dp_if_stage_mux_n1, ZN => 
                           dp_if_stage_mux_n64);
   dp_if_stage_mux_U13 : INV_X1 port map( A => dp_if_stage_mux_n64, ZN => 
                           dp_npc_if_o_10_port);
   dp_if_stage_mux_U12 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_11_port, 
                           A2 => dp_if_stage_mux_n2, B1 => DRAM_ADDRESS_11_port
                           , B2 => dp_if_stage_mux_n1, ZN => 
                           dp_if_stage_mux_n63);
   dp_if_stage_mux_U11 : INV_X1 port map( A => dp_if_stage_mux_n63, ZN => 
                           dp_npc_if_o_11_port);
   dp_if_stage_mux_U10 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_9_port, 
                           A2 => dp_if_stage_mux_n5, B1 => dp_if_stage_mux_n1, 
                           B2 => DRAM_ADDRESS_9_port, ZN => dp_if_stage_mux_n34
                           );
   dp_if_stage_mux_U9 : INV_X1 port map( A => dp_if_stage_mux_n34, ZN => 
                           dp_npc_if_o_9_port);
   dp_if_stage_mux_U8 : AOI22_X1 port map( A1 => dp_if_stage_NPC_4_i_7_port, A2
                           => dp_if_stage_mux_n5, B1 => DRAM_ADDRESS_7_port, B2
                           => dp_if_stage_mux_n1, ZN => dp_if_stage_mux_n36);
   dp_if_stage_mux_U7 : INV_X1 port map( A => dp_if_stage_mux_n36, ZN => 
                           dp_npc_if_o_7_port);
   dp_if_stage_mux_U6 : BUF_X1 port map( A => dp_if_stage_mux_n7, Z => 
                           dp_if_stage_mux_n6);
   dp_if_stage_mux_U5 : BUF_X1 port map( A => dp_if_stage_mux_n7, Z => 
                           dp_if_stage_mux_n2);
   dp_if_stage_mux_U4 : BUF_X1 port map( A => dp_if_stage_mux_n7, Z => 
                           dp_if_stage_mux_n3);
   dp_if_stage_mux_U3 : BUF_X1 port map( A => dp_if_stage_mux_n7, Z => 
                           dp_if_stage_mux_n4);
   dp_if_stage_mux_U2 : BUF_X1 port map( A => dp_if_stage_mux_n7, Z => 
                           dp_if_stage_mux_n5);
   dp_if_stage_mux_U1 : INV_X1 port map( A => dp_if_stage_mux_n6, ZN => 
                           dp_if_stage_mux_n1);
   dp_if_stage_add_77_U91 : XNOR2_X1 port map( A => dp_if_stage_add_77_n58, B 
                           => dp_if_stage_add_77_n56, ZN => 
                           dp_if_stage_NPC_4_i_10_port);
   dp_if_stage_add_77_U90 : XNOR2_X1 port map( A => dp_if_stage_add_77_n57, B 
                           => dp_if_stage_add_77_n55, ZN => 
                           dp_if_stage_NPC_4_i_11_port);
   dp_if_stage_add_77_U89 : INV_X1 port map( A => dp_if_stage_add_77_n11, ZN =>
                           dp_if_stage_add_77_n54);
   dp_if_stage_add_77_U88 : XNOR2_X1 port map( A => dp_if_stage_add_77_n52, B 
                           => dp_if_stage_add_77_n51, ZN => 
                           dp_if_stage_NPC_4_i_13_port);
   dp_if_stage_add_77_U87 : XNOR2_X1 port map( A => dp_if_stage_add_77_n50, B 
                           => dp_if_stage_add_77_n48, ZN => 
                           dp_if_stage_NPC_4_i_15_port);
   dp_if_stage_add_77_U86 : INV_X1 port map( A => dp_if_stage_add_77_n47, ZN =>
                           dp_if_stage_add_77_n44);
   dp_if_stage_add_77_U85 : NAND3_X1 port map( A1 => IRAM_ADDRESS_18_port, A2 
                           => IRAM_ADDRESS_19_port, A3 => IRAM_ADDRESS_17_port,
                           ZN => dp_if_stage_add_77_n38);
   dp_if_stage_add_77_U84 : NAND3_X1 port map( A1 => IRAM_ADDRESS_22_port, A2 
                           => IRAM_ADDRESS_23_port, A3 => IRAM_ADDRESS_21_port,
                           ZN => dp_if_stage_add_77_n32);
   dp_if_stage_add_77_U83 : NAND3_X1 port map( A1 => IRAM_ADDRESS_26_port, A2 
                           => IRAM_ADDRESS_27_port, A3 => IRAM_ADDRESS_25_port,
                           ZN => dp_if_stage_add_77_n26);
   dp_if_stage_add_77_U82 : XNOR2_X1 port map( A => dp_if_stage_add_77_n14, B 
                           => dp_if_stage_add_77_n13, ZN => 
                           dp_if_stage_NPC_4_i_5_port);
   dp_if_stage_add_77_U81 : XNOR2_X1 port map( A => dp_if_stage_add_77_n59, B 
                           => dp_if_stage_add_77_n11, ZN => 
                           dp_if_stage_NPC_4_i_8_port);
   dp_if_stage_add_77_U80 : XNOR2_X1 port map( A => dp_if_stage_add_77_n10, B 
                           => IRAM_ADDRESS_9_port, ZN => 
                           dp_if_stage_NPC_4_i_9_port);
   dp_if_stage_add_77_U79 : INV_X1 port map( A => IRAM_ADDRESS_31_port, ZN => 
                           dp_if_stage_add_77_n18);
   dp_if_stage_add_77_U78 : INV_X1 port map( A => IRAM_ADDRESS_9_port, ZN => 
                           dp_if_stage_add_77_n61);
   dp_if_stage_add_77_U77 : INV_X1 port map( A => IRAM_ADDRESS_19_port, ZN => 
                           dp_if_stage_add_77_n39);
   dp_if_stage_add_77_U76 : INV_X1 port map( A => IRAM_ADDRESS_23_port, ZN => 
                           dp_if_stage_add_77_n33);
   dp_if_stage_add_77_U75 : INV_X1 port map( A => IRAM_ADDRESS_27_port, ZN => 
                           dp_if_stage_add_77_n27);
   dp_if_stage_add_77_U74 : INV_X1 port map( A => IRAM_ADDRESS_29_port, ZN => 
                           dp_if_stage_add_77_n23);
   dp_if_stage_add_77_U73 : INV_X1 port map( A => IRAM_ADDRESS_11_port, ZN => 
                           dp_if_stage_add_77_n57);
   dp_if_stage_add_77_U72 : INV_X1 port map( A => IRAM_ADDRESS_30_port, ZN => 
                           dp_if_stage_add_77_n20);
   dp_if_stage_add_77_U71 : INV_X1 port map( A => IRAM_ADDRESS_28_port, ZN => 
                           dp_if_stage_add_77_n24);
   dp_if_stage_add_77_U70 : INV_X1 port map( A => IRAM_ADDRESS_20_port, ZN => 
                           dp_if_stage_add_77_n36);
   dp_if_stage_add_77_U69 : INV_X1 port map( A => IRAM_ADDRESS_24_port, ZN => 
                           dp_if_stage_add_77_n30);
   dp_if_stage_add_77_U68 : INV_X1 port map( A => IRAM_ADDRESS_5_port, ZN => 
                           dp_if_stage_add_77_n14);
   dp_if_stage_add_77_U67 : INV_X1 port map( A => IRAM_ADDRESS_13_port, ZN => 
                           dp_if_stage_add_77_n52);
   dp_if_stage_add_77_U66 : INV_X1 port map( A => IRAM_ADDRESS_15_port, ZN => 
                           dp_if_stage_add_77_n50);
   dp_if_stage_add_77_U65 : INV_X1 port map( A => IRAM_ADDRESS_10_port, ZN => 
                           dp_if_stage_add_77_n58);
   dp_if_stage_add_77_U64 : INV_X1 port map( A => IRAM_ADDRESS_4_port, ZN => 
                           dp_if_stage_add_77_n60);
   dp_if_stage_add_77_U63 : XNOR2_X1 port map( A => dp_if_stage_add_77_n35, B 
                           => dp_if_stage_add_77_n36, ZN => 
                           dp_if_stage_NPC_4_i_20_port);
   dp_if_stage_add_77_U62 : XNOR2_X1 port map( A => dp_if_stage_add_77_n29, B 
                           => dp_if_stage_add_77_n30, ZN => 
                           dp_if_stage_NPC_4_i_24_port);
   dp_if_stage_add_77_U61 : XNOR2_X1 port map( A => dp_if_stage_add_77_n22, B 
                           => dp_if_stage_add_77_n24, ZN => 
                           dp_if_stage_NPC_4_i_28_port);
   dp_if_stage_add_77_U60 : XNOR2_X1 port map( A => dp_if_stage_add_77_n19, B 
                           => dp_if_stage_add_77_n20, ZN => 
                           dp_if_stage_NPC_4_i_30_port);
   dp_if_stage_add_77_U59 : XOR2_X1 port map( A => dp_if_stage_add_77_n7, B => 
                           IRAM_ADDRESS_18_port, Z => 
                           dp_if_stage_NPC_4_i_18_port);
   dp_if_stage_add_77_U58 : AND2_X1 port map( A1 => IRAM_ADDRESS_18_port, A2 =>
                           dp_if_stage_add_77_n7, ZN => dp_if_stage_add_77_n9);
   dp_if_stage_add_77_U57 : XNOR2_X1 port map( A => dp_if_stage_add_77_n9, B =>
                           dp_if_stage_add_77_n39, ZN => 
                           dp_if_stage_NPC_4_i_19_port);
   dp_if_stage_add_77_U56 : XOR2_X1 port map( A => IRAM_ADDRESS_21_port, B => 
                           dp_if_stage_add_77_n34, Z => 
                           dp_if_stage_NPC_4_i_21_port);
   dp_if_stage_add_77_U55 : XOR2_X1 port map( A => IRAM_ADDRESS_16_port, B => 
                           dp_if_stage_add_77_n41, Z => 
                           dp_if_stage_NPC_4_i_16_port);
   dp_if_stage_add_77_U54 : XOR2_X1 port map( A => IRAM_ADDRESS_17_port, B => 
                           dp_if_stage_add_77_n40, Z => 
                           dp_if_stage_NPC_4_i_17_port);
   dp_if_stage_add_77_U53 : XOR2_X1 port map( A => dp_if_stage_add_77_n6, B => 
                           IRAM_ADDRESS_22_port, Z => 
                           dp_if_stage_NPC_4_i_22_port);
   dp_if_stage_add_77_U52 : XOR2_X1 port map( A => IRAM_ADDRESS_25_port, B => 
                           dp_if_stage_add_77_n28, Z => 
                           dp_if_stage_NPC_4_i_25_port);
   dp_if_stage_add_77_U51 : XOR2_X1 port map( A => dp_if_stage_add_77_n5, B => 
                           IRAM_ADDRESS_26_port, Z => 
                           dp_if_stage_NPC_4_i_26_port);
   dp_if_stage_add_77_U50 : XNOR2_X1 port map( A => IRAM_ADDRESS_29_port, B => 
                           dp_if_stage_add_77_n21, ZN => 
                           dp_if_stage_NPC_4_i_29_port);
   dp_if_stage_add_77_U49 : INV_X1 port map( A => IRAM_ADDRESS_2_port, ZN => 
                           dp_if_stage_NPC_4_i_2_port);
   dp_if_stage_add_77_U48 : INV_X1 port map( A => IRAM_ADDRESS_8_port, ZN => 
                           dp_if_stage_add_77_n59);
   dp_if_stage_add_77_U47 : INV_X1 port map( A => IRAM_ADDRESS_3_port, ZN => 
                           dp_if_stage_add_77_n16);
   dp_if_stage_add_77_U46 : AND2_X1 port map( A1 => IRAM_ADDRESS_6_port, A2 => 
                           dp_if_stage_add_77_n12, ZN => dp_if_stage_add_77_n8)
                           ;
   dp_if_stage_add_77_U45 : AND2_X1 port map( A1 => IRAM_ADDRESS_17_port, A2 =>
                           dp_if_stage_add_77_n40, ZN => dp_if_stage_add_77_n7)
                           ;
   dp_if_stage_add_77_U44 : AND2_X1 port map( A1 => IRAM_ADDRESS_21_port, A2 =>
                           dp_if_stage_add_77_n34, ZN => dp_if_stage_add_77_n6)
                           ;
   dp_if_stage_add_77_U43 : AND2_X1 port map( A1 => IRAM_ADDRESS_25_port, A2 =>
                           dp_if_stage_add_77_n28, ZN => dp_if_stage_add_77_n5)
                           ;
   dp_if_stage_add_77_U42 : NAND2_X1 port map( A1 => dp_if_stage_add_77_n11, A2
                           => IRAM_ADDRESS_8_port, ZN => dp_if_stage_add_77_n10
                           );
   dp_if_stage_add_77_U41 : NAND2_X1 port map( A1 => dp_if_stage_add_77_n29, A2
                           => IRAM_ADDRESS_24_port, ZN => 
                           dp_if_stage_add_77_n25);
   dp_if_stage_add_77_U40 : NAND2_X1 port map( A1 => dp_if_stage_add_77_n35, A2
                           => IRAM_ADDRESS_20_port, ZN => 
                           dp_if_stage_add_77_n31);
   dp_if_stage_add_77_U39 : NAND2_X1 port map( A1 => dp_if_stage_add_77_n41, A2
                           => IRAM_ADDRESS_16_port, ZN => 
                           dp_if_stage_add_77_n37);
   dp_if_stage_add_77_U38 : NAND2_X1 port map( A1 => dp_if_stage_add_77_n22, A2
                           => IRAM_ADDRESS_28_port, ZN => 
                           dp_if_stage_add_77_n21);
   dp_if_stage_add_77_U37 : AND2_X1 port map( A1 => dp_if_stage_add_77_n56, A2 
                           => IRAM_ADDRESS_10_port, ZN => 
                           dp_if_stage_add_77_n55);
   dp_if_stage_add_77_U36 : AND2_X1 port map( A1 => dp_if_stage_add_77_n49, A2 
                           => IRAM_ADDRESS_14_port, ZN => 
                           dp_if_stage_add_77_n48);
   dp_if_stage_add_77_U35 : OR2_X1 port map( A1 => dp_if_stage_NPC_4_i_2_port, 
                           A2 => dp_if_stage_add_77_n16, ZN => 
                           dp_if_stage_add_77_n4);
   dp_if_stage_add_77_U34 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n60, A2 
                           => dp_if_stage_add_77_n4, ZN => 
                           dp_if_stage_add_77_n13);
   dp_if_stage_add_77_U33 : AND2_X1 port map( A1 => IRAM_ADDRESS_12_port, A2 =>
                           dp_if_stage_add_77_n53, ZN => dp_if_stage_add_77_n51
                           );
   dp_if_stage_add_77_U32 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n23, A2 
                           => dp_if_stage_add_77_n21, ZN => 
                           dp_if_stage_add_77_n19);
   dp_if_stage_add_77_U31 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n25, A2 
                           => dp_if_stage_add_77_n26, ZN => 
                           dp_if_stage_add_77_n22);
   dp_if_stage_add_77_U30 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n31, A2 
                           => dp_if_stage_add_77_n32, ZN => 
                           dp_if_stage_add_77_n29);
   dp_if_stage_add_77_U29 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n37, A2 
                           => dp_if_stage_add_77_n38, ZN => 
                           dp_if_stage_add_77_n35);
   dp_if_stage_add_77_U28 : NAND4_X1 port map( A1 => IRAM_ADDRESS_11_port, A2 
                           => IRAM_ADDRESS_10_port, A3 => IRAM_ADDRESS_9_port, 
                           A4 => IRAM_ADDRESS_8_port, ZN => 
                           dp_if_stage_add_77_n47);
   dp_if_stage_add_77_U27 : NAND2_X1 port map( A1 => dp_if_stage_add_77_n44, A2
                           => dp_if_stage_add_77_n45, ZN => 
                           dp_if_stage_add_77_n42);
   dp_if_stage_add_77_U26 : NAND4_X1 port map( A1 => IRAM_ADDRESS_12_port, A2 
                           => IRAM_ADDRESS_13_port, A3 => IRAM_ADDRESS_14_port,
                           A4 => IRAM_ADDRESS_15_port, ZN => 
                           dp_if_stage_add_77_n43);
   dp_if_stage_add_77_U25 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n42, A2 
                           => dp_if_stage_add_77_n43, ZN => 
                           dp_if_stage_add_77_n41);
   dp_if_stage_add_77_U24 : NAND4_X1 port map( A1 => IRAM_ADDRESS_4_port, A2 =>
                           IRAM_ADDRESS_5_port, A3 => IRAM_ADDRESS_6_port, A4 
                           => IRAM_ADDRESS_7_port, ZN => dp_if_stage_add_77_n46
                           );
   dp_if_stage_add_77_U23 : AND2_X1 port map( A1 => dp_if_stage_add_77_n51, A2 
                           => IRAM_ADDRESS_13_port, ZN => 
                           dp_if_stage_add_77_n49);
   dp_if_stage_add_77_U22 : AND2_X1 port map( A1 => dp_if_stage_add_77_n13, A2 
                           => IRAM_ADDRESS_5_port, ZN => dp_if_stage_add_77_n12
                           );
   dp_if_stage_add_77_U21 : INV_X1 port map( A => dp_if_stage_add_77_n4, ZN => 
                           dp_if_stage_add_77_n15);
   dp_if_stage_add_77_U20 : INV_X1 port map( A => dp_if_stage_add_77_n31, ZN =>
                           dp_if_stage_add_77_n34);
   dp_if_stage_add_77_U19 : INV_X1 port map( A => dp_if_stage_add_77_n25, ZN =>
                           dp_if_stage_add_77_n28);
   dp_if_stage_add_77_U18 : INV_X1 port map( A => dp_if_stage_add_77_n37, ZN =>
                           dp_if_stage_add_77_n40);
   dp_if_stage_add_77_U17 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n4, A2 
                           => dp_if_stage_add_77_n46, ZN => 
                           dp_if_stage_add_77_n45);
   dp_if_stage_add_77_U16 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n61, A2 
                           => dp_if_stage_add_77_n10, ZN => 
                           dp_if_stage_add_77_n56);
   dp_if_stage_add_77_U15 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n54, A2 
                           => dp_if_stage_add_77_n47, ZN => 
                           dp_if_stage_add_77_n53);
   dp_if_stage_add_77_U14 : NOR2_X1 port map( A1 => dp_if_stage_add_77_n4, A2 
                           => dp_if_stage_add_77_n46, ZN => 
                           dp_if_stage_add_77_n11);
   dp_if_stage_add_77_U13 : XOR2_X1 port map( A => dp_if_stage_add_77_n16, B =>
                           dp_if_stage_NPC_4_i_2_port, Z => 
                           dp_if_stage_NPC_4_i_3_port);
   dp_if_stage_add_77_U12 : XOR2_X1 port map( A => IRAM_ADDRESS_4_port, B => 
                           dp_if_stage_add_77_n15, Z => 
                           dp_if_stage_NPC_4_i_4_port);
   dp_if_stage_add_77_U11 : XOR2_X1 port map( A => IRAM_ADDRESS_6_port, B => 
                           dp_if_stage_add_77_n12, Z => 
                           dp_if_stage_NPC_4_i_6_port);
   dp_if_stage_add_77_U10 : XOR2_X1 port map( A => IRAM_ADDRESS_7_port, B => 
                           dp_if_stage_add_77_n8, Z => 
                           dp_if_stage_NPC_4_i_7_port);
   dp_if_stage_add_77_U9 : XOR2_X1 port map( A => IRAM_ADDRESS_12_port, B => 
                           dp_if_stage_add_77_n53, Z => 
                           dp_if_stage_NPC_4_i_12_port);
   dp_if_stage_add_77_U8 : XOR2_X1 port map( A => IRAM_ADDRESS_14_port, B => 
                           dp_if_stage_add_77_n49, Z => 
                           dp_if_stage_NPC_4_i_14_port);
   dp_if_stage_add_77_U7 : NAND2_X1 port map( A1 => IRAM_ADDRESS_22_port, A2 =>
                           dp_if_stage_add_77_n6, ZN => dp_if_stage_add_77_n3);
   dp_if_stage_add_77_U6 : XOR2_X1 port map( A => dp_if_stage_add_77_n3, B => 
                           dp_if_stage_add_77_n33, Z => 
                           dp_if_stage_NPC_4_i_23_port);
   dp_if_stage_add_77_U5 : NAND2_X1 port map( A1 => IRAM_ADDRESS_26_port, A2 =>
                           dp_if_stage_add_77_n5, ZN => dp_if_stage_add_77_n2);
   dp_if_stage_add_77_U4 : XOR2_X1 port map( A => dp_if_stage_add_77_n2, B => 
                           dp_if_stage_add_77_n27, Z => 
                           dp_if_stage_NPC_4_i_27_port);
   dp_if_stage_add_77_U3 : NAND2_X1 port map( A1 => dp_if_stage_add_77_n19, A2 
                           => IRAM_ADDRESS_30_port, ZN => dp_if_stage_add_77_n1
                           );
   dp_if_stage_add_77_U2 : XOR2_X1 port map( A => dp_if_stage_add_77_n1, B => 
                           dp_if_stage_add_77_n18, Z => 
                           dp_if_stage_NPC_4_i_31_port);
   dp_id_stage_U147 : XOR2_X1 port map( A => dp_rd_fwd_wb_i_4_port, B => 
                           dp_id_stage_n27, Z => dp_id_stage_p_addr_wRD_4_port)
                           ;
   dp_id_stage_U146 : NOR2_X1 port map( A1 => dp_rd_fwd_wb_i_3_port, A2 => 
                           dp_id_stage_n26, ZN => dp_id_stage_n27);
   dp_id_stage_U145 : XNOR2_X1 port map( A => dp_rd_fwd_wb_i_3_port, B => 
                           dp_id_stage_n26, ZN => dp_id_stage_p_addr_wRD_3_port
                           );
   dp_id_stage_U144 : OAI21_X1 port map( B1 => dp_id_stage_n25, B2 => 
                           dp_id_stage_n28, A => dp_id_stage_n26, ZN => 
                           dp_id_stage_p_addr_wRD_2_port);
   dp_id_stage_U143 : NAND2_X1 port map( A1 => dp_id_stage_n25, A2 => 
                           dp_id_stage_n28, ZN => dp_id_stage_n26);
   dp_id_stage_U142 : AOI21_X1 port map( B1 => dp_rd_fwd_wb_i_0_port, B2 => 
                           dp_rd_fwd_wb_i_1_port, A => dp_id_stage_n25, ZN => 
                           dp_id_stage_n24);
   dp_id_stage_U141 : NOR2_X1 port map( A1 => dp_rd_fwd_wb_i_1_port, A2 => 
                           dp_rd_fwd_wb_i_0_port, ZN => dp_id_stage_n25);
   dp_id_stage_U140 : XOR2_X1 port map( A => dp_ir_20_port, B => 
                           dp_id_stage_n15, Z => dp_id_stage_p_addr_wRS2_4_port
                           );
   dp_id_stage_U139 : NOR2_X1 port map( A1 => dp_ir_19_port, A2 => 
                           dp_id_stage_n14, ZN => dp_id_stage_n15);
   dp_id_stage_U138 : XNOR2_X1 port map( A => dp_ir_19_port, B => 
                           dp_id_stage_n14, ZN => 
                           dp_id_stage_p_addr_wRS2_3_port);
   dp_id_stage_U137 : OAI21_X1 port map( B1 => dp_id_stage_n13, B2 => 
                           dp_id_stage_n16, A => dp_id_stage_n14, ZN => 
                           dp_id_stage_p_addr_wRS2_2_port);
   dp_id_stage_U136 : NAND2_X1 port map( A1 => dp_id_stage_n13, A2 => 
                           dp_id_stage_n16, ZN => dp_id_stage_n14);
   dp_id_stage_U135 : AOI21_X1 port map( B1 => dp_ir_16_port, B2 => 
                           dp_ir_17_port, A => dp_id_stage_n13, ZN => 
                           dp_id_stage_n12);
   dp_id_stage_U134 : NOR2_X1 port map( A1 => dp_ir_17_port, A2 => 
                           dp_ir_16_port, ZN => dp_id_stage_n13);
   dp_id_stage_U133 : XOR2_X1 port map( A => dp_ir_25_port, B => 
                           dp_id_stage_n10, Z => dp_id_stage_p_addr_wRS1_4_port
                           );
   dp_id_stage_U132 : NOR2_X1 port map( A1 => dp_ir_24_port, A2 => 
                           dp_id_stage_n9, ZN => dp_id_stage_n10);
   dp_id_stage_U131 : XNOR2_X1 port map( A => dp_ir_24_port, B => 
                           dp_id_stage_n9, ZN => dp_id_stage_p_addr_wRS1_3_port
                           );
   dp_id_stage_U130 : OAI21_X1 port map( B1 => dp_id_stage_n8, B2 => 
                           dp_id_stage_n11, A => dp_id_stage_n9, ZN => 
                           dp_id_stage_p_addr_wRS1_2_port);
   dp_id_stage_U129 : NAND2_X1 port map( A1 => dp_id_stage_n8, A2 => 
                           dp_id_stage_n11, ZN => dp_id_stage_n9);
   dp_id_stage_U128 : AOI21_X1 port map( B1 => dp_ir_21_port, B2 => 
                           dp_ir_22_port, A => dp_id_stage_n8, ZN => 
                           dp_id_stage_n7);
   dp_id_stage_U127 : NOR2_X1 port map( A1 => dp_ir_22_port, A2 => 
                           dp_ir_21_port, ZN => dp_id_stage_n8);
   dp_id_stage_U126 : INV_X1 port map( A => dp_ir_23_port, ZN => 
                           dp_id_stage_n11);
   dp_id_stage_U125 : INV_X1 port map( A => dp_ir_18_port, ZN => 
                           dp_id_stage_n16);
   dp_id_stage_U124 : INV_X1 port map( A => dp_id_stage_n7, ZN => 
                           dp_id_stage_p_addr_wRS1_1_port);
   dp_id_stage_U123 : INV_X1 port map( A => dp_ir_21_port, ZN => 
                           dp_id_stage_p_addr_wRS1_0_port);
   dp_id_stage_U122 : INV_X1 port map( A => dp_id_stage_n12, ZN => 
                           dp_id_stage_p_addr_wRS2_1_port);
   dp_id_stage_U121 : INV_X1 port map( A => dp_ir_16_port, ZN => 
                           dp_id_stage_p_addr_wRS2_0_port);
   dp_id_stage_U120 : INV_X1 port map( A => dp_rd_fwd_wb_i_2_port, ZN => 
                           dp_id_stage_n28);
   dp_id_stage_U119 : INV_X1 port map( A => dp_rd_fwd_wb_i_0_port, ZN => 
                           dp_id_stage_p_addr_wRD_0_port);
   dp_id_stage_U118 : OR3_X1 port map( A1 => dp_ir_20_port, A2 => dp_ir_19_port
                           , A3 => dp_ir_18_port, ZN => dp_id_stage_n18);
   dp_id_stage_U117 : OR3_X1 port map( A1 => dp_ir_17_port, A2 => dp_ir_16_port
                           , A3 => dp_id_stage_n18, ZN => dp_id_stage_n17);
   dp_id_stage_U116 : OR3_X1 port map( A1 => dp_ir_25_port, A2 => dp_ir_24_port
                           , A3 => dp_ir_23_port, ZN => dp_id_stage_n20);
   dp_id_stage_U115 : OR3_X1 port map( A1 => dp_ir_22_port, A2 => dp_ir_21_port
                           , A3 => dp_id_stage_n20, ZN => dp_id_stage_n19);
   dp_id_stage_U114 : INV_X1 port map( A => dp_id_stage_n24, ZN => 
                           dp_id_stage_p_addr_wRD_1_port);
   dp_id_stage_U113 : INV_X1 port map( A => imm_uns_i, ZN => dp_id_stage_n39);
   dp_id_stage_U112 : INV_X1 port map( A => dp_ir_22_port, ZN => 
                           dp_id_stage_n35);
   dp_id_stage_U111 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n35, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_22_port);
   dp_id_stage_U110 : AND2_X1 port map( A1 => dp_id_stage_out2_i_3_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_3_port);
   dp_id_stage_U109 : AND2_X1 port map( A1 => dp_id_stage_out2_i_4_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_4_port);
   dp_id_stage_U108 : AND2_X1 port map( A1 => dp_id_stage_out2_i_5_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_5_port);
   dp_id_stage_U107 : AND2_X1 port map( A1 => dp_id_stage_out2_i_6_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_6_port);
   dp_id_stage_U106 : AND2_X1 port map( A1 => dp_id_stage_out2_i_7_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_7_port);
   dp_id_stage_U105 : AND2_X1 port map( A1 => dp_id_stage_out2_i_8_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_8_port);
   dp_id_stage_U104 : AND2_X1 port map( A1 => dp_id_stage_out2_i_9_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_9_port);
   dp_id_stage_U103 : AND2_X1 port map( A1 => dp_id_stage_out2_i_10_port, A2 =>
                           dp_id_stage_n6, ZN => dp_rf_out2_id_o_10_port);
   dp_id_stage_U102 : AND2_X1 port map( A1 => dp_id_stage_out2_i_11_port, A2 =>
                           dp_id_stage_n6, ZN => dp_rf_out2_id_o_11_port);
   dp_id_stage_U101 : AND2_X1 port map( A1 => dp_id_stage_out2_i_12_port, A2 =>
                           dp_id_stage_n6, ZN => dp_rf_out2_id_o_12_port);
   dp_id_stage_U100 : AND2_X1 port map( A1 => dp_id_stage_out2_i_13_port, A2 =>
                           dp_id_stage_n6, ZN => dp_rf_out2_id_o_13_port);
   dp_id_stage_U99 : AND2_X1 port map( A1 => dp_id_stage_out2_i_14_port, A2 => 
                           dp_id_stage_n6, ZN => dp_rf_out2_id_o_14_port);
   dp_id_stage_U98 : AND2_X1 port map( A1 => dp_id_stage_out2_i_15_port, A2 => 
                           dp_id_stage_n6, ZN => dp_rf_out2_id_o_15_port);
   dp_id_stage_U97 : AND2_X1 port map( A1 => dp_id_stage_out2_i_16_port, A2 => 
                           dp_id_stage_n6, ZN => dp_rf_out2_id_o_16_port);
   dp_id_stage_U96 : AND2_X1 port map( A1 => dp_id_stage_out2_i_17_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_17_port);
   dp_id_stage_U95 : AND2_X1 port map( A1 => dp_id_stage_out2_i_18_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_18_port);
   dp_id_stage_U94 : AND2_X1 port map( A1 => dp_id_stage_out2_i_19_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_19_port);
   dp_id_stage_U93 : AND2_X1 port map( A1 => dp_id_stage_out2_i_20_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_20_port);
   dp_id_stage_U92 : AND2_X1 port map( A1 => dp_id_stage_out2_i_21_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_21_port);
   dp_id_stage_U91 : AND2_X1 port map( A1 => dp_id_stage_out1_i_0_port, A2 => 
                           dp_id_stage_n3, ZN => dp_rf_out1_id_o_0_port);
   dp_id_stage_U90 : AND2_X1 port map( A1 => dp_id_stage_out2_i_22_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_22_port);
   dp_id_stage_U89 : AND2_X1 port map( A1 => dp_id_stage_out2_i_23_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_23_port);
   dp_id_stage_U88 : AND2_X1 port map( A1 => dp_id_stage_out2_i_24_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_24_port);
   dp_id_stage_U87 : AND2_X1 port map( A1 => dp_id_stage_out2_i_25_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_25_port);
   dp_id_stage_U86 : AND2_X1 port map( A1 => dp_id_stage_out2_i_26_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_26_port);
   dp_id_stage_U85 : AND2_X1 port map( A1 => dp_id_stage_out2_i_27_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_27_port);
   dp_id_stage_U84 : AND2_X1 port map( A1 => dp_id_stage_out2_i_28_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_28_port);
   dp_id_stage_U83 : AND2_X1 port map( A1 => dp_id_stage_out2_i_29_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_29_port);
   dp_id_stage_U82 : AND2_X1 port map( A1 => dp_id_stage_out2_i_30_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_30_port);
   dp_id_stage_U81 : AND2_X1 port map( A1 => dp_id_stage_out2_i_31_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_31_port);
   dp_id_stage_U80 : AND2_X1 port map( A1 => dp_id_stage_out1_i_1_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_1_port);
   dp_id_stage_U79 : AND2_X1 port map( A1 => dp_id_stage_out1_i_2_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_2_port);
   dp_id_stage_U78 : AND2_X1 port map( A1 => dp_id_stage_out1_i_3_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_3_port);
   dp_id_stage_U77 : AND2_X1 port map( A1 => dp_id_stage_out1_i_4_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_4_port);
   dp_id_stage_U76 : AND2_X1 port map( A1 => dp_id_stage_out1_i_5_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_5_port);
   dp_id_stage_U75 : AND2_X1 port map( A1 => dp_id_stage_out1_i_6_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_6_port);
   dp_id_stage_U74 : AND2_X1 port map( A1 => dp_id_stage_out1_i_7_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_7_port);
   dp_id_stage_U73 : AND2_X1 port map( A1 => dp_id_stage_out1_i_8_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_8_port);
   dp_id_stage_U72 : AND2_X1 port map( A1 => dp_id_stage_out1_i_9_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_9_port);
   dp_id_stage_U71 : AND2_X1 port map( A1 => dp_id_stage_out1_i_10_port, A2 => 
                           dp_id_stage_n3, ZN => dp_rf_out1_id_o_10_port);
   dp_id_stage_U70 : AND2_X1 port map( A1 => dp_id_stage_out1_i_11_port, A2 => 
                           dp_id_stage_n3, ZN => dp_rf_out1_id_o_11_port);
   dp_id_stage_U69 : AND2_X1 port map( A1 => dp_id_stage_out1_i_12_port, A2 => 
                           dp_id_stage_n3, ZN => dp_rf_out1_id_o_12_port);
   dp_id_stage_U68 : AND2_X1 port map( A1 => dp_id_stage_out1_i_13_port, A2 => 
                           dp_id_stage_n3, ZN => dp_rf_out1_id_o_13_port);
   dp_id_stage_U67 : AND2_X1 port map( A1 => dp_id_stage_out1_i_14_port, A2 => 
                           dp_id_stage_n3, ZN => dp_rf_out1_id_o_14_port);
   dp_id_stage_U66 : AND2_X1 port map( A1 => dp_id_stage_out1_i_15_port, A2 => 
                           dp_id_stage_n3, ZN => dp_rf_out1_id_o_15_port);
   dp_id_stage_U65 : AND2_X1 port map( A1 => dp_id_stage_out1_i_16_port, A2 => 
                           dp_id_stage_n3, ZN => dp_rf_out1_id_o_16_port);
   dp_id_stage_U64 : AND2_X1 port map( A1 => dp_id_stage_out1_i_17_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_17_port);
   dp_id_stage_U63 : AND2_X1 port map( A1 => dp_id_stage_out1_i_18_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_18_port);
   dp_id_stage_U62 : AND2_X1 port map( A1 => dp_id_stage_out1_i_19_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_19_port);
   dp_id_stage_U61 : AND2_X1 port map( A1 => dp_id_stage_out1_i_20_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_20_port);
   dp_id_stage_U60 : AND2_X1 port map( A1 => dp_id_stage_out1_i_21_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_21_port);
   dp_id_stage_U59 : AND2_X1 port map( A1 => dp_id_stage_out1_i_22_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_22_port);
   dp_id_stage_U58 : AND2_X1 port map( A1 => dp_id_stage_out1_i_23_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_23_port);
   dp_id_stage_U57 : AND2_X1 port map( A1 => dp_id_stage_out1_i_24_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_24_port);
   dp_id_stage_U56 : INV_X1 port map( A => dp_ir_16_port, ZN => dp_id_stage_n29
                           );
   dp_id_stage_U55 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n29, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_16_port);
   dp_id_stage_U54 : INV_X1 port map( A => dp_ir_19_port, ZN => dp_id_stage_n32
                           );
   dp_id_stage_U53 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n32, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_19_port);
   dp_id_stage_U52 : INV_X1 port map( A => dp_ir_20_port, ZN => dp_id_stage_n33
                           );
   dp_id_stage_U51 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n33, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_20_port);
   dp_id_stage_U50 : INV_X1 port map( A => dp_ir_23_port, ZN => dp_id_stage_n36
                           );
   dp_id_stage_U49 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n36, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_23_port);
   dp_id_stage_U48 : INV_X1 port map( A => dp_ir_18_port, ZN => dp_id_stage_n31
                           );
   dp_id_stage_U47 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n31, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_18_port);
   dp_id_stage_U46 : INV_X1 port map( A => dp_ir_21_port, ZN => dp_id_stage_n34
                           );
   dp_id_stage_U45 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n34, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_21_port);
   dp_id_stage_U44 : INV_X1 port map( A => dp_ir_24_port, ZN => dp_id_stage_n37
                           );
   dp_id_stage_U43 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n37, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_24_port);
   dp_id_stage_U42 : INV_X1 port map( A => dp_ir_17_port, ZN => dp_id_stage_n30
                           );
   dp_id_stage_U41 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n30, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_17_port);
   dp_id_stage_U40 : AND2_X1 port map( A1 => dp_id_stage_out1_i_31_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_31_port);
   dp_id_stage_U39 : AND2_X1 port map( A1 => dp_id_stage_out1_i_26_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_26_port);
   dp_id_stage_U38 : AND2_X1 port map( A1 => dp_id_stage_out1_i_29_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_29_port);
   dp_id_stage_U37 : AND2_X1 port map( A1 => dp_id_stage_out1_i_25_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_25_port);
   dp_id_stage_U36 : AND2_X1 port map( A1 => dp_id_stage_out1_i_27_port, A2 => 
                           dp_id_stage_n2, ZN => dp_rf_out1_id_o_27_port);
   dp_id_stage_U35 : AND2_X1 port map( A1 => dp_id_stage_out1_i_28_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_28_port);
   dp_id_stage_U34 : AND2_X1 port map( A1 => dp_id_stage_out1_i_30_port, A2 => 
                           dp_id_stage_n1, ZN => dp_rf_out1_id_o_30_port);
   dp_id_stage_U33 : AND2_X1 port map( A1 => dp_id_stage_out2_i_0_port, A2 => 
                           dp_id_stage_n6, ZN => dp_rf_out2_id_o_0_port);
   dp_id_stage_U32 : AND2_X1 port map( A1 => dp_id_stage_out2_i_1_port, A2 => 
                           dp_id_stage_n5, ZN => dp_rf_out2_id_o_1_port);
   dp_id_stage_U31 : AND2_X1 port map( A1 => dp_id_stage_out2_i_2_port, A2 => 
                           dp_id_stage_n4, ZN => dp_rf_out2_id_o_2_port);
   dp_id_stage_U30 : AND2_X1 port map( A1 => dp_ir_14_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_14_port);
   dp_id_stage_U29 : AND2_X1 port map( A1 => dp_ir_1_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_1_port);
   dp_id_stage_U28 : AND2_X1 port map( A1 => dp_ir_2_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_2_port);
   dp_id_stage_U27 : AND2_X1 port map( A1 => dp_ir_4_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_4_port);
   dp_id_stage_U26 : AND2_X1 port map( A1 => dp_ir_5_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_5_port);
   dp_id_stage_U25 : AND2_X1 port map( A1 => dp_ir_7_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_7_port);
   dp_id_stage_U24 : AND2_X1 port map( A1 => dp_ir_11_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_11_port);
   dp_id_stage_U23 : AND2_X1 port map( A1 => dp_ir_0_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_0_port);
   dp_id_stage_U22 : AND2_X1 port map( A1 => dp_ir_3_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_3_port);
   dp_id_stage_U21 : AND2_X1 port map( A1 => dp_ir_6_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_6_port);
   dp_id_stage_U20 : AND2_X1 port map( A1 => dp_ir_8_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_8_port);
   dp_id_stage_U19 : AND2_X1 port map( A1 => dp_ir_9_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_9_port);
   dp_id_stage_U18 : AND2_X1 port map( A1 => dp_ir_10_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_10_port);
   dp_id_stage_U17 : AND2_X1 port map( A1 => dp_ir_12_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_12_port);
   dp_id_stage_U16 : AND2_X1 port map( A1 => dp_ir_13_port, A2 => 
                           dp_id_stage_n21, ZN => dp_imm_id_o_13_port);
   dp_id_stage_U15 : AND2_X1 port map( A1 => dp_id_stage_n21, A2 => 
                           dp_ir_15_port, ZN => dp_imm_id_o_15_port);
   dp_id_stage_U14 : NAND2_X1 port map( A1 => imm_isoff_i, A2 => 
                           dp_id_stage_n22, ZN => dp_id_stage_n21);
   dp_id_stage_U13 : NAND2_X1 port map( A1 => imm_isoff_i, A2 => 
                           dp_id_stage_n39, ZN => dp_id_stage_n22);
   dp_id_stage_U12 : INV_X1 port map( A => imm_isoff_i, ZN => dp_id_stage_n40);
   dp_id_stage_U11 : NAND3_X1 port map( A1 => dp_id_stage_n40, A2 => 
                           dp_id_stage_n39, A3 => dp_ir_15_port, ZN => 
                           dp_id_stage_n23);
   dp_id_stage_U10 : INV_X1 port map( A => dp_ir_25_port, ZN => dp_id_stage_n38
                           );
   dp_id_stage_U9 : OAI21_X1 port map( B1 => dp_id_stage_n22, B2 => 
                           dp_id_stage_n38, A => dp_id_stage_n23, ZN => 
                           dp_imm_id_o_31_port);
   dp_id_stage_U8 : BUF_X1 port map( A => dp_id_stage_n17, Z => dp_id_stage_n6)
                           ;
   dp_id_stage_U7 : BUF_X1 port map( A => dp_id_stage_n19, Z => dp_id_stage_n3)
                           ;
   dp_id_stage_U6 : BUF_X1 port map( A => dp_id_stage_n17, Z => dp_id_stage_n5)
                           ;
   dp_id_stage_U5 : BUF_X1 port map( A => dp_id_stage_n17, Z => dp_id_stage_n4)
                           ;
   dp_id_stage_U4 : BUF_X1 port map( A => dp_id_stage_n19, Z => dp_id_stage_n2)
                           ;
   dp_id_stage_U3 : BUF_X1 port map( A => dp_id_stage_n19, Z => dp_id_stage_n1)
                           ;
   dp_id_stage_regfile_ControlUnit_U46 : INV_X1 port map( A => rf_call_i, ZN =>
                           dp_id_stage_regfile_ControlUnit_n41);
   dp_id_stage_regfile_ControlUnit_U45 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_canrestore, A2 => rf_ret_i, ZN 
                           => dp_id_stage_regfile_ControlUnit_n24);
   dp_id_stage_regfile_ControlUnit_U44 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_cansave, A2 => 
                           dp_id_stage_regfile_ControlUnit_n41, B1 => rf_call_i
                           , B2 => dp_id_stage_regfile_ControlUnit_n24, ZN => 
                           dp_id_stage_regfile_ControlUnit_n23);
   dp_id_stage_regfile_ControlUnit_U43 : INV_X1 port map( A => 
                           dp_id_stage_regfile_end_sf, ZN => 
                           dp_id_stage_regfile_ControlUnit_n16);
   dp_id_stage_regfile_ControlUnit_U42 : AND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n13, A2 => 
                           dp_id_stage_regfile_ControlUnit_n12, A3 => 
                           dp_id_stage_regfile_ControlUnit_current_state_3_port
                           , ZN => dp_id_stage_regfile_cnt_swp);
   dp_id_stage_regfile_ControlUnit_U41 : NAND2_X1 port map( A1 => rf_call_i, A2
                           => dp_id_stage_regfile_ControlUnit_n6, ZN => 
                           dp_id_stage_regfile_ControlUnit_n19);
   dp_id_stage_regfile_ControlUnit_U40 : AOI21_X1 port map( B1 => 
                           dp_id_stage_regfile_ControlUnit_n17, B2 => 
                           dp_id_stage_regfile_ControlUnit_n19, A => RST, ZN =>
                           dp_id_stage_regfile_ControlUnit_next_state_1_port);
   dp_id_stage_regfile_ControlUnit_U39 : AOI21_X1 port map( B1 => 
                           dp_id_stage_regfile_ControlUnit_n17, B2 => 
                           dp_id_stage_regfile_ControlUnit_n18, A => RST, ZN =>
                           dp_id_stage_regfile_ControlUnit_next_state_2_port);
   dp_id_stage_regfile_ControlUnit_U38 : INV_X1 port map( A => 
                           dp_id_stage_regfile_ControlUnit_n26, ZN => 
                           dp_id_stage_regfile_ControlUnit_n15);
   dp_id_stage_regfile_ControlUnit_U37 : AOI21_X1 port map( B1 => 
                           dp_id_stage_regfile_ControlUnit_n6, B2 => 
                           dp_id_stage_regfile_ControlUnit_n23, A => 
                           dp_id_stage_regfile_rd_cu, ZN => 
                           dp_id_stage_regfile_ControlUnit_n22);
   dp_id_stage_regfile_ControlUnit_U36 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n15, A2 => 
                           dp_id_stage_regfile_ControlUnit_n12, B1 => 
                           dp_id_stage_regfile_ControlUnit_n25, B2 => 
                           dp_id_stage_regfile_ControlUnit_n14, ZN => 
                           dp_id_stage_regfile_ControlUnit_n21);
   dp_id_stage_regfile_ControlUnit_U35 : AOI21_X1 port map( B1 => 
                           dp_id_stage_regfile_ControlUnit_n21, B2 => 
                           dp_id_stage_regfile_ControlUnit_n22, A => RST, ZN =>
                           dp_id_stage_regfile_ControlUnit_next_state_0_port);
   dp_id_stage_regfile_ControlUnit_U34 : NOR3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n16, A2 => RST, A3 
                           => dp_id_stage_regfile_ControlUnit_n9, ZN => 
                           dp_id_stage_regfile_ControlUnit_next_state_3_port);
   dp_id_stage_regfile_ControlUnit_U33 : AOI21_X1 port map( B1 => 
                           dp_id_stage_regfile_ControlUnit_n13, B2 => 
                           dp_id_stage_regfile_ControlUnit_current_state_3_port
                           , A => dp_id_stage_regfile_ControlUnit_n27, ZN => 
                           dp_id_stage_regfile_ControlUnit_n26);
   dp_id_stage_regfile_ControlUnit_U32 : INV_X1 port map( A => 
                           dp_id_stage_regfile_ControlUnit_n29, ZN => 
                           dp_id_stage_regfile_wr_cu);
   dp_id_stage_regfile_ControlUnit_U31 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n14, A2 => 
                           dp_id_stage_regfile_ControlUnit_current_state_2_port
                           , ZN => dp_id_stage_regfile_ControlUnit_n40);
   dp_id_stage_regfile_ControlUnit_U30 : AND2_X2 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n1, A2 => 
                           dp_id_stage_regfile_ControlUnit_n13, ZN => 
                           dp_id_stage_regfile_ControlUnit_n25);
   dp_id_stage_regfile_ControlUnit_U29 : INV_X1 port map( A => 
                           dp_id_stage_regfile_up_dwn_cwp, ZN => 
                           dp_id_stage_regfile_ControlUnit_n5);
   dp_id_stage_regfile_ControlUnit_U28 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n35, A2 => 
                           dp_id_stage_regfile_ControlUnit_n5, ZN => 
                           dp_id_stage_regfile_up_dwn_rest);
   dp_id_stage_regfile_ControlUnit_U27 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n35, A2 => 
                           dp_id_stage_regfile_ControlUnit_n29, ZN => rf_fill_i
                           );
   dp_id_stage_regfile_ControlUnit_U26 : AND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n38, A2 => 
                           dp_id_stage_regfile_ControlUnit_n32, A3 => 
                           dp_id_stage_regfile_ControlUnit_n39, ZN => 
                           dp_id_stage_regfile_ControlUnit_n34);
   dp_id_stage_regfile_ControlUnit_U25 : NAND4_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n30, A2 => 
                           dp_id_stage_regfile_ControlUnit_n31, A3 => 
                           dp_id_stage_regfile_ControlUnit_n32, A4 => 
                           dp_id_stage_regfile_ControlUnit_n9, ZN => 
                           dp_id_stage_regfile_up_dwn_swp);
   dp_id_stage_regfile_ControlUnit_U24 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n37, A2 => 
                           dp_id_stage_regfile_ControlUnit_n28, ZN => 
                           rf_spill_i);
   dp_id_stage_regfile_ControlUnit_U23 : INV_X1 port map( A => rf_spill_i, ZN 
                           => dp_id_stage_regfile_ControlUnit_n4);
   dp_id_stage_regfile_ControlUnit_U22 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n30, A2 => 
                           dp_id_stage_regfile_ControlUnit_n4, ZN => 
                           dp_id_stage_regfile_sel_wp);
   dp_id_stage_regfile_ControlUnit_U21 : INV_X1 port map( A => 
                           dp_id_stage_regfile_ControlUnit_n28, ZN => 
                           dp_id_stage_regfile_rd_cu);
   dp_id_stage_regfile_ControlUnit_U20 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n40, A2 => 
                           dp_id_stage_regfile_ControlUnit_n25, ZN => 
                           dp_id_stage_regfile_ControlUnit_n38);
   dp_id_stage_regfile_ControlUnit_U19 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n36, A2 => 
                           dp_id_stage_regfile_ControlUnit_n33, ZN => 
                           dp_id_stage_regfile_cnt_save);
   dp_id_stage_regfile_ControlUnit_U18 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n37, A2 => 
                           dp_id_stage_regfile_ControlUnit_n35, ZN => 
                           dp_id_stage_regfile_ControlUnit_n20);
   dp_id_stage_regfile_ControlUnit_U17 : INV_X1 port map( A => 
                           dp_id_stage_regfile_ControlUnit_n32, ZN => 
                           dp_id_stage_regfile_rst_rf);
   dp_id_stage_regfile_ControlUnit_U16 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n40, A2 => 
                           dp_id_stage_regfile_ControlUnit_n27, ZN => 
                           dp_id_stage_regfile_ControlUnit_n37);
   dp_id_stage_regfile_ControlUnit_U15 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_cnt_swp, A2 => 
                           dp_id_stage_regfile_rf_enable, ZN => 
                           dp_id_stage_regfile_ControlUnit_n39);
   dp_id_stage_regfile_ControlUnit_U14 : AOI21_X1 port map( B1 => 
                           dp_id_stage_regfile_ControlUnit_n16, B2 => 
                           dp_id_stage_regfile_rf_enable, A => 
                           dp_id_stage_regfile_ControlUnit_n20, ZN => 
                           dp_id_stage_regfile_ControlUnit_n17);
   dp_id_stage_regfile_ControlUnit_U13 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n29, A2 => 
                           dp_id_stage_regfile_ControlUnit_n28, ZN => 
                           dp_id_stage_regfile_rf_enable);
   dp_id_stage_regfile_ControlUnit_U12 : INV_X1 port map( A => 
                           dp_id_stage_regfile_ControlUnit_n20, ZN => 
                           dp_id_stage_regfile_ControlUnit_n3);
   dp_id_stage_regfile_ControlUnit_U11 : INV_X1 port map( A => 
                           dp_id_stage_regfile_cnt_save, ZN => 
                           dp_id_stage_regfile_ControlUnit_n10);
   dp_id_stage_regfile_ControlUnit_U10 : INV_X1 port map( A => 
                           dp_id_stage_regfile_rf_enable, ZN => 
                           dp_id_stage_regfile_ControlUnit_n9);
   dp_id_stage_regfile_ControlUnit_U9 : INV_X1 port map( A => 
                           dp_id_stage_regfile_ControlUnit_n38, ZN => 
                           dp_id_stage_regfile_ControlUnit_n6);
   dp_id_stage_regfile_ControlUnit_U8 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n39, A2 => 
                           dp_id_stage_regfile_ControlUnit_n31, ZN => 
                           dp_id_stage_regfile_rst_swp);
   dp_id_stage_regfile_ControlUnit_U7 : NAND4_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n39, A2 => 
                           dp_id_stage_regfile_ControlUnit_n37, A3 => 
                           dp_id_stage_regfile_ControlUnit_n38, A4 => 
                           dp_id_stage_regfile_ControlUnit_n10, ZN => 
                           dp_id_stage_regfile_rst_spill_fill);
   dp_id_stage_regfile_ControlUnit_U6 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n3, A2 => 
                           dp_id_stage_regfile_ControlUnit_n10, ZN => 
                           dp_id_stage_regfile_cnt_cwp);
   dp_id_stage_regfile_ControlUnit_U5 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n6, A2 => 
                           dp_id_stage_regfile_cnt_cwp, ZN => 
                           dp_id_stage_regfile_ControlUnit_n31);
   dp_id_stage_regfile_ControlUnit_U4 : INV_X2 port map( A => 
                           dp_id_stage_regfile_ControlUnit_n31, ZN => 
                           dp_id_stage_regfile_cpu_work);
   dp_id_stage_regfile_ControlUnit_U3 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n13, A2 => 
                           dp_id_stage_regfile_ControlUnit_current_state_3_port
                           , ZN => dp_id_stage_regfile_ControlUnit_n27);
   dp_id_stage_regfile_ControlUnit_U56 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_current_state_2_port
                           , A2 => 
                           dp_id_stage_regfile_ControlUnit_current_state_0_port
                           , A3 => dp_id_stage_regfile_ControlUnit_n25, ZN => 
                           dp_id_stage_regfile_ControlUnit_n35);
   dp_id_stage_regfile_ControlUnit_U55 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n14, A2 => 
                           dp_id_stage_regfile_ControlUnit_n12, A3 => 
                           dp_id_stage_regfile_ControlUnit_n27, ZN => 
                           dp_id_stage_regfile_ControlUnit_n36);
   dp_id_stage_regfile_ControlUnit_U54 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_current_state_2_port
                           , A2 => dp_id_stage_regfile_ControlUnit_n14, A3 => 
                           dp_id_stage_regfile_ControlUnit_n25, ZN => 
                           dp_id_stage_regfile_ControlUnit_n33);
   dp_id_stage_regfile_ControlUnit_U53 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n27, A2 => 
                           dp_id_stage_regfile_ControlUnit_n14, A3 => 
                           dp_id_stage_regfile_ControlUnit_current_state_2_port
                           , ZN => dp_id_stage_regfile_ControlUnit_n29);
   dp_id_stage_regfile_ControlUnit_U52 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n14, A2 => 
                           dp_id_stage_regfile_ControlUnit_n12, A3 => 
                           dp_id_stage_regfile_ControlUnit_n25, ZN => 
                           dp_id_stage_regfile_ControlUnit_n32);
   dp_id_stage_regfile_ControlUnit_U51 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_current_state_0_port
                           , A2 => dp_id_stage_regfile_ControlUnit_n27, A3 => 
                           dp_id_stage_regfile_ControlUnit_current_state_2_port
                           , ZN => dp_id_stage_regfile_ControlUnit_n28);
   dp_id_stage_regfile_ControlUnit_U50 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n40, A2 => 
                           dp_id_stage_regfile_ControlUnit_n13, A3 => 
                           dp_id_stage_regfile_ControlUnit_current_state_3_port
                           , ZN => dp_id_stage_regfile_ControlUnit_n30);
   dp_id_stage_regfile_ControlUnit_U49 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n36, A2 => 
                           dp_id_stage_regfile_ControlUnit_n37, A3 => 
                           dp_id_stage_regfile_ControlUnit_n34, ZN => 
                           dp_id_stage_regfile_up_dwn_cwp);
   dp_id_stage_regfile_ControlUnit_U48 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n3, A2 => 
                           dp_id_stage_regfile_ControlUnit_n33, A3 => 
                           dp_id_stage_regfile_ControlUnit_n34, ZN => 
                           dp_id_stage_regfile_up_dwn_save);
   dp_id_stage_regfile_ControlUnit_U47 : NAND3_X1 port map( A1 => 
                           dp_id_stage_regfile_ControlUnit_n6, A2 => 
                           dp_id_stage_regfile_ControlUnit_n41, A3 => rf_ret_i,
                           ZN => dp_id_stage_regfile_ControlUnit_n18);
   dp_id_stage_regfile_ControlUnit_current_state_reg_3_inst : DFF_X1 port map( 
                           D => 
                           dp_id_stage_regfile_ControlUnit_next_state_3_port, 
                           CK => CLK, Q => 
                           dp_id_stage_regfile_ControlUnit_current_state_3_port
                           , QN => dp_id_stage_regfile_ControlUnit_n1);
   dp_id_stage_regfile_ControlUnit_current_state_reg_2_inst : DFF_X1 port map( 
                           D => 
                           dp_id_stage_regfile_ControlUnit_next_state_2_port, 
                           CK => CLK, Q => 
                           dp_id_stage_regfile_ControlUnit_current_state_2_port
                           , QN => dp_id_stage_regfile_ControlUnit_n12);
   dp_id_stage_regfile_ControlUnit_current_state_reg_1_inst : DFF_X1 port map( 
                           D => 
                           dp_id_stage_regfile_ControlUnit_next_state_1_port, 
                           CK => CLK, Q => n_1156, QN => 
                           dp_id_stage_regfile_ControlUnit_n13);
   dp_id_stage_regfile_ControlUnit_current_state_reg_0_inst : DFF_X1 port map( 
                           D => 
                           dp_id_stage_regfile_ControlUnit_next_state_0_port, 
                           CK => CLK, Q => 
                           dp_id_stage_regfile_ControlUnit_current_state_0_port
                           , QN => dp_id_stage_regfile_ControlUnit_n14);
   dp_id_stage_regfile_DataPath_U4 : AND3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_1_port, A2 
                           => dp_id_stage_regfile_DataPath_addr_sf_in_0_port, 
                           A3 => dp_id_stage_regfile_DataPath_addr_sf_in_2_port
                           , ZN => dp_id_stage_regfile_end_sf);
   dp_id_stage_regfile_DataPath_U3 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_CWP_0_port, ZN => 
                           dp_id_stage_regfile_DataPath_cwp_1_0_port);
   dp_id_stage_regfile_DataPath_Logic0_port <= '0';
   dp_id_stage_regfile_DataPath_Logic1_port <= '1';
   dp_id_stage_regfile_DataPath_Conv_RD1_U20 : AOI21_X1 port map( B1 => 
                           dp_id_stage_p_addr_wRS1_3_port, B2 => 
                           dp_id_stage_p_addr_wRS1_2_port, A => 
                           dp_id_stage_p_addr_wRS1_4_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_N1_port);
   dp_id_stage_regfile_DataPath_Conv_RD1_U19 : XNOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRS1_3_port, B => 
                           dp_id_stage_regfile_DataPath_CWP_0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n18);
   dp_id_stage_regfile_DataPath_Conv_RD1_U18 : XOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRS1_3_port, B => 
                           dp_id_stage_p_addr_wRS1_2_port, Z => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n4);
   dp_id_stage_regfile_DataPath_Conv_RD1_U17 : AND2_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRS1_3_port, A2 => 
                           dp_id_stage_p_addr_wRS1_2_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n3);
   dp_id_stage_regfile_DataPath_Conv_RD1_U16 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_N5, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n8, B1 => 
                           dp_id_stage_p_addr_wRS1_2_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_N1_port, ZN =>
                           dp_id_stage_regfile_DataPath_Conv_RD1_n20);
   dp_id_stage_regfile_DataPath_Conv_RD1_U15 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n20, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_2_port);
   dp_id_stage_regfile_DataPath_Conv_RD1_U14 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n1, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n8, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_4_port);
   dp_id_stage_regfile_DataPath_Conv_RD1_U13 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n2, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n8, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_5_port);
   dp_id_stage_regfile_DataPath_Conv_RD1_U12 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n4, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n8, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n19);
   dp_id_stage_regfile_DataPath_Conv_RD1_U11 : OAI21_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n18, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n8, A => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n19, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_3_port);
   dp_id_stage_regfile_DataPath_Conv_RD1_U10 : AOI22_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRS1_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n8, B1 => 
                           dp_id_stage_p_addr_wRS1_1_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_N1_port, ZN =>
                           dp_id_stage_regfile_DataPath_Conv_RD1_n21);
   dp_id_stage_regfile_DataPath_Conv_RD1_U9 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n21, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_1_port);
   dp_id_stage_regfile_DataPath_Conv_RD1_U8 : AOI22_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRS1_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n8, B1 => 
                           dp_id_stage_p_addr_wRS1_0_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_N1_port, ZN =>
                           dp_id_stage_regfile_DataPath_Conv_RD1_n22);
   dp_id_stage_regfile_DataPath_Conv_RD1_U7 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n22, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_0_port);
   dp_id_stage_regfile_DataPath_Conv_RD1_U6 : INV_X1 port map( A => 
                           dp_id_stage_p_addr_wRS1_2_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_N5);
   dp_id_stage_regfile_DataPath_Conv_RD1_U5 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_N1_port, ZN =>
                           dp_id_stage_regfile_DataPath_Conv_RD1_n8);
   dp_id_stage_regfile_DataPath_Conv_RD1_U4 : AND2_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRS1_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n3, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n2);
   dp_id_stage_regfile_DataPath_Conv_RD1_U3 : XOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRS1_4_port, B => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n3, Z => 
                           dp_id_stage_regfile_DataPath_Conv_RD1_n1);
   dp_id_stage_regfile_DataPath_Conv_RD2_U20 : AOI21_X1 port map( B1 => 
                           dp_id_stage_p_addr_wRS2_3_port, B2 => 
                           dp_id_stage_p_addr_wRS2_2_port, A => 
                           dp_id_stage_p_addr_wRS2_4_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_N1_port);
   dp_id_stage_regfile_DataPath_Conv_RD2_U19 : AOI22_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRS2_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n8, B1 => 
                           dp_id_stage_p_addr_wRS2_1_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_N1_port, ZN =>
                           dp_id_stage_regfile_DataPath_Conv_RD2_n10);
   dp_id_stage_regfile_DataPath_Conv_RD2_U18 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n10, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_1_port);
   dp_id_stage_regfile_DataPath_Conv_RD2_U17 : AOI22_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRS2_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n8, B1 => 
                           dp_id_stage_p_addr_wRS2_0_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_N1_port, ZN =>
                           dp_id_stage_regfile_DataPath_Conv_RD2_n9);
   dp_id_stage_regfile_DataPath_Conv_RD2_U16 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n9, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_0_port);
   dp_id_stage_regfile_DataPath_Conv_RD2_U15 : XNOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRS2_3_port, B => 
                           dp_id_stage_regfile_DataPath_CWP_0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n13);
   dp_id_stage_regfile_DataPath_Conv_RD2_U14 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n1, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n8, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n12);
   dp_id_stage_regfile_DataPath_Conv_RD2_U13 : OAI21_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n13, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n8, A => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n12, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_3_port);
   dp_id_stage_regfile_DataPath_Conv_RD2_U12 : AND2_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRS2_3_port, A2 => 
                           dp_id_stage_p_addr_wRS2_2_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n4);
   dp_id_stage_regfile_DataPath_Conv_RD2_U11 : AND2_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRS2_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n4, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n3);
   dp_id_stage_regfile_DataPath_Conv_RD2_U10 : XOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRS2_4_port, B => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n4, Z => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n2);
   dp_id_stage_regfile_DataPath_Conv_RD2_U9 : INV_X1 port map( A => 
                           dp_id_stage_p_addr_wRS2_2_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_N5);
   dp_id_stage_regfile_DataPath_Conv_RD2_U8 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_N5, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n8, B1 => 
                           dp_id_stage_p_addr_wRS2_2_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_N1_port, ZN =>
                           dp_id_stage_regfile_DataPath_Conv_RD2_n11);
   dp_id_stage_regfile_DataPath_Conv_RD2_U7 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n11, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_2_port);
   dp_id_stage_regfile_DataPath_Conv_RD2_U6 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_N1_port, ZN =>
                           dp_id_stage_regfile_DataPath_Conv_RD2_n8);
   dp_id_stage_regfile_DataPath_Conv_RD2_U5 : XOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRS2_3_port, B => 
                           dp_id_stage_p_addr_wRS2_2_port, Z => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n1);
   dp_id_stage_regfile_DataPath_Conv_RD2_U4 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n3, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n8, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_5_port);
   dp_id_stage_regfile_DataPath_Conv_RD2_U3 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n2, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_RD2_n8, ZN => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_4_port);
   dp_id_stage_regfile_DataPath_Conv_W_U20 : AOI21_X1 port map( B1 => 
                           dp_id_stage_p_addr_wRD_3_port, B2 => 
                           dp_id_stage_p_addr_wRD_2_port, A => 
                           dp_id_stage_p_addr_wRD_4_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_N1_port);
   dp_id_stage_regfile_DataPath_Conv_W_U19 : XNOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRD_3_port, B => 
                           dp_id_stage_regfile_DataPath_CWP_0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_n13);
   dp_id_stage_regfile_DataPath_Conv_W_U18 : OAI21_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n13, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n8, A => 
                           dp_id_stage_regfile_DataPath_Conv_W_n12, ZN => 
                           dp_id_stage_regfile_DataPath_addr_w_p_3_port);
   dp_id_stage_regfile_DataPath_Conv_W_U17 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n3, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n8, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_n12);
   dp_id_stage_regfile_DataPath_Conv_W_U16 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n2, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n8, ZN => 
                           dp_id_stage_regfile_DataPath_addr_w_p_5_port);
   dp_id_stage_regfile_DataPath_Conv_W_U15 : AND2_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRD_3_port, A2 => 
                           dp_id_stage_p_addr_wRD_2_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_n4);
   dp_id_stage_regfile_DataPath_Conv_W_U14 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n1, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n8, ZN => 
                           dp_id_stage_regfile_DataPath_addr_w_p_4_port);
   dp_id_stage_regfile_DataPath_Conv_W_U13 : AOI22_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRD_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n8, B1 => 
                           dp_id_stage_p_addr_wRD_1_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_N1_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_n10);
   dp_id_stage_regfile_DataPath_Conv_W_U12 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_W_n10, ZN => 
                           dp_id_stage_regfile_DataPath_addr_w_p_1_port);
   dp_id_stage_regfile_DataPath_Conv_W_U11 : AOI22_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRD_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n8, B1 => 
                           dp_id_stage_p_addr_wRD_0_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_N1_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_n9);
   dp_id_stage_regfile_DataPath_Conv_W_U10 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_W_n9, ZN => 
                           dp_id_stage_regfile_DataPath_addr_w_p_0_port);
   dp_id_stage_regfile_DataPath_Conv_W_U9 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Conv_W_N5, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n8, B1 => 
                           dp_id_stage_p_addr_wRD_2_port, B2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_N1_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_n11);
   dp_id_stage_regfile_DataPath_Conv_W_U8 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_W_n11, ZN => 
                           dp_id_stage_regfile_DataPath_addr_w_p_2_port);
   dp_id_stage_regfile_DataPath_Conv_W_U7 : INV_X1 port map( A => 
                           dp_id_stage_p_addr_wRD_2_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_N5);
   dp_id_stage_regfile_DataPath_Conv_W_U6 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Conv_W_N1_port, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_n8);
   dp_id_stage_regfile_DataPath_Conv_W_U5 : XOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRD_3_port, B => 
                           dp_id_stage_p_addr_wRD_2_port, Z => 
                           dp_id_stage_regfile_DataPath_Conv_W_n3);
   dp_id_stage_regfile_DataPath_Conv_W_U4 : AND2_X1 port map( A1 => 
                           dp_id_stage_p_addr_wRD_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Conv_W_n4, ZN => 
                           dp_id_stage_regfile_DataPath_Conv_W_n2);
   dp_id_stage_regfile_DataPath_Conv_W_U3 : XOR2_X1 port map( A => 
                           dp_id_stage_p_addr_wRD_4_port, B => 
                           dp_id_stage_regfile_DataPath_Conv_W_n4, Z => 
                           dp_id_stage_regfile_DataPath_Conv_W_n1);
   dp_id_stage_regfile_DataPath_SF_converter_U20 : AOI21_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, B2 => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_2_port, A =>
                           dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_SF_converter_N1_port);
   dp_id_stage_regfile_DataPath_SF_converter_U19 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, A2 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n2, ZN => 
                           dp_id_stage_regfile_DataPath_SF_converter_n4);
   dp_id_stage_regfile_DataPath_SF_converter_U18 : XOR2_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Logic0_port, B => 
                           dp_id_stage_regfile_DataPath_SF_converter_n2, Z => 
                           dp_id_stage_regfile_DataPath_SF_converter_n3);
   dp_id_stage_regfile_DataPath_SF_converter_U17 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, A2 => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_2_port, ZN 
                           => dp_id_stage_regfile_DataPath_SF_converter_n2);
   dp_id_stage_regfile_DataPath_SF_converter_U16 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_2_port, ZN 
                           => dp_id_stage_regfile_DataPath_SF_converter_N5_port
                           );
   dp_id_stage_regfile_DataPath_SF_converter_U15 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_SF_converter_N5_port, 
                           A2 => dp_id_stage_regfile_DataPath_SF_converter_n10,
                           B1 => dp_id_stage_regfile_DataPath_addr_sf_in_2_port
                           , B2 => 
                           dp_id_stage_regfile_DataPath_SF_converter_N1_port, 
                           ZN => dp_id_stage_regfile_DataPath_SF_converter_n7);
   dp_id_stage_regfile_DataPath_SF_converter_U14 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_SF_converter_n7, ZN => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_2_port)
                           ;
   dp_id_stage_regfile_DataPath_SF_converter_U13 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_1_port, A2 
                           => dp_id_stage_regfile_DataPath_SF_converter_n10, B1
                           => dp_id_stage_regfile_DataPath_addr_sf_in_1_port, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_SF_converter_N1_port, 
                           ZN => dp_id_stage_regfile_DataPath_SF_converter_n6);
   dp_id_stage_regfile_DataPath_SF_converter_U12 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_SF_converter_n6, ZN => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_1_port)
                           ;
   dp_id_stage_regfile_DataPath_SF_converter_U11 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_0_port, A2 
                           => dp_id_stage_regfile_DataPath_SF_converter_n10, B1
                           => dp_id_stage_regfile_DataPath_addr_sf_in_0_port, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_SF_converter_N1_port, 
                           ZN => dp_id_stage_regfile_DataPath_SF_converter_n5);
   dp_id_stage_regfile_DataPath_SF_converter_U10 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_SF_converter_n5, ZN => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_0_port)
                           ;
   dp_id_stage_regfile_DataPath_SF_converter_U9 : XNOR2_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Logic0_port, B => 
                           dp_id_stage_regfile_DataPath_sf_wp_0_port, ZN => 
                           dp_id_stage_regfile_DataPath_SF_converter_n9);
   dp_id_stage_regfile_DataPath_SF_converter_U8 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n1, A2 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n10, ZN =>
                           dp_id_stage_regfile_DataPath_SF_converter_n8);
   dp_id_stage_regfile_DataPath_SF_converter_U7 : OAI21_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n9, B2 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n10, A => 
                           dp_id_stage_regfile_DataPath_SF_converter_n8, ZN => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_3_port)
                           ;
   dp_id_stage_regfile_DataPath_SF_converter_U6 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_SF_converter_N1_port, 
                           ZN => dp_id_stage_regfile_DataPath_SF_converter_n10)
                           ;
   dp_id_stage_regfile_DataPath_SF_converter_U5 : XOR2_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Logic0_port, B => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_2_port, Z =>
                           dp_id_stage_regfile_DataPath_SF_converter_n1);
   dp_id_stage_regfile_DataPath_SF_converter_U4 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n3, A2 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n10, ZN =>
                           dp_id_stage_regfile_DataPath_spill_fill_addr_4_port)
                           ;
   dp_id_stage_regfile_DataPath_SF_converter_U3 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n4, A2 => 
                           dp_id_stage_regfile_DataPath_SF_converter_n10, ZN =>
                           dp_id_stage_regfile_DataPath_spill_fill_addr_5_port)
                           ;
   dp_id_stage_regfile_DataPath_Cwp_counter_U6 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n2);
   dp_id_stage_regfile_DataPath_Cwp_counter_U5 : INV_X1 port map( A => 
                           dp_id_stage_regfile_rst_swp, ZN => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n4);
   dp_id_stage_regfile_DataPath_Cwp_counter_U4 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n3, A2 => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n2, B1 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, B2 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n1);
   dp_id_stage_regfile_DataPath_Cwp_counter_U3 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n1, A2 => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n4, ZN => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n5);
   dp_id_stage_regfile_DataPath_Cwp_counter_U7 : XOR2_X1 port map( A => 
                           dp_id_stage_regfile_cnt_cwp, B => 
                           dp_id_stage_regfile_DataPath_CWP_0_port, Z => 
                           dp_id_stage_regfile_DataPath_Cwp_counter_n3);
   dp_id_stage_regfile_DataPath_Cwp_counter_Q_reg_0_inst : DFF_X1 port map( D 
                           => dp_id_stage_regfile_DataPath_Cwp_counter_n5, CK 
                           => CLK, Q => dp_id_stage_regfile_DataPath_CWP_0_port
                           , QN => n_1157);
   dp_id_stage_regfile_DataPath_Swp_counter_U6 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Swp_counter_n2);
   dp_id_stage_regfile_DataPath_Swp_counter_U5 : INV_X1 port map( A => 
                           dp_id_stage_regfile_rst_swp, ZN => 
                           dp_id_stage_regfile_DataPath_Swp_counter_n4);
   dp_id_stage_regfile_DataPath_Swp_counter_U4 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Swp_counter_n7, A2 => 
                           dp_id_stage_regfile_DataPath_Swp_counter_n2, B1 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, B2 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Swp_counter_n8);
   dp_id_stage_regfile_DataPath_Swp_counter_U3 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Swp_counter_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Swp_counter_n4, ZN => 
                           dp_id_stage_regfile_DataPath_Swp_counter_n6);
   dp_id_stage_regfile_DataPath_Swp_counter_U7 : XOR2_X1 port map( A => 
                           dp_id_stage_regfile_cnt_swp, B => 
                           dp_id_stage_regfile_DataPath_Swp_counter_Q_0_port, Z
                           => dp_id_stage_regfile_DataPath_Swp_counter_n7);
   dp_id_stage_regfile_DataPath_Swp_counter_Q_reg_0_inst : DFF_X1 port map( D 
                           => dp_id_stage_regfile_DataPath_Swp_counter_n6, CK 
                           => CLK, Q => 
                           dp_id_stage_regfile_DataPath_Swp_counter_Q_0_port, 
                           QN => n_1158);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U18 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n4);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U17 : XNOR2_X1 port map( A 
                           => dp_id_stage_regfile_DataPath_Logic1_port, B => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n11,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n10)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U16 : AOI22_X1 port map( A1 
                           => dp_id_stage_regfile_DataPath_addr_sf_in_1_port, 
                           A2 => dp_id_stage_regfile_DataPath_addr_sf_in_0_port
                           , B1 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n11,
                           B2 => dp_id_stage_regfile_DataPath_Logic1_port, ZN 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n9);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U15 : XNOR2_X1 port map( A 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n9, 
                           B => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n10,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n7);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U14 : AOI22_X1 port map( A1 
                           => dp_id_stage_regfile_DataPath_Logic0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, B1 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n1, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n4, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n18)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U13 : OR2_X1 port map( A1 =>
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n14,
                           A2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n18,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n17)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U12 : OAI22_X1 port map( A1 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n1, 
                           A2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n12,
                           B1 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n16,
                           B2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n17,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n21)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U11 : AOI22_X1 port map( A1 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n10,
                           A2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n4, 
                           B1 => dp_id_stage_regfile_DataPath_Logic0_port, B2 
                           => dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n15)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U10 : OR2_X1 port map( A1 =>
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n14,
                           A2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n15,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n13)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U9 : OAI22_X1 port map( A1 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n3, 
                           A2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n12,
                           B1 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n16,
                           B2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n13,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n20)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U8 : OAI21_X1 port map( B1 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n7, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n2, 
                           A => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n8, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n6);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U7 : AOI22_X1 port map( A1 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n6, 
                           A2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n4, 
                           B1 => dp_id_stage_regfile_DataPath_Logic0_port, B2 
                           => dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n5);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U6 : OAI22_X1 port map( A1 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n2, 
                           A2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n12,
                           B1 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n5, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n16,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n19)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U5 : NOR3_X1 port map( A1 =>
                           dp_id_stage_regfile_rf_enable, A2 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, A3 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n16,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n14)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U4 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n14,
                           ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n12)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U3 : INV_X1 port map( A => 
                           dp_id_stage_regfile_rst_spill_fill, ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n16)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U23 : XOR2_X1 port map( A =>
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n3, 
                           B => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n1, 
                           Z => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n11)
                           ;
   dp_id_stage_regfile_DataPath_Spill_fill_counter_U22 : NAND3_X1 port map( A1 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n7, 
                           A2 => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n2, 
                           A3 => dp_id_stage_regfile_rf_enable, ZN => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n8);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_Q_reg_2_inst : DFF_X1 port 
                           map( D => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n19,
                           CK => CLK, Q => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_2_port, QN 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n2);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_Q_reg_1_inst : DFF_X1 port 
                           map( D => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n20,
                           CK => CLK, Q => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_1_port, QN 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n3);
   dp_id_stage_regfile_DataPath_Spill_fill_counter_Q_reg_0_inst : DFF_X1 port 
                           map( D => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n21,
                           CK => CLK, Q => 
                           dp_id_stage_regfile_DataPath_addr_sf_in_0_port, QN 
                           => 
                           dp_id_stage_regfile_DataPath_Spill_fill_counter_n1);
   dp_id_stage_regfile_DataPath_CANSAVE_counter_U6 : INV_X1 port map( A => 
                           dp_id_stage_regfile_rst_rf, ZN => 
                           dp_id_stage_regfile_DataPath_CANSAVE_counter_n4);
   dp_id_stage_regfile_DataPath_CANSAVE_counter_U5 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_CANSAVE_counter_n7, A2 
                           => dp_id_stage_regfile_DataPath_CANSAVE_counter_n4, 
                           B1 => dp_id_stage_regfile_rst_rf, B2 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_CANSAVE_counter_n8);
   dp_id_stage_regfile_DataPath_CANSAVE_counter_U4 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Logic1_port, ZN => 
                           dp_id_stage_regfile_DataPath_CANSAVE_counter_n2);
   dp_id_stage_regfile_DataPath_CANSAVE_counter_U3 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_CANSAVE_counter_n8, A2 
                           => dp_id_stage_regfile_DataPath_CANSAVE_counter_n2, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_CANSAVE_counter_n6);
   dp_id_stage_regfile_DataPath_CANSAVE_counter_U7 : XOR2_X1 port map( A => 
                           dp_id_stage_regfile_cnt_save, B => 
                           dp_id_stage_regfile_cansave, Z => 
                           dp_id_stage_regfile_DataPath_CANSAVE_counter_n7);
   dp_id_stage_regfile_DataPath_CANSAVE_counter_Q_reg_0_inst : DFF_X1 port map(
                           D => dp_id_stage_regfile_DataPath_CANSAVE_counter_n6
                           , CK => CLK, Q => dp_id_stage_regfile_cansave, QN =>
                           n_1159);
   dp_id_stage_regfile_DataPath_CANRESTORE_counter_U6 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n2);
   dp_id_stage_regfile_DataPath_CANRESTORE_counter_U5 : INV_X1 port map( A => 
                           dp_id_stage_regfile_rst_swp, ZN => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n4);
   dp_id_stage_regfile_DataPath_CANRESTORE_counter_U4 : AOI22_X1 port map( A1 
                           => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n7, 
                           A2 => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n2, 
                           B1 => dp_id_stage_regfile_DataPath_Logic0_port, B2 
                           => dp_id_stage_regfile_DataPath_Logic0_port, ZN => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n8);
   dp_id_stage_regfile_DataPath_CANRESTORE_counter_U3 : NOR2_X1 port map( A1 =>
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n8, 
                           A2 => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n4, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n6);
   dp_id_stage_regfile_DataPath_CANRESTORE_counter_U7 : XOR2_X1 port map( A => 
                           dp_id_stage_regfile_cnt_save, B => 
                           dp_id_stage_regfile_canrestore, Z => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n7);
   dp_id_stage_regfile_DataPath_CANRESTORE_counter_Q_reg_0_inst : DFF_X1 port 
                           map( D => 
                           dp_id_stage_regfile_DataPath_CANRESTORE_counter_n6, 
                           CK => CLK, Q => dp_id_stage_regfile_canrestore, QN 
                           => n_1160);
   dp_id_stage_regfile_DataPath_Mux_rd_U13 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_2_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_rd_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_2_port, B2 
                           => dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n11);
   dp_id_stage_regfile_DataPath_Mux_rd_U12 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n11, ZN => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_2_port);
   dp_id_stage_regfile_DataPath_Mux_rd_U11 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_4_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_rd_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_4_port, B2 
                           => dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n9);
   dp_id_stage_regfile_DataPath_Mux_rd_U10 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n9, ZN => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_4_port);
   dp_id_stage_regfile_DataPath_Mux_rd_U9 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_5_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_rd_n1, B1 => 
                           dp_id_stage_regfile_cpu_work, B2 => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_5_port, ZN 
                           => dp_id_stage_regfile_DataPath_Mux_rd_n8);
   dp_id_stage_regfile_DataPath_Mux_rd_U8 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n8, ZN => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_5_port);
   dp_id_stage_regfile_DataPath_Mux_rd_U7 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_3_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_rd_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_3_port, B2 
                           => dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n10);
   dp_id_stage_regfile_DataPath_Mux_rd_U6 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n10, ZN => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_3_port);
   dp_id_stage_regfile_DataPath_Mux_rd_U5 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_1_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_rd_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_1_port, B2 
                           => dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n12);
   dp_id_stage_regfile_DataPath_Mux_rd_U4 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n12, ZN => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_1_port);
   dp_id_stage_regfile_DataPath_Mux_rd_U3 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_0_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_rd_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_rd1_p_0_port, B2 
                           => dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n13);
   dp_id_stage_regfile_DataPath_Mux_rd_U2 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n13, ZN => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_0_port);
   dp_id_stage_regfile_DataPath_Mux_rd_U1 : INV_X1 port map( A => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd_n1);
   dp_id_stage_regfile_DataPath_Mux_wr_U13 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_3_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_wr_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_w_p_3_port, B2 => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n5);
   dp_id_stage_regfile_DataPath_Mux_wr_U12 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n5, ZN => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_3_port);
   dp_id_stage_regfile_DataPath_Mux_wr_U11 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_5_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_wr_n1, B1 => 
                           dp_id_stage_regfile_cpu_work, B2 => 
                           dp_id_stage_regfile_DataPath_addr_w_p_5_port, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n7);
   dp_id_stage_regfile_DataPath_Mux_wr_U10 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n7, ZN => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_5_port);
   dp_id_stage_regfile_DataPath_Mux_wr_U9 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_4_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_wr_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_w_p_4_port, B2 => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n6);
   dp_id_stage_regfile_DataPath_Mux_wr_U8 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n6, ZN => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_4_port);
   dp_id_stage_regfile_DataPath_Mux_wr_U7 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_1_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_wr_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_w_p_1_port, B2 => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n3);
   dp_id_stage_regfile_DataPath_Mux_wr_U6 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_0_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_wr_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_w_p_0_port, B2 => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n2);
   dp_id_stage_regfile_DataPath_Mux_wr_U5 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_spill_fill_addr_2_port,
                           A2 => dp_id_stage_regfile_DataPath_Mux_wr_n1, B1 => 
                           dp_id_stage_regfile_DataPath_addr_w_p_2_port, B2 => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n4);
   dp_id_stage_regfile_DataPath_Mux_wr_U4 : INV_X1 port map( A => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n1);
   dp_id_stage_regfile_DataPath_Mux_wr_U3 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n4, ZN => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_2_port);
   dp_id_stage_regfile_DataPath_Mux_wr_U2 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n3, ZN => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_1_port);
   dp_id_stage_regfile_DataPath_Mux_wr_U1 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_wr_n2, ZN => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_0_port);
   dp_id_stage_regfile_DataPath_Mux_sf_U3 : INV_X1 port map( A => 
                           dp_id_stage_regfile_sel_wp, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_sf_n1);
   dp_id_stage_regfile_DataPath_Mux_sf_U2 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_CWP_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Mux_sf_n1, B1 => 
                           dp_id_stage_regfile_sel_wp, B2 => 
                           dp_id_stage_regfile_DataPath_cwp_1_0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_sf_n3);
   dp_id_stage_regfile_DataPath_Mux_sf_U1 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_sf_n3, ZN => 
                           dp_id_stage_regfile_DataPath_sf_wp_0_port);
   dp_id_stage_regfile_DataPath_Mux_rd1_control_U3 : INV_X1 port map( A => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd1_control_n2);
   dp_id_stage_regfile_DataPath_Mux_rd1_control_U2 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_rd_cu, A2 => 
                           dp_id_stage_regfile_DataPath_Mux_rd1_control_n2, B1 
                           => dp_id_stage_regfile_cpu_work, B2 => rf_rs1_en_i, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd1_control_n3);
   dp_id_stage_regfile_DataPath_Mux_rd1_control_U1 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_rd1_control_n3, ZN 
                           => dp_id_stage_regfile_DataPath_mux_rd1_control_out)
                           ;
   dp_id_stage_regfile_DataPath_Mux_rd2_control_U3 : INV_X1 port map( A => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd2_control_n2);
   dp_id_stage_regfile_DataPath_Mux_rd2_control_U2 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Logic0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Mux_rd2_control_n2, B1 
                           => dp_id_stage_regfile_cpu_work, B2 => rf_rs2_en_i, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Mux_rd2_control_n4);
   dp_id_stage_regfile_DataPath_Mux_rd2_control_U1 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_rd2_control_n4, ZN 
                           => dp_id_stage_regfile_DataPath_mux_rd2_control_out)
                           ;
   dp_id_stage_regfile_DataPath_Mux_wr_control_U3 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_wr_cu, A2 => 
                           dp_id_stage_regfile_DataPath_Mux_wr_control_n2, B1 
                           => dp_id_stage_regfile_cpu_work, B2 => rf_we_i, ZN 
                           => dp_id_stage_regfile_DataPath_Mux_wr_control_n4);
   dp_id_stage_regfile_DataPath_Mux_wr_control_U2 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_wr_control_n4, ZN 
                           => dp_id_stage_regfile_DataPath_mux_wr_control_out);
   dp_id_stage_regfile_DataPath_Mux_wr_control_U1 : INV_X1 port map( A => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_wr_control_n2);
   dp_id_stage_regfile_DataPath_Mux_en_control_U3 : INV_X1 port map( A => 
                           dp_id_stage_regfile_cpu_work, ZN => 
                           dp_id_stage_regfile_DataPath_Mux_en_control_n2);
   dp_id_stage_regfile_DataPath_Mux_en_control_U2 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_rf_enable, A2 => 
                           dp_id_stage_regfile_DataPath_Mux_en_control_n2, B1 
                           => dp_id_stage_regfile_cpu_work, B2 => rf_en_i, ZN 
                           => dp_id_stage_regfile_DataPath_Mux_en_control_n4);
   dp_id_stage_regfile_DataPath_Mux_en_control_U1 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Mux_en_control_n4, ZN 
                           => dp_id_stage_regfile_DataPath_mux_en_control_out);
   dp_id_stage_regfile_DataPath_Physical_RF_U3825 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4227, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4220);
   dp_id_stage_regfile_DataPath_Physical_RF_U3824 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4217, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4210);
   dp_id_stage_regfile_DataPath_Physical_RF_U3823 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4207, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4200);
   dp_id_stage_regfile_DataPath_Physical_RF_U3822 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4144, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4137);
   dp_id_stage_regfile_DataPath_Physical_RF_U3821 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4134, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4127);
   dp_id_stage_regfile_DataPath_Physical_RF_U3820 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4124, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4117);
   dp_id_stage_regfile_DataPath_Physical_RF_U3819 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4114, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4107);
   dp_id_stage_regfile_DataPath_Physical_RF_U3818 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4042, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4035);
   dp_id_stage_regfile_DataPath_Physical_RF_U3817 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4032, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4025);
   dp_id_stage_regfile_DataPath_Physical_RF_U3816 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3982, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3975);
   dp_id_stage_regfile_DataPath_Physical_RF_U3815 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3950, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3943);
   dp_id_stage_regfile_DataPath_Physical_RF_U3814 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3900, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3893);
   dp_id_stage_regfile_DataPath_Physical_RF_U3813 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3890, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3883);
   dp_id_stage_regfile_DataPath_Physical_RF_U3812 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1189, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1188);
   dp_id_stage_regfile_DataPath_Physical_RF_U3811 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1189, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187);
   dp_id_stage_regfile_DataPath_Physical_RF_U3810 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1189, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186);
   dp_id_stage_regfile_DataPath_Physical_RF_U3809 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1189, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1185);
   dp_id_stage_regfile_DataPath_Physical_RF_U3808 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1200, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184);
   dp_id_stage_regfile_DataPath_Physical_RF_U3807 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1200, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183);
   dp_id_stage_regfile_DataPath_Physical_RF_U3806 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1200, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182);
   dp_id_stage_regfile_DataPath_Physical_RF_U3805 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1200, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181);
   dp_id_stage_regfile_DataPath_Physical_RF_U3804 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1200, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180);
   dp_id_stage_regfile_DataPath_Physical_RF_U3803 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1200, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1179);
   dp_id_stage_regfile_DataPath_Physical_RF_U3802 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1202, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178);
   dp_id_stage_regfile_DataPath_Physical_RF_U3801 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1202, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177);
   dp_id_stage_regfile_DataPath_Physical_RF_U3800 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1202, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1176);
   dp_id_stage_regfile_DataPath_Physical_RF_U3799 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1202, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175);
   dp_id_stage_regfile_DataPath_Physical_RF_U3798 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1202, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174);
   dp_id_stage_regfile_DataPath_Physical_RF_U3797 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_rd2_control_out, A2
                           => dp_id_stage_regfile_DataPath_mux_en_control_out, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N429_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3796 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_rd1_control_out, A2
                           => dp_id_stage_regfile_DataPath_mux_en_control_out, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N428_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3795 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n450, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n418, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2553, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2541
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3794 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2523, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2524, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2525
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2526, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2522);
   dp_id_stage_regfile_DataPath_Physical_RF_U3793 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2541, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2542, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2543
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2544, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2521);
   dp_id_stage_regfile_DataPath_Physical_RF_U3792 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2521, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2522, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N396_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3791 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n450, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n418, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3180, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3168
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3790 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3150, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3151, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3152
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3153, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3149);
   dp_id_stage_regfile_DataPath_Physical_RF_U3789 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3168, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3169, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3170
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3171, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3148);
   dp_id_stage_regfile_DataPath_Physical_RF_U3788 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3148, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3149, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N328_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3787 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n451, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n419, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2520, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2513
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3786 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2505, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2506, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2507
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2508, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2504);
   dp_id_stage_regfile_DataPath_Physical_RF_U3785 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2513, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2514, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2515
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2516, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2503);
   dp_id_stage_regfile_DataPath_Physical_RF_U3784 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2503, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2504, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N397_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3783 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n451, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n419, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3147, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3140
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3782 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3132, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3133, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3134
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3135, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3131);
   dp_id_stage_regfile_DataPath_Physical_RF_U3781 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3140, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3141, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3142
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3143, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3130);
   dp_id_stage_regfile_DataPath_Physical_RF_U3780 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3130, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3131, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N329_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3779 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n452, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n420, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2502, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2495
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3778 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2487, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2488, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2489
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2490, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2486);
   dp_id_stage_regfile_DataPath_Physical_RF_U3777 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2495, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2496, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2497
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2498, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2485);
   dp_id_stage_regfile_DataPath_Physical_RF_U3776 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2485, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2486, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N398_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3775 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n452, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n420, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3129, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3122
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3774 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3114, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3115, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3116
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3117, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3113);
   dp_id_stage_regfile_DataPath_Physical_RF_U3773 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3122, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3123, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3124
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3125, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3112);
   dp_id_stage_regfile_DataPath_Physical_RF_U3772 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3112, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3113, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N330_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3771 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n453, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n421, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2484, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2477
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3770 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2469, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2470, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2471
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2472, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2468);
   dp_id_stage_regfile_DataPath_Physical_RF_U3769 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2477, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2478, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2479
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2480, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2467);
   dp_id_stage_regfile_DataPath_Physical_RF_U3768 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2467, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2468, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N399_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3767 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n453, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n421, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3111, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3104
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3766 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3096, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3097, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3098
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3099, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3095);
   dp_id_stage_regfile_DataPath_Physical_RF_U3765 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3104, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3105, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3106
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3107, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3094);
   dp_id_stage_regfile_DataPath_Physical_RF_U3764 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3094, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3095, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N331_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3763 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n454, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n422, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2466, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2459
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3762 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2451, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2452, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2453
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2454, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2450);
   dp_id_stage_regfile_DataPath_Physical_RF_U3761 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2459, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2460, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2461
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2462, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2449);
   dp_id_stage_regfile_DataPath_Physical_RF_U3760 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2449, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2450, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N400_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3759 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n454, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n422, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3093, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3086
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3758 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3078, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3079, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3080
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3081, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3077);
   dp_id_stage_regfile_DataPath_Physical_RF_U3757 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3086, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3087, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3088
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3089, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3076);
   dp_id_stage_regfile_DataPath_Physical_RF_U3756 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3076, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3077, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N332_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3755 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n455, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n423, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2448, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2441
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3754 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2433, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2434, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2435
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2436, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2432);
   dp_id_stage_regfile_DataPath_Physical_RF_U3753 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2441, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2442, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2443
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2444, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2431);
   dp_id_stage_regfile_DataPath_Physical_RF_U3752 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2431, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2432, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N401_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3751 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n455, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n423, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3075, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3068
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3750 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3060, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3061, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3062
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3063, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3059);
   dp_id_stage_regfile_DataPath_Physical_RF_U3749 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3068, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3069, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3070
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3071, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3058);
   dp_id_stage_regfile_DataPath_Physical_RF_U3748 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3058, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3059, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N333_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3747 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n456, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n424, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2430, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2423
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3746 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2415, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2416, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2417
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2418, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2414);
   dp_id_stage_regfile_DataPath_Physical_RF_U3745 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2423, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2424, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2425
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2426, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2413);
   dp_id_stage_regfile_DataPath_Physical_RF_U3744 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2413, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2414, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N402_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3743 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n456, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n424, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3057, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3050
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3742 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3042, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3043, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3044
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3045, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3041);
   dp_id_stage_regfile_DataPath_Physical_RF_U3741 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3050, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3051, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3052
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3053, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3040);
   dp_id_stage_regfile_DataPath_Physical_RF_U3740 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3040, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3041, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N334_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3739 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n457, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n425, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2412, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2405
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3738 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2397, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2398, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2399
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2400, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2396);
   dp_id_stage_regfile_DataPath_Physical_RF_U3737 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2405, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2406, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2407
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2408, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2395);
   dp_id_stage_regfile_DataPath_Physical_RF_U3736 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2395, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2396, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N403_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3735 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n457, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n425, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3039, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3032
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3734 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3024, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3025, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3026
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3027, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3023);
   dp_id_stage_regfile_DataPath_Physical_RF_U3733 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3032, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3033, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3034
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3035, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3022);
   dp_id_stage_regfile_DataPath_Physical_RF_U3732 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3022, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3023, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N335_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3731 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n458, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n426, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2394, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2387
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3730 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2379, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2380, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2381
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2382, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2378);
   dp_id_stage_regfile_DataPath_Physical_RF_U3729 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2387, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2388, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2389
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2390, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2377);
   dp_id_stage_regfile_DataPath_Physical_RF_U3728 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2377, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2378, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N404_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3727 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n458, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n426, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3021, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3014
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3726 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3006, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3007, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3008
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3009, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3005);
   dp_id_stage_regfile_DataPath_Physical_RF_U3725 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3014, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3015, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n3016
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3017, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3004);
   dp_id_stage_regfile_DataPath_Physical_RF_U3724 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3004, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3005, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N336_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3723 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n459, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n427, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2376, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2369
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3722 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2361, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2362, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2363
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2364, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2360);
   dp_id_stage_regfile_DataPath_Physical_RF_U3721 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2369, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2370, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2371
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2372, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2359);
   dp_id_stage_regfile_DataPath_Physical_RF_U3720 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2359, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2360, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N405_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3719 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n459, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n427, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3003, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2996
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3718 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2988, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2989, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2990
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2991, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2987);
   dp_id_stage_regfile_DataPath_Physical_RF_U3717 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2996, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2997, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2998
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2999, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2986);
   dp_id_stage_regfile_DataPath_Physical_RF_U3716 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2986, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2987, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N337_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3715 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n460, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n428, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2358, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2351
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3714 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2343, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2344, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2345
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2346, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2342);
   dp_id_stage_regfile_DataPath_Physical_RF_U3713 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2351, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2352, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2353
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2354, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2341);
   dp_id_stage_regfile_DataPath_Physical_RF_U3712 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2341, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2342, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N406_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3711 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n460, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n428, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2985, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2978
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3710 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2970, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2971, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2972
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2973, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2969);
   dp_id_stage_regfile_DataPath_Physical_RF_U3709 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2978, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2979, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2980
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2981, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2968);
   dp_id_stage_regfile_DataPath_Physical_RF_U3708 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2968, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2969, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N338_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3707 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n461, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n429, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3760, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2340, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2333
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3706 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2325, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2326, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2327
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2328, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2324);
   dp_id_stage_regfile_DataPath_Physical_RF_U3705 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2333, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2334, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2335
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2336, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2323);
   dp_id_stage_regfile_DataPath_Physical_RF_U3704 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2323, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2324, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N407_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3703 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n461, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n429, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1212, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2967, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2960
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3702 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2952, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2953, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2954
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2955, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2951);
   dp_id_stage_regfile_DataPath_Physical_RF_U3701 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2960, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2961, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2962
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2963, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2950);
   dp_id_stage_regfile_DataPath_Physical_RF_U3700 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2950, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2951, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N339_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3699 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n462, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n430, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2322, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2315
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3698 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2307, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2308, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2309
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2310, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2306);
   dp_id_stage_regfile_DataPath_Physical_RF_U3697 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2315, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2316, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2317
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2318, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2305);
   dp_id_stage_regfile_DataPath_Physical_RF_U3696 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2305, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2306, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N408_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3695 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n462, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n430, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2949, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2942
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3694 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2934, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2935, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2936
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2937, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2933);
   dp_id_stage_regfile_DataPath_Physical_RF_U3693 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2942, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2943, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2944
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2945, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2932);
   dp_id_stage_regfile_DataPath_Physical_RF_U3692 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2932, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2933, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N340_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3691 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n463, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n431, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2304, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2297
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3690 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2289, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2290, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2291
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2292, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2288);
   dp_id_stage_regfile_DataPath_Physical_RF_U3689 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2297, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2298, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2299
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2300, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2287);
   dp_id_stage_regfile_DataPath_Physical_RF_U3688 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2287, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2288, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N409_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3687 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n463, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n431, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2931, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2924
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3686 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2916, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2917, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2918
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2919, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2915);
   dp_id_stage_regfile_DataPath_Physical_RF_U3685 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2924, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2925, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2926
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2927, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2914);
   dp_id_stage_regfile_DataPath_Physical_RF_U3684 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2914, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2915, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N341_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3683 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n464, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n432, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2286, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2279
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3682 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2271, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2272, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2273
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2274, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2270);
   dp_id_stage_regfile_DataPath_Physical_RF_U3681 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2279, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2280, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2281
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2282, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2269);
   dp_id_stage_regfile_DataPath_Physical_RF_U3680 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2270, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N410_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3679 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n464, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n432, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2913, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2906
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3678 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2898, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2899, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2900
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2901, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2897);
   dp_id_stage_regfile_DataPath_Physical_RF_U3677 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2906, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2907, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2908
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2909, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2896);
   dp_id_stage_regfile_DataPath_Physical_RF_U3676 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2896, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2897, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N342_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3675 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n465, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n433, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2268, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2261
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3674 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2254, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2255
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2256, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2252);
   dp_id_stage_regfile_DataPath_Physical_RF_U3673 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2262, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2263
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2264, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2251);
   dp_id_stage_regfile_DataPath_Physical_RF_U3672 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2252, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N411_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3671 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n465, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n433, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2895, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2888
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3670 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2880, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2881, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2882
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2883, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2879);
   dp_id_stage_regfile_DataPath_Physical_RF_U3669 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2888, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2889, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2890
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2891, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2878);
   dp_id_stage_regfile_DataPath_Physical_RF_U3668 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2878, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2879, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N343_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3667 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n466, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n434, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2250, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2243
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3666 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2235, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2236, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2237
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2238, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2234);
   dp_id_stage_regfile_DataPath_Physical_RF_U3665 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2244, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2245
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2246, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2233);
   dp_id_stage_regfile_DataPath_Physical_RF_U3664 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2233, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2234, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N412_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3663 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n466, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n434, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2877, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2870
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3662 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2862, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2863, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2864
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2865, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2861);
   dp_id_stage_regfile_DataPath_Physical_RF_U3661 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2870, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2871, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2872
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2873, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2860);
   dp_id_stage_regfile_DataPath_Physical_RF_U3660 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2860, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2861, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N344_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3659 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n467, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n435, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2232, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2225
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3658 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2217, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2218, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2219
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2220, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2216);
   dp_id_stage_regfile_DataPath_Physical_RF_U3657 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2225, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2226, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2227
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2228, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2215);
   dp_id_stage_regfile_DataPath_Physical_RF_U3656 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2215, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2216, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N413_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3655 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n467, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n435, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2859, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2852
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3654 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2844, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2845, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2846
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2847, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2843);
   dp_id_stage_regfile_DataPath_Physical_RF_U3653 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2852, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2853, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2854
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2855, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2842);
   dp_id_stage_regfile_DataPath_Physical_RF_U3652 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2842, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2843, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N345_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3651 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n468, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n436, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2214, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2207
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3650 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2199, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2200, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2201
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2202, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2198);
   dp_id_stage_regfile_DataPath_Physical_RF_U3649 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2207, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2208, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2209
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2210, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2197);
   dp_id_stage_regfile_DataPath_Physical_RF_U3648 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2197, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2198, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N414_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3647 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n468, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n436, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2841, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2834
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3646 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2826, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2827, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2828
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2829, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2825);
   dp_id_stage_regfile_DataPath_Physical_RF_U3645 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2834, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2835, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2836
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2837, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2824);
   dp_id_stage_regfile_DataPath_Physical_RF_U3644 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2824, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2825, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N346_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3643 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n469, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n437, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2196, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2189
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3642 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2181, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2182, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2183
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2184, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2180);
   dp_id_stage_regfile_DataPath_Physical_RF_U3641 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2189, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2190, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2191
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2192, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2179);
   dp_id_stage_regfile_DataPath_Physical_RF_U3640 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2179, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2180, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N415_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3639 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n469, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n437, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2823, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2816
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3638 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2808, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2809, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2810
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2811, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2807);
   dp_id_stage_regfile_DataPath_Physical_RF_U3637 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2816, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2817, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2818
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2819, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2806);
   dp_id_stage_regfile_DataPath_Physical_RF_U3636 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2806, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2807, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N347_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3635 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n470, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n438, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2178, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2171
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3634 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2163, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2164, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2165
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2166, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2162);
   dp_id_stage_regfile_DataPath_Physical_RF_U3633 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2171, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2172, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2173
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2174, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2161);
   dp_id_stage_regfile_DataPath_Physical_RF_U3632 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2161, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2162, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N416_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3631 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n470, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n438, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2805, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2798
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3630 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2790, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2791, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2792
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2793, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2789);
   dp_id_stage_regfile_DataPath_Physical_RF_U3629 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2798, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2799, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2800
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2801, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2788);
   dp_id_stage_regfile_DataPath_Physical_RF_U3628 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2788, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2789, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N348_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3627 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n471, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n439, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2153
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3626 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2145, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2146, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2147
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2148, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2144);
   dp_id_stage_regfile_DataPath_Physical_RF_U3625 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2153, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2154, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2155
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2156, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2143);
   dp_id_stage_regfile_DataPath_Physical_RF_U3624 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2143, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2144, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N417_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3623 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n471, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n439, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2787, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2780
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3622 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2772, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2773, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2774
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2775, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2771);
   dp_id_stage_regfile_DataPath_Physical_RF_U3621 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2780, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2781, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2782
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2783, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2770);
   dp_id_stage_regfile_DataPath_Physical_RF_U3620 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2770, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2771, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N349_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3619 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n472, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n440, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2142, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2135
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3618 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2127, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2128, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2129
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2130, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2126);
   dp_id_stage_regfile_DataPath_Physical_RF_U3617 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2135, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2136, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2137
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2138, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2125);
   dp_id_stage_regfile_DataPath_Physical_RF_U3616 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2125, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2126, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N418_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3615 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n472, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n440, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2769, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2762
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3614 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2754, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2755, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2756
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2757, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2753);
   dp_id_stage_regfile_DataPath_Physical_RF_U3613 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2762, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2763, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2764
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2765, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2752);
   dp_id_stage_regfile_DataPath_Physical_RF_U3612 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2752, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2753, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N350_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3611 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n473, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n441, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3761, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2124, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2117
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3610 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2109, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2110, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2111
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2112, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2108);
   dp_id_stage_regfile_DataPath_Physical_RF_U3609 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2117, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2118, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2119
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2120, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2107);
   dp_id_stage_regfile_DataPath_Physical_RF_U3608 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2107, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2108, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N419_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3607 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n473, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n441, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1213, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2751, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2744
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3606 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2736, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2737, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2738
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2739, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2735);
   dp_id_stage_regfile_DataPath_Physical_RF_U3605 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2744, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2745, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2746
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2747, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2734);
   dp_id_stage_regfile_DataPath_Physical_RF_U3604 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2734, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2735, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N351_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3603 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n474, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n442, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3762, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2106, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2099
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3602 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2091, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2092, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2093
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2094, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2090);
   dp_id_stage_regfile_DataPath_Physical_RF_U3601 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2099, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2100, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2101
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2102, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2089);
   dp_id_stage_regfile_DataPath_Physical_RF_U3600 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2089, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2090, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N420_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3599 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n474, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n442, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1214, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2733, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2726
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3598 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2718, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2719, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2720
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2721, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2717);
   dp_id_stage_regfile_DataPath_Physical_RF_U3597 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2726, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2727, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2728
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2729, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2716);
   dp_id_stage_regfile_DataPath_Physical_RF_U3596 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2716, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2717, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N352_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3595 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n475, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n443, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3762, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2088, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2081
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3594 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2073, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2074, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2075
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2076, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2072);
   dp_id_stage_regfile_DataPath_Physical_RF_U3593 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2081, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2082, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2083
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2084, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2071);
   dp_id_stage_regfile_DataPath_Physical_RF_U3592 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2071, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2072, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N421_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3591 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n475, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n443, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1214, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2715, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2708
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3590 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2700, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2701, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2702
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2703, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2699);
   dp_id_stage_regfile_DataPath_Physical_RF_U3589 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2708, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2709, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2710
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2711, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2698);
   dp_id_stage_regfile_DataPath_Physical_RF_U3588 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2698, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2699, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N353_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3587 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n476, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n444, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3762, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2070, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2063
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3586 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2055, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2056, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2057
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2058, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2054);
   dp_id_stage_regfile_DataPath_Physical_RF_U3585 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2063, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2064, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2065
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2066, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2053);
   dp_id_stage_regfile_DataPath_Physical_RF_U3584 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2053, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2054, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N422_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3583 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n476, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n444, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1214, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2697, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2690
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3582 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2682, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2683, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2684
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2685, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2681);
   dp_id_stage_regfile_DataPath_Physical_RF_U3581 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2690, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2691, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2692
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2693, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2680);
   dp_id_stage_regfile_DataPath_Physical_RF_U3580 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2680, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2681, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N354_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3579 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n477, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n445, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3762, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2052, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2045
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3578 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2037, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2038, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2039
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2040, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2036);
   dp_id_stage_regfile_DataPath_Physical_RF_U3577 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2045, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2046, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2047
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2048, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2035);
   dp_id_stage_regfile_DataPath_Physical_RF_U3576 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2035, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2036, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N423_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3575 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n477, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n445, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1214, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2679, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2672
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3574 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2664, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2665, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2666
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2667, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2663);
   dp_id_stage_regfile_DataPath_Physical_RF_U3573 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2672, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2673, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2674
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2675, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2662);
   dp_id_stage_regfile_DataPath_Physical_RF_U3572 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2662, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2663, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N355_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3571 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n478, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n446, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3762, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2034, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2027
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3570 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2019, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2020, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2021
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2022, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2018);
   dp_id_stage_regfile_DataPath_Physical_RF_U3569 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2027, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2028, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2029
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2030, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2017);
   dp_id_stage_regfile_DataPath_Physical_RF_U3568 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2017, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2018, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N424_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3567 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n478, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n446, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1214, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2661, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2654
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3566 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2646, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2647, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2648
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2649, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2645);
   dp_id_stage_regfile_DataPath_Physical_RF_U3565 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2654, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2655, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2656
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2657, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2644);
   dp_id_stage_regfile_DataPath_Physical_RF_U3564 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2644, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2645, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N356_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3563 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n479, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n447, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3762, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2016, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2009
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3562 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2001, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2002, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2003
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2004, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2000);
   dp_id_stage_regfile_DataPath_Physical_RF_U3561 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2009, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2010, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2011
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2012, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1999);
   dp_id_stage_regfile_DataPath_Physical_RF_U3560 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1999, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2000, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N425_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3559 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n479, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n447, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1214, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2643, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2636
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3558 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2628, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2629, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2630
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2631, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2627);
   dp_id_stage_regfile_DataPath_Physical_RF_U3557 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2636, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2637, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2638
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2639, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2626);
   dp_id_stage_regfile_DataPath_Physical_RF_U3556 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2626, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2627, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N357_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3555 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n480, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n448, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3762, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1998, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1991
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3554 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1983, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1984, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1985
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1986, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1982);
   dp_id_stage_regfile_DataPath_Physical_RF_U3553 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1991, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1992, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1993
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1994, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1981);
   dp_id_stage_regfile_DataPath_Physical_RF_U3552 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1981, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1982, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N426_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3551 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n480, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n448, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1214, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2625, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2618
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3550 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2610, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2611, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2612
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2613, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2609);
   dp_id_stage_regfile_DataPath_Physical_RF_U3549 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2618, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2619, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2620
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2621, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2608);
   dp_id_stage_regfile_DataPath_Physical_RF_U3548 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2608, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2609, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N358_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3547 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n481, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n449, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3762, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1977, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1955
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3546 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1929, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1930, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1931
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1932, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1928);
   dp_id_stage_regfile_DataPath_Physical_RF_U3545 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1955, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1956, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1957
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1958, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1927);
   dp_id_stage_regfile_DataPath_Physical_RF_U3544 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1927, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1928, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N427_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3543 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n481, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n449, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1214, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2604, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2582
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3542 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2556, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2557, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2558
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2559, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2555);
   dp_id_stage_regfile_DataPath_Physical_RF_U3541 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2582, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2583, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n2584
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2585, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2554);
   dp_id_stage_regfile_DataPath_Physical_RF_U3540 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2554, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2555, 
                           ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N359_port);
   dp_id_stage_regfile_DataPath_Physical_RF_U3539 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3810
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_31_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3807
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2540
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3538 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1026, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n994,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3814
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2540, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2523);
   dp_id_stage_regfile_DataPath_Physical_RF_U3537 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3702
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_31_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3699
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3167
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3536 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1026, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n994,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3706
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3167, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3150);
   dp_id_stage_regfile_DataPath_Physical_RF_U3535 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3810
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_30_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3807
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2512
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3534 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1027, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n995,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3814
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2512, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2505);
   dp_id_stage_regfile_DataPath_Physical_RF_U3533 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3702
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_30_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3699
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3139
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3532 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1027, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n995,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3706
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3139, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3132);
   dp_id_stage_regfile_DataPath_Physical_RF_U3531 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3810
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_29_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3807
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2494
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3530 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1028, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n996,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3814
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2494, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2487);
   dp_id_stage_regfile_DataPath_Physical_RF_U3529 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3702
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_29_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3699
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3121
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3528 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1028, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n996,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3706
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3121, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3114);
   dp_id_stage_regfile_DataPath_Physical_RF_U3527 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3810
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_28_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3807
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2476
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3526 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1029, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n997,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3814
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2476, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2469);
   dp_id_stage_regfile_DataPath_Physical_RF_U3525 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3702
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_28_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3699
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3103
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3524 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1029, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n997,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3706
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3103, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3096);
   dp_id_stage_regfile_DataPath_Physical_RF_U3523 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3810
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_27_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3807
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2458
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3522 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1030, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n998,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3814
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2458, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2451);
   dp_id_stage_regfile_DataPath_Physical_RF_U3521 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3702
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_27_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3699
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3085
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3520 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1030, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n998,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3706
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3085, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3078);
   dp_id_stage_regfile_DataPath_Physical_RF_U3519 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3810
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_26_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3807
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2440
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3518 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1031, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n999,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3814
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2440, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2433);
   dp_id_stage_regfile_DataPath_Physical_RF_U3517 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3702
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_26_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3699
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3067
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3516 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1031, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n999,
                           C2 => dp_id_stage_regfile_DataPath_Physical_RF_n3706
                           , A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3067, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3060);
   dp_id_stage_regfile_DataPath_Physical_RF_U3515 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3810
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_25_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3807
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2422
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3514 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1032, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1000
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3814, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2422, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2415);
   dp_id_stage_regfile_DataPath_Physical_RF_U3513 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3702
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_25_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3699
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3049
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3512 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1032, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1000
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3706, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3049, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3042);
   dp_id_stage_regfile_DataPath_Physical_RF_U3511 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3810
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_24_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3807
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2404
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3510 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1033, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1001
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3814, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2404, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2397);
   dp_id_stage_regfile_DataPath_Physical_RF_U3509 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3702
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_24_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3699
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3031
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3508 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1033, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1001
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3706, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3031, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3024);
   dp_id_stage_regfile_DataPath_Physical_RF_U3507 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_23_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2386
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3506 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1034, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1002
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3814, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2386, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2379);
   dp_id_stage_regfile_DataPath_Physical_RF_U3505 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_23_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3013
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3504 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1034, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1002
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3706, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3013, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3006);
   dp_id_stage_regfile_DataPath_Physical_RF_U3503 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_22_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2368
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3502 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1035, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1003
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3814, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2368, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2361);
   dp_id_stage_regfile_DataPath_Physical_RF_U3501 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_22_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2995
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3500 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1035, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1003
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3706, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2995, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2988);
   dp_id_stage_regfile_DataPath_Physical_RF_U3499 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_21_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2350
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3498 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1036, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1004
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3814, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2350, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2343);
   dp_id_stage_regfile_DataPath_Physical_RF_U3497 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_21_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2977
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3496 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1036, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1004
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3706, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2977, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2970);
   dp_id_stage_regfile_DataPath_Physical_RF_U3495 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_20_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2332
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3494 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1037, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3817, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1005
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3814, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2332, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2325);
   dp_id_stage_regfile_DataPath_Physical_RF_U3493 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_20_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2959
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3492 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1037, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3709, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1005
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3706, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2959, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2952);
   dp_id_stage_regfile_DataPath_Physical_RF_U3491 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_19_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2314
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3490 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1038, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1006
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2314, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2307);
   dp_id_stage_regfile_DataPath_Physical_RF_U3489 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_19_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2941
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3488 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1038, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1006
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2941, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2934);
   dp_id_stage_regfile_DataPath_Physical_RF_U3487 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_18_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2296
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3486 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1039, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1007
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2296, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2289);
   dp_id_stage_regfile_DataPath_Physical_RF_U3485 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_18_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2923
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3484 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1039, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1007
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2923, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2916);
   dp_id_stage_regfile_DataPath_Physical_RF_U3483 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_17_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2278
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3482 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1040, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1008
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2278, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2271);
   dp_id_stage_regfile_DataPath_Physical_RF_U3481 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_17_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2905
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3480 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1040, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1008
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2905, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2898);
   dp_id_stage_regfile_DataPath_Physical_RF_U3479 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_16_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2260
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3478 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1041, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1009
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2260, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2253);
   dp_id_stage_regfile_DataPath_Physical_RF_U3477 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_16_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2887
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3476 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1041, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1009
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2887, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2880);
   dp_id_stage_regfile_DataPath_Physical_RF_U3475 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_15_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2242
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3474 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1042, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1010
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2242, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2235);
   dp_id_stage_regfile_DataPath_Physical_RF_U3473 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_15_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2869
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3472 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1042, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1010
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2869, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2862);
   dp_id_stage_regfile_DataPath_Physical_RF_U3471 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_14_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2224
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3470 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1043, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1011
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2224, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2217);
   dp_id_stage_regfile_DataPath_Physical_RF_U3469 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_14_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2851
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3468 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1043, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1011
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2851, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2844);
   dp_id_stage_regfile_DataPath_Physical_RF_U3467 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_13_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2206
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3466 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1044, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1012
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2206, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2199);
   dp_id_stage_regfile_DataPath_Physical_RF_U3465 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_13_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2833
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3464 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1044, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1012
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2833, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2826);
   dp_id_stage_regfile_DataPath_Physical_RF_U3463 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3809
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_12_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3806
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2188
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3462 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1045, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1013
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2188, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2181);
   dp_id_stage_regfile_DataPath_Physical_RF_U3461 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3701
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_12_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3698
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2815
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3460 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1045, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1013
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2815, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2808);
   dp_id_stage_regfile_DataPath_Physical_RF_U3459 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_11_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2170
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3458 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1046, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1014
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2170, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2163);
   dp_id_stage_regfile_DataPath_Physical_RF_U3457 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_11_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2797
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3456 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1046, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1014
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2797, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2790);
   dp_id_stage_regfile_DataPath_Physical_RF_U3455 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_10_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2152
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3454 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1047, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1015
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2152, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2145);
   dp_id_stage_regfile_DataPath_Physical_RF_U3453 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_10_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2779
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3452 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1047, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1015
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2779, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2772);
   dp_id_stage_regfile_DataPath_Physical_RF_U3451 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_9_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2134
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3450 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1048, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1016
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2134, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2127);
   dp_id_stage_regfile_DataPath_Physical_RF_U3449 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_9_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2761
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3448 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1048, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1016
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2761, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2754);
   dp_id_stage_regfile_DataPath_Physical_RF_U3447 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_8_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2116
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3446 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1049, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3818, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1017
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2116, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2109);
   dp_id_stage_regfile_DataPath_Physical_RF_U3445 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_8_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2743
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3444 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1049, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3710, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1017
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2743, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2736);
   dp_id_stage_regfile_DataPath_Physical_RF_U3443 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_7_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2098
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3442 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1050, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1018
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2098, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2091);
   dp_id_stage_regfile_DataPath_Physical_RF_U3441 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_7_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2725
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3440 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1050, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1018
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2725, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2718);
   dp_id_stage_regfile_DataPath_Physical_RF_U3439 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_6_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2080
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3438 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1051, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1019
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2080, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2073);
   dp_id_stage_regfile_DataPath_Physical_RF_U3437 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_6_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2707
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3436 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1051, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1019
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2707, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2700);
   dp_id_stage_regfile_DataPath_Physical_RF_U3435 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_5_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2062
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3434 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1052, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1020
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2062, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2055);
   dp_id_stage_regfile_DataPath_Physical_RF_U3433 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_5_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2689
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3432 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1052, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1020
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2689, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2682);
   dp_id_stage_regfile_DataPath_Physical_RF_U3431 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_4_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2044
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3430 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1053, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1021
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2044, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2037);
   dp_id_stage_regfile_DataPath_Physical_RF_U3429 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_4_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2671
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3428 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1053, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1021
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2671, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2664);
   dp_id_stage_regfile_DataPath_Physical_RF_U3427 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_3_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2026
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3426 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1054, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1022
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2026, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2019);
   dp_id_stage_regfile_DataPath_Physical_RF_U3425 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_3_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2653
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3424 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1054, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1022
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2653, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2646);
   dp_id_stage_regfile_DataPath_Physical_RF_U3423 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_2_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2008
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3422 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1055, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1023
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2008, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2001);
   dp_id_stage_regfile_DataPath_Physical_RF_U3421 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_2_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2635
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3420 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1055, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1023
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2635, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2628);
   dp_id_stage_regfile_DataPath_Physical_RF_U3419 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_1_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1990
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3418 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1056, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1024
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1990, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1983);
   dp_id_stage_regfile_DataPath_Physical_RF_U3417 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_1_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2617
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3416 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1056, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1024
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2617, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2610);
   dp_id_stage_regfile_DataPath_Physical_RF_U3415 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3808
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_0_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3805
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1951
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3414 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1057, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3819, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1025
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1951, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1929);
   dp_id_stage_regfile_DataPath_Physical_RF_U3413 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3700
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_0_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3697
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2578
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3412 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1057, B2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3711, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1025
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708, A =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n2578, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2556);
   dp_id_stage_regfile_DataPath_Physical_RF_U3411 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3768
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2550
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3410 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n322, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n290, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2550, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2542
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3409 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3822
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2537
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3408 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n962, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n930, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2537, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2524
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3407 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1220
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3177
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3406 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n322, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n290, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3177, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3169
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3405 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3714
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3164
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3404 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n962, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n930, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3164, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3151
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3403 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3768
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2519
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3402 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n323, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n291, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2519, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2514
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3401 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3822
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2511
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3400 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n963, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n931, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2511, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2506
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3399 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1220
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3146
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3398 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n323, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n291, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3146, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3141
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3397 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3714
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3138
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3396 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n963, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n931, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3138, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3133
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3395 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3768
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2501
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3394 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n324, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n292, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2501, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2496
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3393 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3822
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2493
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3392 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n964, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n932, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2493, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2488
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3391 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1220
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3128
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3390 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n324, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n292, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3128, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3123
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3389 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3714
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3120
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3388 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n964, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n932, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3120, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3115
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3387 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3768
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2483
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3386 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n325, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n293, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2483, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2478
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3385 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3822
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2475
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3384 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n965, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n933, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2475, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2470
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3383 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1220
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3110
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3382 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n325, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n293, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3110, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3105
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3381 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3714
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3102
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3380 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n965, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n933, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3102, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3097
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3379 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3768
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2465
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3378 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n326, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n294, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2465, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2460
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3377 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3822
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2457
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3376 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n966, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n934, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2457, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2452
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3375 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1220
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3092
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3374 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n326, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n294, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3092, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3087
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3373 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3714
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3084
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3372 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n966, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n934, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3084, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3079
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3371 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3768
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2447
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3370 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n327, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n295, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2447, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2442
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3369 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3822
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2439
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3368 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n967, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n935, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2439, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2434
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3367 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1220
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3074
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3366 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n327, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n295, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3074, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3069
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3365 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3714
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3066
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3364 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n967, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n935, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3066, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3061
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3363 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3768
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2429
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3362 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n328, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n296, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2429, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2424
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3361 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3822
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2421
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3360 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n968, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n936, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2421, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2416
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3359 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1220
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3056
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3358 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n328, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n296, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3056, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3051
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3357 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3714
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3048
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3356 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n968, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n936, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3048, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3043
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3355 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3768
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2411
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3354 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n329, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n297, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2411, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2406
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3353 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3822
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2403
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3352 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n969, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n937, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2403, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2398
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3351 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1220
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3038
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3350 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n329, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n297, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3038, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3033
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3349 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3714
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3030
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3348 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n969, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n937, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3030, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3025
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3347 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2393
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3346 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n330, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n298, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2393, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2388
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3345 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2385
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3344 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n970, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n938, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2385, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2380
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3343 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3020
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3342 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n330, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n298, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3020, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3015
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3341 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3012
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3340 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n970, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n938, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3012, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3007
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3339 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2375
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3338 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n331, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n299, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2375, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2370
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3337 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2367
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3336 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n971, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n939, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2367, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2362
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3335 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3002
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3334 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n331, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n299, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3002, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2997
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3333 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2994
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3332 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n971, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n939, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2994, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2989
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3331 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2357
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3330 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n332, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n300, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2357, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2352
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3329 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2349
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3328 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n972, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n940, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2349, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2344
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3327 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2984
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3326 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n332, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n300, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2984, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2979
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3325 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2976
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3324 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n972, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n940, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2976, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2971
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3323 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2339
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3322 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n333, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n301, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3772, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2339, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2334
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3321 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2331
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3320 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n973, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n941, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3826, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2331, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2326
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3319 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2966
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3318 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n333, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n301, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1224, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2966, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2961
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3317 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2958
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3316 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n973, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n941, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3718, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2958, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2953
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3315 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2321
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3314 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n334, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n302, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2321, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2316
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3313 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2313
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3312 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n974, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n942, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2313, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2308
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3311 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2948
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3310 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n334, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n302, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2948, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2943
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3309 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2940
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3308 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n974, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n942, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2940, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2935
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3307 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2303
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3306 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n335, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n303, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2303, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2298
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3305 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2295
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3304 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n975, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n943, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2295, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2290
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3303 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2930
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3302 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n335, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n303, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2930, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2925
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3301 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2922
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3300 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n975, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n943, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2922, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2917
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3299 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2285
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3298 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n336, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n304, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2285, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2280
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3297 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2277
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3296 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n976, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n944, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2277, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2272
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3295 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2912
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3294 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n336, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n304, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2912, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2907
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3293 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2904
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3292 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n976, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n944, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2904, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2899
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3291 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2267
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3290 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n337, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n305, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2267, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2262
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3289 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2259
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3288 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n977, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n945, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2259, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2254
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3287 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2894
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3286 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n337, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n305, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2894, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2889
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3285 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2886
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3284 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n977, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n945, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2886, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2881
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3283 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2249
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3282 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n338, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n306, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2249, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2244
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3281 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2241
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3280 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n978, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n946, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2241, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2236
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3279 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2876
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3278 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n338, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n306, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2876, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2871
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3277 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2868
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3276 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n978, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n946, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2868, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2863
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3275 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2231
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3274 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n339, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n307, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2231, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2226
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3273 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2223
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3272 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n979, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n947, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2223, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2218
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3271 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2858
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3270 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n339, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n307, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2858, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2853
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3269 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2850
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3268 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n979, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n947, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2850, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2845
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3267 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2213
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3266 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n340, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n308, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2213, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2208
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3265 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2205
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3264 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n980, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n948, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2205, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2200
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3263 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2840
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3262 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n340, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n308, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2840, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2835
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3261 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2832
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3260 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n980, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n948, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2832, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2827
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3259 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3767
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2195
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3258 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n341, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n309, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2195, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2190
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3257 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3821
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2187
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3256 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n981, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n949, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2187, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2182
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3255 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1219
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2822
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3254 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n341, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n309, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2822, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2817
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3253 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3713
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2814
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3252 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n981, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n949, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2814, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2809
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3251 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2177
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3250 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n342, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n310, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2177, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2172
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3249 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2169
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3248 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n982, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n950, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2169, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2164
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3247 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2804
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3246 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n342, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n310, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2804, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2799
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3245 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2796
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3244 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n982, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n950, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2796, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2791
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3243 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2159
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3242 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n343, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n311, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2154
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3241 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2151
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3240 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n983, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n951, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2151, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2146
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3239 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2786
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3238 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n343, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n311, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2786, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2781
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3237 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2778
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3236 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n983, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n951, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2778, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2773
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3235 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2141
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3234 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n344, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n312, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2141, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2136
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3233 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2133
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3232 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n984, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n952, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2133, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2128
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3231 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2768
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3230 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n344, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n312, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2768, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2763
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3229 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2760
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3228 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n984, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n952, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2760, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2755
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3227 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2123
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3226 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n345, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n313, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3773, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2123, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2118
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3225 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2115
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3224 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n985, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n953, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3827, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2115, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2110
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3223 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2750
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3222 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n345, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n313, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1225, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2750, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2745
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3221 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2742
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3220 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n985, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n953, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3719, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2742, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2737
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3219 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2105
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3218 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n346, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n314, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3774, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2105, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2100
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3217 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2097
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3216 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n986, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n954, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3828, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2097, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2092
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3215 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2732
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3214 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n346, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n314, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1226, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2732, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2727
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3213 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2724
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3212 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n986, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n954, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3720, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2724, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2719
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3211 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2087
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3210 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n347, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n315, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3774, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2087, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2082
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3209 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2079
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3208 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n987, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n955, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3828, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2079, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2074
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3207 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2714
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3206 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n347, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n315, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1226, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2714, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2709
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3205 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2706
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3204 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n987, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n955, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3720, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2706, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2701
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3203 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2069
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3202 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n348, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n316, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3774, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2069, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2064
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3201 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2061
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3200 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n988, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n956, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3828, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2061, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2056
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3199 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2696
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3198 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n348, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n316, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1226, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2696, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2691
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3197 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2688
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3196 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n988, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n956, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3720, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2688, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2683
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3195 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2051
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3194 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n349, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n317, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3774, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2051, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2046
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3193 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2043
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3192 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n989, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n957, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3828, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2043, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2038
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3191 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2678
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3190 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n349, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n317, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1226, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2678, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2673
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3189 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2670
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3188 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n989, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n957, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3720, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2670, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2665
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3187 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2033
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3186 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n350, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n318, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3774, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2033, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2028
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3185 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2025
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3184 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n990, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n958, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3828, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2025, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2020
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3183 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2660
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3182 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n350, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n318, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1226, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2660, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2655
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3181 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2652
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3180 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n990, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n958, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3720, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2652, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2647
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3179 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2015
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3178 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n351, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n319, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3774, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2015, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2010
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3177 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2007
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3176 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n991, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n959, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3828, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2007, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2002
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3175 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2642
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3174 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n351, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n319, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1226, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2642, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2637
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3173 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2634
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3172 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n991, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n959, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3720, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2634, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2629
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3171 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1997
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3170 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n352, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n320, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3774, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1997, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1992
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3169 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1989
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3168 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n992, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n960, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3828, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1989, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1984
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3167 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2624
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3166 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n352, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n320, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1226, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2624, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2619
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3165 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2616
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3164 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n992, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n960, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3720, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2616, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2611
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3163 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3766
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1972
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3162 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n353, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n321, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3774, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1972, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1956
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3161 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3820
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1946
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3160 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n993, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n961, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3828, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1946, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1930
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3159 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1218
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2599
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3158 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n353, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n321, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1226, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2599, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2583
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3157 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3712
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2573
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3156 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n993, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n961, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3720, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2573, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2557
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3155 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3783
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_31_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3780
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2547
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3154 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n162, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n130, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2547, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2543
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3153 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3837
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_31_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3834
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2534
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3152 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n738, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n706, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2534, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2525
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3151 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1235
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_31_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1232
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3174
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3150 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n162, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n130, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3174, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3170
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3149 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3729
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_31_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3726
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3161
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3148 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n738, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n706, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3161, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3152
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3147 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3783
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_30_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3780
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2518
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3146 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n163, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n131, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2518, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2515
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3145 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3837
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_30_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3834
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2510
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3144 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n739, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n707, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2510, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2507
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3143 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1235
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_30_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1232
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3145
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3142 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n163, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n131, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3145, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3142
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3141 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3729
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_30_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3726
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3137
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3140 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n739, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n707, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3137, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3134
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3139 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3783
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_29_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3780
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2500
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3138 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n164, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n132, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2500, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2497
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3137 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3837
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_29_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3834
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2492
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3136 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n740, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n708, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2492, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2489
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3135 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1235
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_29_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1232
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3127
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3134 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n164, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n132, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3127, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3124
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3133 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3729
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_29_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3726
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3119
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3132 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n740, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n708, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3119, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3116
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3131 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3783
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_28_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3780
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2482
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3130 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n165, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n133, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2482, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2479
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3129 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3837
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_28_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3834
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2474
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3128 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n741, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n709, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2474, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2471
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3127 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1235
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_28_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1232
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3109
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3126 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n165, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n133, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3109, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3106
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3125 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3729
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_28_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3726
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3101
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3124 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n741, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n709, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3101, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3098
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3123 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3783
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_27_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3780
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2464
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3122 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n166, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n134, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2464, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2461
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3121 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3837
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_27_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3834
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2456
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3120 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n742, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n710, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2456, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2453
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3119 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1235
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_27_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1232
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3091
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3118 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n166, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n134, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3091, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3088
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3117 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3729
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_27_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3726
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3083
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3116 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n742, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n710, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3083, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3080
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3115 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3783
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_26_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3780
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2446
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3114 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n167, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n135, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2446, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2443
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3113 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3837
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_26_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3834
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2438
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3112 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n743, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n711, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2438, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2435
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3111 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1235
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_26_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1232
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3073
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3110 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n167, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n135, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3073, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3070
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3109 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3729
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_26_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3726
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3065
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3108 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n743, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n711, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3065, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3062
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3107 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3783
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_25_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3780
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2428
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3106 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n168, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n136, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2428, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2425
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3105 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3837
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_25_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3834
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2420
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3104 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n744, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n712, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2420, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2417
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3103 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1235
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_25_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1232
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3055
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3102 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n168, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n136, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3055, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3052
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3101 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3729
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_25_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3726
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3047
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3100 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n744, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n712, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3047, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3044
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3099 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3783
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_24_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3780
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2410
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3098 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n169, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n137, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2410, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2407
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3097 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3837
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_24_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3834
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2402
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3096 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n745, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n713, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2402, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2399
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3095 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1235
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_24_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1232
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3037
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3094 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n169, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n137, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3037, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3034
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3093 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3729
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_24_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3726
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3029
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3092 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n745, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n713, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3029, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3026
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3091 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_23_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2392
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3090 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n170, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n138, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2392, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2389
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3089 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_23_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2384
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3088 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n746, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n714, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2384, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2381
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3087 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_23_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3019
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3086 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n170, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n138, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3019, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3016
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3085 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_23_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3011
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3084 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n746, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n714, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3011, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3008
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3083 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_22_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2374
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3082 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n171, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n139, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2374, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2371
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3081 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_22_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2366
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3080 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n747, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n715, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2366, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2363
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3079 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_22_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3001
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3078 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n171, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n139, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3001, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2998
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3077 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_22_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2993
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3076 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n747, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n715, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2993, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2990
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3075 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_21_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2356
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3074 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n172, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n140, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2356, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2353
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3073 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_21_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2348
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3072 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n748, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n716, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2348, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2345
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3071 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_21_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2983
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3070 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n172, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n140, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2983, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2980
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3069 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_21_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2975
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3068 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n748, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n716, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2975, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2972
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3067 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_20_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2338
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3066 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n173, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n141, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3787, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2338, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2335
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3065 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_20_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2330
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3064 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n749, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n717, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3841, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2330, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2327
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3063 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_20_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2965
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3062 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n173, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n141, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1346, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2965, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2962
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3061 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_20_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2957
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3060 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n749, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n717, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3733, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2957, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2954
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3059 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_19_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2320
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3058 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n174, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n142, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2320, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2317
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3057 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_19_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2312
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3056 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n750, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n718, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2312, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2309
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3055 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_19_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2947
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3054 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n174, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n142, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2947, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2944
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3053 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_19_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2939
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3052 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n750, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n718, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2939, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2936
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3051 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_18_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2302
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3050 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n175, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n143, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2302, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2299
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3049 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_18_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2294
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3048 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n751, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n719, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2294, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2291
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3047 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_18_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2929
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3046 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n175, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n143, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2929, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2926
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3045 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_18_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2921
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3044 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n751, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n719, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2921, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2918
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3043 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_17_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2284
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3042 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n176, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n144, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2284, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2281
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3041 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_17_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2276
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3040 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n752, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n720, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2276, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2273
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3039 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_17_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2911
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3038 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n176, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n144, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2911, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2908
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3037 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_17_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2903
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3036 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n752, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n720, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2903, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2900
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3035 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_16_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2266
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3034 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n177, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n145, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2266, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2263
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3033 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_16_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2258
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3032 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n753, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n721, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2258, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2255
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3031 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_16_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2893
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3030 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n177, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n145, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2893, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2890
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3029 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_16_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2885
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3028 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n753, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n721, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2885, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2882
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3027 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_15_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2248
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3026 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n178, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n146, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2248, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2245
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3025 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_15_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2240
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3024 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n754, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n722, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2240, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2237
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3023 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_15_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2875
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3022 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n178, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n146, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2875, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2872
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3021 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_15_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2867
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3020 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n754, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n722, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2867, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2864
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3019 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_14_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2230
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3018 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n179, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n147, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2230, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2227
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3017 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_14_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2222
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3016 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n755, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n723, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2222, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2219
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3015 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_14_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2857
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3014 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n179, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n147, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2857, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2854
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3013 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_14_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2849
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3012 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n755, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n723, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2849, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2846
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3011 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_13_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2212
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3010 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n180, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n148, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2212, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2209
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3009 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_13_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2204
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3008 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n756, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n724, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2204, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2201
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3007 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_13_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2839
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3006 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n180, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n148, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2839, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2836
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3005 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_13_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2831
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3004 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n756, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n724, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2831, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2828
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3003 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3782
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_12_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3779
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2194
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3002 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n181, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n149, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2194, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2191
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3001 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3836
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_12_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3833
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2186
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U3000 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n757, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n725, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2186, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2183
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2999 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1234
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_12_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1231
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2821
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2998 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n181, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n149, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2821, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2818
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2997 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3728
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_12_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3725
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2813
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2996 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n757, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n725, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2813, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2810
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2995 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_11_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2176
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2994 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n182, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n150, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2176, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2173
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2993 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_11_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2168
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2992 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n758, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n726, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2168, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2165
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2991 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_11_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2803
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2990 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n182, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n150, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2803, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2800
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2989 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_11_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2795
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2988 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n758, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n726, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2795, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2792
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2987 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_10_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2158
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2986 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n183, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n151, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2158, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2155
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2985 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_10_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2150
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2984 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n759, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n727, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2150, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2147
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2983 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_10_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2785
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2982 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n183, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n151, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2785, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2782
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2981 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_10_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2777
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2980 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n759, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n727, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2777, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2774
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2979 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_9_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2140
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2978 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n184, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n152, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2140, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2137
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2977 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_9_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2132
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2976 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n760, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n728, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2132, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2129
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2975 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_9_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2767
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2974 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n184, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n152, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2767, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2764
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2973 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_9_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2759
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2972 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n760, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n728, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2759, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2756
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2971 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_8_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2122
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2970 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n185, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n153, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3788, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2122, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2119
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2969 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_8_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2114
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2968 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n761, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n729, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3842, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2114, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2111
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2967 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_8_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2749
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2966 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n185, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n153, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1348, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2749, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2746
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2965 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_8_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2741
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2964 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n761, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n729, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3734, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2741, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2738
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2963 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_7_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2104
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2962 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n186, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n154, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3789, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2104, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2101
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2961 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_7_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2096
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2960 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n762, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n730, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3843, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2096, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2093
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2959 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_7_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2731
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2958 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n186, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n154, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1516, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2731, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2728
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2957 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_7_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2723
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2956 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n762, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n730, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3735, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2723, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2720
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2955 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_6_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2086
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2954 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n187, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n155, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3789, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2086, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2083
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2953 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_6_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2078
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2952 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n763, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n731, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3843, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2078, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2075
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2951 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_6_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2713
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2950 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n187, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n155, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1516, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2713, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2710
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2949 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_6_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2705
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2948 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n763, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n731, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3735, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2705, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2702
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2947 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_5_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2068
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2946 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n188, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n156, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3789, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2068, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2065
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2945 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_5_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2060
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2944 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n764, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n732, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3843, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2060, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2057
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2943 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_5_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2695
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2942 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n188, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n156, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1516, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2695, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2692
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2941 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_5_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2687
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2940 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n764, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n732, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3735, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2687, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2684
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2939 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_4_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2050
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2938 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n189, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n157, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3789, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2050, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2047
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2937 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_4_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2042
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2936 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n765, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n733, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3843, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2042, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2039
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2935 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_4_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2677
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2934 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n189, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n157, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1516, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2677, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2674
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2933 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_4_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2669
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2932 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n765, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n733, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3735, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2669, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2666
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2931 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_3_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2032
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2930 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n190, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n158, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3789, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2032, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2029
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2929 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_3_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2024
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2928 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n766, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n734, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3843, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2024, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2021
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2927 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_3_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2659
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2926 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n190, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n158, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1516, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2659, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2656
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2925 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_3_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2651
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2924 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n766, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n734, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3735, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2651, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2648
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2923 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_2_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2014
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2922 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n191, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n159, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3789, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2014, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2011
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2921 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_2_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2006
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2920 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n767, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n735, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3843, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2006, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2003
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2919 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_2_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2641
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2918 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n191, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n159, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1516, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2641, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2638
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2917 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_2_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2633
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2916 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n767, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n735, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3735, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2633, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2630
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2915 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_1_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1996
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2914 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n192, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n160, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3789, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1996, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1993
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2913 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_1_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1988
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2912 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n768, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n736, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3843, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1988, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1985
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2911 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_1_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2623
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2910 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n192, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n160, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1516, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2623, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2620
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2909 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_1_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2615
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2908 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n768, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n736, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3735, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2615, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2612
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2907 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3781
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_0_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3778
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1966
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2906 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n193, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n161, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3789, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1966, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1957
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2905 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3835
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_0_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3832
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1940
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2904 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n769, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n737, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3843, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1940, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1931
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2903 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1233
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_0_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1230
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2593
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2902 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n193, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n161, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1516, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2593, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2584
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2901 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3727
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_0_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3724
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2567
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2900 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n769, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n737, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3735, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2567, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2558
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2899 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3795
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2545
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2898 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n34, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2545, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2544
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2897 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3849
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2527
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2896 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n610, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n578, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2527, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2526
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2895 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3172
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2894 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n34, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3172, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3171
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2893 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3741
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3154
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2892 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n610, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n578, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3154, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3153
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2891 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3795
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2517
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2890 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n35, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2517, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2516
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2889 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3849
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2509
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2888 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n611, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n579, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2509, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2508
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2887 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3144
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2886 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n35, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3144, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3143
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2885 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3741
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3136
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2884 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n611, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n579, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3136, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3135
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2883 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3795
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2499
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2882 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n36, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2499, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2498
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2881 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3849
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2491
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2880 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n612, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n580, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2491, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2490
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2879 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3126
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2878 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n36, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3126, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3125
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2877 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3741
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3118
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2876 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n612, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n580, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3118, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3117
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2875 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3795
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2481
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2874 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n37, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n5, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2481, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2480
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2873 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3849
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2473
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2872 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n613, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n581, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2473, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2472
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2871 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3108
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2870 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n37, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n5, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3108, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3107
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2869 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3741
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3100
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2868 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n613, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n581, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3100, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3099
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2867 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3795
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2463
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2866 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n38, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n6, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2463, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2462
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2865 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3849
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2455
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2864 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n614, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n582, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2455, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2454
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2863 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3090
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2862 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n38, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n6, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3090, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3089
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2861 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3741
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3082
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2860 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n614, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n582, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3082, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3081
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2859 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3795
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2445
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2858 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n39, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n7, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2445, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2444
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2857 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3849
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2437
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2856 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n615, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n583, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2437, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2436
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2855 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3072
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2854 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n39, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n7, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3072, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3071
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2853 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3741
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3064
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2852 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n615, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n583, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3064, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3063
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2851 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3795
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2427
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2850 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n40, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n8, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2427, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2426
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2849 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3849
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2419
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2848 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n616, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n584, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2419, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2418
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2847 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3054
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2846 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n40, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n8, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3054, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3053
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2845 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3741
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3046
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2844 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n616, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n584, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3046, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3045
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2843 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3795
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2409
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2842 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n41, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n9, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2409, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2408
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2841 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3849
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2401
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2840 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n617, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n585, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2401, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2400
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2839 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3036
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2838 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n41, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n9, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3036, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3035
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2837 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3741
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3028
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2836 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n617, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n585, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3028, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3027
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2835 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2391
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2834 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n42, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n10, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2391, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2390
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2833 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2383
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2832 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n618, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n586, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2383, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2382
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2831 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3018
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2830 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n42, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n10, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3018, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3017
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2829 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3010
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2828 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n618, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n586, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3010, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3009
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2827 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2373
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2826 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n43, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n11, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2373, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2372
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2825 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2365
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2824 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n619, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n587, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2365, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2364
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2823 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3000
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2822 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n43, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n11, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3000, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2999
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2821 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2992
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2820 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n619, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n587, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2992, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2991
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2819 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2355
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2818 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n44, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n12, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2355, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2354
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2817 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2347
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2816 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n620, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n588, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2347, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2346
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2815 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2982
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2814 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n44, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n12, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2982, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2981
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2813 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2974
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2812 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n620, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n588, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2974, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2973
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2811 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2337
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2810 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n45, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n13, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3799, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2337, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2336
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2809 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2329
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2808 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n621, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n589, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3853, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2329, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2328
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2807 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2964
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2806 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n45, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n13, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1925, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2964, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2963
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2805 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2956
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2804 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n621, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n589, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3745, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2956, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2955
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2803 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2319
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2802 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n46, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n14, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2319, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2318
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2801 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2311
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2800 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n622, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n590, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2311, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2310
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2799 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2946
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2798 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n46, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n14, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2946, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2945
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2797 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2938
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2796 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n622, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n590, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2938, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2937
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2795 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2301
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2794 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n47, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n15, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2301, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2300
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2793 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2293
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2792 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n623, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n591, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2293, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2292
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2791 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2928
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2790 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n47, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n15, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2928, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2927
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2789 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2920
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2788 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n623, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n591, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2920, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2919
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2787 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2283
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2786 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n48, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n16, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2283, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2282
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2785 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2275
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2784 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n624, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n592, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2275, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2274
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2783 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2910
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2782 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n48, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n16, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2910, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2909
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2781 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2902
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2780 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n624, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n592, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2902, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2901
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2779 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2265
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2778 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n49, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n17, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2265, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2264
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2777 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2257
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2776 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n625, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n593, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2257, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2256
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2775 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2892
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2774 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n49, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n17, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2892, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2891
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2773 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2884
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2772 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n625, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n593, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2884, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2883
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2771 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2247
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2770 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n50, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n18, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2247, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2246
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2769 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2239
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2768 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n626, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n594, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2239, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2238
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2767 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2874
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2766 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n50, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n18, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2874, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2873
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2765 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2866
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2764 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n626, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n594, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2866, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2865
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2763 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2229
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2762 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n51, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n19, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2229, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2228
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2761 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2221
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2760 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n627, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n595, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2221, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2220
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2759 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2856
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2758 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n51, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n19, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2856, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2855
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2757 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2848
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2756 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n627, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n595, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2848, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2847
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2755 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2211
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2754 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n52, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n20, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2211, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2210
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2753 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2203
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2752 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n628, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n596, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2203, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2202
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2751 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2838
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2750 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n52, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n20, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2838, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2837
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2749 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2830
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2748 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n628, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n596, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2830, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2829
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2747 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3794
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2193
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2746 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n53, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n21, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2193, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2192
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2745 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3848
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2185
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2744 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n629, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n597, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2185, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2184
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2743 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1688
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2820
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2742 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n53, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n21, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2820, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2819
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2741 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3740
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2812
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2740 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n629, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n597, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2812, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2811
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2739 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2175
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2738 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n54, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n22, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2175, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2174
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2737 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2167
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2736 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n630, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n598, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2167, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2166
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2735 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2802
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2734 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n54, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n22, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2802, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2801
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2733 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2794
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2732 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n630, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n598, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2794, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2793
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2731 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2157
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2730 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n55, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n23, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2156
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2729 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2149
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2728 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n631, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n599, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2149, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2148
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2727 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2784
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2726 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n55, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n23, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2784, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2783
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2725 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2776
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2724 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n631, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n599, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2776, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2775
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2723 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2139
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2722 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n56, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n24, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2139, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2138
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2721 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2131
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2720 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n632, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n600, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2131, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2130
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2719 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2766
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2718 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n56, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n24, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2766, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2765
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2717 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2758
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2716 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n632, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n600, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2758, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2757
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2715 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2121
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2714 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n57, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n25, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3800, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2121, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2120
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2713 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2113
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2712 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n633, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n601, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3854, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2113, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2112
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2711 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2748
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2710 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n57, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n25, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1926, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2748, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2747
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2709 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2740
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2708 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n633, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n601, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3746, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2740, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2739
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2707 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2103
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2706 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n58, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n26, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3801, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2103, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2102
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2705 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2095
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2704 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n634, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n602, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3855, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2095, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2094
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2703 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2730
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2702 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n58, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n26, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3693, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2730, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2729
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2701 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2722
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2700 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n634, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n602, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3747, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2722, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2721
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2699 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2085
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2698 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n59, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n27, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3801, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2085, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2084
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2697 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2077
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2696 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n635, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n603, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3855, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2077, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2076
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2695 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2712
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2694 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n59, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n27, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3693, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2712, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2711
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2693 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2704
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2692 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n635, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n603, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3747, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2704, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2703
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2691 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2067
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2690 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n60, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n28, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3801, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2067, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2066
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2689 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2059
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2688 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n636, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n604, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3855, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2059, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2058
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2687 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2694
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2686 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n60, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n28, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3693, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2694, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2693
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2685 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2686
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2684 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n636, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n604, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3747, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2686, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2685
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2683 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2049
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2682 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n61, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n29, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3801, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2049, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2048
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2681 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2041
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2680 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n637, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n605, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3855, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2041, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2040
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2679 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2676
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2678 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n61, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n29, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3693, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2676, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2675
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2677 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2668
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2676 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n637, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n605, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3747, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2668, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2667
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2675 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2031
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2674 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n62, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n30, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3801, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2031, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2030
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2673 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2023
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2672 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n638, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n606, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3855, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2023, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2022
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2671 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2658
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2670 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n62, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n30, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3693, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2658, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2657
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2669 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2650
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2668 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n638, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n606, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3747, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2650, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2649
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2667 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2013
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2666 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n63, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n31, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3801, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2013, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2012
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2665 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2005
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2664 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n639, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n607, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3855, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2005, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2004
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2663 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2640
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2662 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n63, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n31, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3693, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2640, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2639
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2661 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2632
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2660 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n639, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n607, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3747, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2632, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2631
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2659 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1995
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2658 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n64, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n32, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3801, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1995, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1994
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2657 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1987
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2656 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n640, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n608, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3855, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1987, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1986
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2655 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2622
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2654 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n64, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n32, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3693, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2622, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2621
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2653 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2614
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2652 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n640, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n608, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3747, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2614, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2613
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2651 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3793
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1961
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2650 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n65, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n33, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3801, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1961, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1958
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2649 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3847
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1935
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2648 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n641, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n609, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3855, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1935, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1932
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2647 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1687
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2588
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2646 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n65, B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n33, C2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3693, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2588, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2585
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2645 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3739
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2562
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2644 : OAI221_X1 port map( B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n641, B2 =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750, C1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n609, C2
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3747, A
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2562, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2559
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2643 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3756
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_31_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3753
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2553
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2642 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_31_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1208
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_31_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1205
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3180
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2641 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3756
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_30_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3753
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2520
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2640 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_30_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1208
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_30_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1205
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3147
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2639 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3756
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_29_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3753
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2502
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2638 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_29_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1208
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_29_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1205
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3129
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2637 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3756
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_28_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3753
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2484
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2636 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_28_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1208
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_28_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1205
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3111
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2635 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3756
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_27_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3753
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2466
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2634 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_27_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1208
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_27_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1205
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3093
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2633 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3756
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_26_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3753
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2448
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2632 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_26_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1208
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_26_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1205
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3075
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2631 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3756
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_25_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3753
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2430
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2630 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_25_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1208
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_25_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1205
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3057
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2629 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3756
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_24_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3753
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2412
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2628 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_24_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1208
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_24_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1205
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3039
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2627 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_23_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2394
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2626 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_23_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_23_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3021
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2625 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_22_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2376
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2624 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_22_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_22_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3003
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2623 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_21_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2358
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2622 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_21_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_21_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2985
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2621 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_20_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2340
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2620 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_20_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_20_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2967
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2619 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_19_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2322
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2618 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_19_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_19_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2949
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2617 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_18_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2304
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2616 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_18_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_18_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2931
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2615 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_17_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2286
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2614 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_17_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_17_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2913
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2613 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_16_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2268
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2612 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_16_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_16_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2895
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2611 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_15_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2250
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2610 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_15_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_15_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2877
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2609 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_14_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2232
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2608 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_14_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_14_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2859
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2607 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_13_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2214
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2606 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_13_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_13_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2841
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2605 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3755
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_12_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3752
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2196
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2604 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_12_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1207
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_12_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1204
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2823
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2603 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_11_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2178
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2602 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_11_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_11_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2805
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2601 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_10_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2160
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2600 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_10_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_10_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2787
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2599 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_9_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2142
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2598 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_9_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_9_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2769
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2597 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_8_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2124
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2596 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_8_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_8_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2751
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2595 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_7_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2106
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2594 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_7_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_7_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2733
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2593 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_6_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2088
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2592 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_6_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_6_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2715
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2591 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_5_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2070
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2590 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_5_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_5_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2697
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2589 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_4_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2052
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2588 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_4_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_4_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2679
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2587 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_3_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2034
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2586 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_3_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_3_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2661
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2585 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_2_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2016
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2584 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_2_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_2_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2643
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2583 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_1_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1998
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2582 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_1_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_1_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2625
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2581 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3754
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_0_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n3751
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1977
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2580 : AOI222_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211, A2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_0_port, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n1206
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_0_port, 
                           C1 => dp_id_stage_regfile_DataPath_Physical_RF_n1203
                           , C2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2604
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2579 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_23_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4225, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1261
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2578 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1261, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1130);
   dp_id_stage_regfile_DataPath_Physical_RF_U2577 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_22_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4225, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1260
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2576 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1260, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1131);
   dp_id_stage_regfile_DataPath_Physical_RF_U2575 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_21_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4225, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1259
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2574 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1259, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1132);
   dp_id_stage_regfile_DataPath_Physical_RF_U2573 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_20_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4225, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1258
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2572 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1258, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1133);
   dp_id_stage_regfile_DataPath_Physical_RF_U2571 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_19_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4224, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1257
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2570 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1257, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1134);
   dp_id_stage_regfile_DataPath_Physical_RF_U2569 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_18_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4224, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1256
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2568 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1256, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1135);
   dp_id_stage_regfile_DataPath_Physical_RF_U2567 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_17_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4224, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1255
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2566 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1255, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1136);
   dp_id_stage_regfile_DataPath_Physical_RF_U2565 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_16_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4224, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1254
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2564 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1254, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1137);
   dp_id_stage_regfile_DataPath_Physical_RF_U2563 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_15_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4224, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1253
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2562 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1253, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1138);
   dp_id_stage_regfile_DataPath_Physical_RF_U2561 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_14_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4223, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1252
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2560 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1252, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1139);
   dp_id_stage_regfile_DataPath_Physical_RF_U2559 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_13_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4223, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1251
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2558 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1251, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1140);
   dp_id_stage_regfile_DataPath_Physical_RF_U2557 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4219, A2 
                           => dp_wr_data_id_i_12_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4223, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1250
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2556 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1250, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1141);
   dp_id_stage_regfile_DataPath_Physical_RF_U2555 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_11_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4223, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1249
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2554 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1249, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1142);
   dp_id_stage_regfile_DataPath_Physical_RF_U2553 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_10_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4223, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1248
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2552 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1248, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1143);
   dp_id_stage_regfile_DataPath_Physical_RF_U2551 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_9_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4222, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1247
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2550 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1247, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1144);
   dp_id_stage_regfile_DataPath_Physical_RF_U2549 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_8_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4222, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1246
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2548 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1246, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1145);
   dp_id_stage_regfile_DataPath_Physical_RF_U2547 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_7_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4222, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1245
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2546 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1245, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1146);
   dp_id_stage_regfile_DataPath_Physical_RF_U2545 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_6_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4222, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1244
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2544 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1244, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1147);
   dp_id_stage_regfile_DataPath_Physical_RF_U2543 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_5_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4222, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1243
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2542 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1243, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1148);
   dp_id_stage_regfile_DataPath_Physical_RF_U2541 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_4_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4221, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1242
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2540 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1242, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1149);
   dp_id_stage_regfile_DataPath_Physical_RF_U2539 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_3_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4221, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1241
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2538 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1241, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1150);
   dp_id_stage_regfile_DataPath_Physical_RF_U2537 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_2_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4221, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1240
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2536 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1240, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1151);
   dp_id_stage_regfile_DataPath_Physical_RF_U2535 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_1_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4221, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1239
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2534 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1239, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1152);
   dp_id_stage_regfile_DataPath_Physical_RF_U2533 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4218, A2 
                           => dp_wr_data_id_i_0_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4221, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1237
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2532 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1237, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1153);
   dp_id_stage_regfile_DataPath_Physical_RF_U2531 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4220, A2 
                           => dp_n12, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4227, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1269
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2530 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1269, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1122);
   dp_id_stage_regfile_DataPath_Physical_RF_U2529 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4220, A2 
                           => dp_n10, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4227, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1268
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2528 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1268, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1123);
   dp_id_stage_regfile_DataPath_Physical_RF_U2527 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4220, A2 
                           => dp_wr_data_id_i_29_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4226, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1267
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2526 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1267, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1124);
   dp_id_stage_regfile_DataPath_Physical_RF_U2525 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4220, A2 
                           => dp_wr_data_id_i_28_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4226, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1266
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2524 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1266, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1125);
   dp_id_stage_regfile_DataPath_Physical_RF_U2523 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4220, A2 
                           => dp_n8, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4226, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1265
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2522 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1265, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1126);
   dp_id_stage_regfile_DataPath_Physical_RF_U2521 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4220, A2 
                           => dp_n6, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4226, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1264
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2520 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1264, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1127);
   dp_id_stage_regfile_DataPath_Physical_RF_U2519 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4220, A2 
                           => dp_wr_data_id_i_25_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4226, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1263
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2518 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1263, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1128);
   dp_id_stage_regfile_DataPath_Physical_RF_U2517 : AOI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4220, A2 
                           => dp_wr_data_id_i_24_port, B1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4225, B2 
                           => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1262
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2516 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1262, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1129);
   dp_id_stage_regfile_DataPath_Physical_RF_U2515 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4020, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1677
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2514 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1677, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n490);
   dp_id_stage_regfile_DataPath_Physical_RF_U2513 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4020, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1676
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2512 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1676, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n491);
   dp_id_stage_regfile_DataPath_Physical_RF_U2511 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4020, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1675
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2510 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1675, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n492);
   dp_id_stage_regfile_DataPath_Physical_RF_U2509 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4020, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1674
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2508 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1674, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n493);
   dp_id_stage_regfile_DataPath_Physical_RF_U2507 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4019, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1673
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2506 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1673, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n494);
   dp_id_stage_regfile_DataPath_Physical_RF_U2505 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4019, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1672
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2504 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1672, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n495);
   dp_id_stage_regfile_DataPath_Physical_RF_U2503 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4019, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1671
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2502 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1671, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n496);
   dp_id_stage_regfile_DataPath_Physical_RF_U2501 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4019, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1670
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2500 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1670, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n497);
   dp_id_stage_regfile_DataPath_Physical_RF_U2499 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4019, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1669
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2498 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1669, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n498);
   dp_id_stage_regfile_DataPath_Physical_RF_U2497 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4018, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1668
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2496 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1668, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n499);
   dp_id_stage_regfile_DataPath_Physical_RF_U2495 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4018, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1667
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2494 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1667, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n500);
   dp_id_stage_regfile_DataPath_Physical_RF_U2493 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4018, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1666
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2492 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1666, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n501);
   dp_id_stage_regfile_DataPath_Physical_RF_U2491 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4018, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1665
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2490 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1665, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n502);
   dp_id_stage_regfile_DataPath_Physical_RF_U2489 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4018, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1664
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2488 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1664, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n503);
   dp_id_stage_regfile_DataPath_Physical_RF_U2487 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4017, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1663
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2486 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1663, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n504);
   dp_id_stage_regfile_DataPath_Physical_RF_U2485 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4017, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1662
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2484 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1662, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n505);
   dp_id_stage_regfile_DataPath_Physical_RF_U2483 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4017, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1661
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2482 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1661, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n506);
   dp_id_stage_regfile_DataPath_Physical_RF_U2481 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4017, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1660
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2480 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1660, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n507);
   dp_id_stage_regfile_DataPath_Physical_RF_U2479 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4017, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1659
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2478 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1659, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n508);
   dp_id_stage_regfile_DataPath_Physical_RF_U2477 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4016, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1658
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2476 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1658, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n509);
   dp_id_stage_regfile_DataPath_Physical_RF_U2475 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4016, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1657
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2474 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1657, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n510);
   dp_id_stage_regfile_DataPath_Physical_RF_U2473 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4016, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1656
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2472 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1656, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n511);
   dp_id_stage_regfile_DataPath_Physical_RF_U2471 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4016, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1655
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2470 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1655, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n512);
   dp_id_stage_regfile_DataPath_Physical_RF_U2469 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4016, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1653
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2468 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1653, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n513);
   dp_id_stage_regfile_DataPath_Physical_RF_U2467 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4022, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1685
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2466 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1685, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n482);
   dp_id_stage_regfile_DataPath_Physical_RF_U2465 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4022, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1684
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2464 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1684, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n483);
   dp_id_stage_regfile_DataPath_Physical_RF_U2463 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4021, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1683
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2462 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1683, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n484);
   dp_id_stage_regfile_DataPath_Physical_RF_U2461 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4021, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1682
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2460 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1682, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n485);
   dp_id_stage_regfile_DataPath_Physical_RF_U2459 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4021, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1681
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2458 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1681, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n486);
   dp_id_stage_regfile_DataPath_Physical_RF_U2457 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4021, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1680
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2456 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1680, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n487);
   dp_id_stage_regfile_DataPath_Physical_RF_U2455 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4015, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4021, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1679
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2454 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1679, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n488);
   dp_id_stage_regfile_DataPath_Physical_RF_U2453 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4014, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4020, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1678
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2452 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1678, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n489);
   dp_id_stage_regfile_DataPath_Physical_RF_U2451 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4151, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1374
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2450 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1374, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n906);
   dp_id_stage_regfile_DataPath_Physical_RF_U2449 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4151, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1373
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2448 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1373, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n907);
   dp_id_stage_regfile_DataPath_Physical_RF_U2447 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4151, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1372
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2446 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1372, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n908);
   dp_id_stage_regfile_DataPath_Physical_RF_U2445 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4151, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1371
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2444 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1371, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n909);
   dp_id_stage_regfile_DataPath_Physical_RF_U2443 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4150, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1370
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2442 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1370, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n910);
   dp_id_stage_regfile_DataPath_Physical_RF_U2441 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4150, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1369
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2440 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1369, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n911);
   dp_id_stage_regfile_DataPath_Physical_RF_U2439 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4150, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1368
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2438 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1368, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n912);
   dp_id_stage_regfile_DataPath_Physical_RF_U2437 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4150, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1367
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2436 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1367, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n913);
   dp_id_stage_regfile_DataPath_Physical_RF_U2435 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4150, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1366
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2434 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1366, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n914);
   dp_id_stage_regfile_DataPath_Physical_RF_U2433 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4149, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1365
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2432 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1365, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n915);
   dp_id_stage_regfile_DataPath_Physical_RF_U2431 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4149, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1364
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2430 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1364, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n916);
   dp_id_stage_regfile_DataPath_Physical_RF_U2429 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4149, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1363
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2428 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1363, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n917);
   dp_id_stage_regfile_DataPath_Physical_RF_U2427 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4149, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1362
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2426 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1362, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n918);
   dp_id_stage_regfile_DataPath_Physical_RF_U2425 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4149, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1361
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2424 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1361, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n919);
   dp_id_stage_regfile_DataPath_Physical_RF_U2423 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4148, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1360
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2422 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1360, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n920);
   dp_id_stage_regfile_DataPath_Physical_RF_U2421 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4148, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1359
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2420 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1359, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n921);
   dp_id_stage_regfile_DataPath_Physical_RF_U2419 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4148, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1358
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2418 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1358, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n922);
   dp_id_stage_regfile_DataPath_Physical_RF_U2417 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4148, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1357
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2416 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1357, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n923);
   dp_id_stage_regfile_DataPath_Physical_RF_U2415 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4148, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1356
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2414 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1356, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n924);
   dp_id_stage_regfile_DataPath_Physical_RF_U2413 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4147, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1355
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2412 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1355, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n925);
   dp_id_stage_regfile_DataPath_Physical_RF_U2411 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4147, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1354
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2410 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1354, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n926);
   dp_id_stage_regfile_DataPath_Physical_RF_U2409 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4147, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1353
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2408 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1353, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n927);
   dp_id_stage_regfile_DataPath_Physical_RF_U2407 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4147, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1352
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2406 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1352, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n928);
   dp_id_stage_regfile_DataPath_Physical_RF_U2405 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4147, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1350
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2404 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1350, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n929);
   dp_id_stage_regfile_DataPath_Physical_RF_U2403 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3989, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1713
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2402 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1713, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n394);
   dp_id_stage_regfile_DataPath_Physical_RF_U2401 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3989, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1712
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2400 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1712, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n395);
   dp_id_stage_regfile_DataPath_Physical_RF_U2399 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3989, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1711
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2398 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1711, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n396);
   dp_id_stage_regfile_DataPath_Physical_RF_U2397 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3989, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1710
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2396 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1710, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n397);
   dp_id_stage_regfile_DataPath_Physical_RF_U2395 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3988, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1709
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2394 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1709, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n398);
   dp_id_stage_regfile_DataPath_Physical_RF_U2393 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3988, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1708
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2392 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1708, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n399);
   dp_id_stage_regfile_DataPath_Physical_RF_U2391 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3988, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1707
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2390 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1707, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n400);
   dp_id_stage_regfile_DataPath_Physical_RF_U2389 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3988, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1706
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2388 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1706, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n401);
   dp_id_stage_regfile_DataPath_Physical_RF_U2387 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3988, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1705
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2386 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1705, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n402);
   dp_id_stage_regfile_DataPath_Physical_RF_U2385 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3987, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1704
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2384 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1704, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n403);
   dp_id_stage_regfile_DataPath_Physical_RF_U2383 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3987, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1703
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2382 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1703, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n404);
   dp_id_stage_regfile_DataPath_Physical_RF_U2381 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3987, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1702
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2380 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1702, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n405);
   dp_id_stage_regfile_DataPath_Physical_RF_U2379 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3987, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1701
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2378 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1701, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n406);
   dp_id_stage_regfile_DataPath_Physical_RF_U2377 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3987, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1700
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2376 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1700, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n407);
   dp_id_stage_regfile_DataPath_Physical_RF_U2375 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3986, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1699
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2374 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1699, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n408);
   dp_id_stage_regfile_DataPath_Physical_RF_U2373 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3986, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1698
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2372 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1698, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n409);
   dp_id_stage_regfile_DataPath_Physical_RF_U2371 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3986, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1697
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2370 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1697, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n410);
   dp_id_stage_regfile_DataPath_Physical_RF_U2369 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3986, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1696
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2368 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1696, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n411);
   dp_id_stage_regfile_DataPath_Physical_RF_U2367 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3986, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1695
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2366 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1695, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n412);
   dp_id_stage_regfile_DataPath_Physical_RF_U2365 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3985, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1694
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2364 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1694, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n413);
   dp_id_stage_regfile_DataPath_Physical_RF_U2363 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3985, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1693
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2362 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1693, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n414);
   dp_id_stage_regfile_DataPath_Physical_RF_U2361 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3985, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1692
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2360 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1692, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n415);
   dp_id_stage_regfile_DataPath_Physical_RF_U2359 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3985, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1691
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2358 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1691, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n416);
   dp_id_stage_regfile_DataPath_Physical_RF_U2357 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3985, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1689
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2356 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1689, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n417);
   dp_id_stage_regfile_DataPath_Physical_RF_U2355 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4153, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1382
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2354 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1382, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n898);
   dp_id_stage_regfile_DataPath_Physical_RF_U2353 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4153, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1381
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2352 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1381, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n899);
   dp_id_stage_regfile_DataPath_Physical_RF_U2351 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4152, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1380
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2350 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1380, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n900);
   dp_id_stage_regfile_DataPath_Physical_RF_U2349 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4152, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1379
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2348 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1379, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n901);
   dp_id_stage_regfile_DataPath_Physical_RF_U2347 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4152, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1378
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2346 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1378, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n902);
   dp_id_stage_regfile_DataPath_Physical_RF_U2345 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4152, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1377
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2344 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1377, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n903);
   dp_id_stage_regfile_DataPath_Physical_RF_U2343 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4146, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4152, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1376
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2342 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1376, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n904);
   dp_id_stage_regfile_DataPath_Physical_RF_U2341 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4145, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4151, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1375
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2340 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1375, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n905);
   dp_id_stage_regfile_DataPath_Physical_RF_U2339 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3991, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1721
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2338 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1721, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n386);
   dp_id_stage_regfile_DataPath_Physical_RF_U2337 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3991, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1720
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2336 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1720, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n387);
   dp_id_stage_regfile_DataPath_Physical_RF_U2335 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3990, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1719
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2334 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1719, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n388);
   dp_id_stage_regfile_DataPath_Physical_RF_U2333 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3990, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1718
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2332 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1718, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n389);
   dp_id_stage_regfile_DataPath_Physical_RF_U2331 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3990, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1717
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2330 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1717, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n390);
   dp_id_stage_regfile_DataPath_Physical_RF_U2329 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3990, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1716
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2328 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1716, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n391);
   dp_id_stage_regfile_DataPath_Physical_RF_U2327 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3984, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3990, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1715
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2326 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1715, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n392);
   dp_id_stage_regfile_DataPath_Physical_RF_U2325 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3983, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3989, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1714
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2324 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1714, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n393);
   dp_id_stage_regfile_DataPath_Physical_RF_U2323 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3929, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1848
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2322 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1848, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n202);
   dp_id_stage_regfile_DataPath_Physical_RF_U2321 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3929, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1847
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2320 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1847, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n203);
   dp_id_stage_regfile_DataPath_Physical_RF_U2319 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3929, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1846
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2318 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1846, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n204);
   dp_id_stage_regfile_DataPath_Physical_RF_U2317 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3929, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1845
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2316 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1845, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n205);
   dp_id_stage_regfile_DataPath_Physical_RF_U2315 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3928, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1844
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2314 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1844, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n206);
   dp_id_stage_regfile_DataPath_Physical_RF_U2313 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3928, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1843
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2312 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1843, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n207);
   dp_id_stage_regfile_DataPath_Physical_RF_U2311 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3928, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1842
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2310 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1842, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n208);
   dp_id_stage_regfile_DataPath_Physical_RF_U2309 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3928, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1841
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2308 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1841, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n209);
   dp_id_stage_regfile_DataPath_Physical_RF_U2307 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3928, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1840
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2306 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1840, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n210);
   dp_id_stage_regfile_DataPath_Physical_RF_U2305 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3927, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1839
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2304 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1839, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n211);
   dp_id_stage_regfile_DataPath_Physical_RF_U2303 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3927, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1838
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2302 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1838, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n212);
   dp_id_stage_regfile_DataPath_Physical_RF_U2301 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3927, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1837
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2300 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1837, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n213);
   dp_id_stage_regfile_DataPath_Physical_RF_U2299 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3927, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1836
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2298 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1836, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n214);
   dp_id_stage_regfile_DataPath_Physical_RF_U2297 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3927, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1835
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2296 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1835, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n215);
   dp_id_stage_regfile_DataPath_Physical_RF_U2295 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3926, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1834
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2294 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1834, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n216);
   dp_id_stage_regfile_DataPath_Physical_RF_U2293 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3926, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1833
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2292 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1833, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n217);
   dp_id_stage_regfile_DataPath_Physical_RF_U2291 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3926, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1832
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2290 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1832, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n218);
   dp_id_stage_regfile_DataPath_Physical_RF_U2289 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3926, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1831
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2288 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1831, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n219);
   dp_id_stage_regfile_DataPath_Physical_RF_U2287 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3926, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1830
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2286 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1830, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n220);
   dp_id_stage_regfile_DataPath_Physical_RF_U2285 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3925, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1829
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2284 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1829, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n221);
   dp_id_stage_regfile_DataPath_Physical_RF_U2283 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3925, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1828
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2282 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1828, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n222);
   dp_id_stage_regfile_DataPath_Physical_RF_U2281 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3925, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1827
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2280 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1827, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n223);
   dp_id_stage_regfile_DataPath_Physical_RF_U2279 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3925, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1826
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2278 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1826, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n224);
   dp_id_stage_regfile_DataPath_Physical_RF_U2277 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3925, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1824
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2276 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1824, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n225);
   dp_id_stage_regfile_DataPath_Physical_RF_U2275 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3938, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1814
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2274 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1814, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n234);
   dp_id_stage_regfile_DataPath_Physical_RF_U2273 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3938, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1813
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2272 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1813, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n235);
   dp_id_stage_regfile_DataPath_Physical_RF_U2271 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3938, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1812
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2270 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1812, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n236);
   dp_id_stage_regfile_DataPath_Physical_RF_U2269 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3938, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1811
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2268 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1811, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n237);
   dp_id_stage_regfile_DataPath_Physical_RF_U2267 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3937, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1810
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2266 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1810, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n238);
   dp_id_stage_regfile_DataPath_Physical_RF_U2265 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3937, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1809
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2264 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1809, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n239);
   dp_id_stage_regfile_DataPath_Physical_RF_U2263 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3937, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1808
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2262 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1808, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n240);
   dp_id_stage_regfile_DataPath_Physical_RF_U2261 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3937, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1807
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2260 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1807, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n241);
   dp_id_stage_regfile_DataPath_Physical_RF_U2259 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3937, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1806
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2258 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1806, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n242);
   dp_id_stage_regfile_DataPath_Physical_RF_U2257 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3936, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1805
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2256 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1805, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n243);
   dp_id_stage_regfile_DataPath_Physical_RF_U2255 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3936, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1804
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2254 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1804, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n244);
   dp_id_stage_regfile_DataPath_Physical_RF_U2253 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3936, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1803
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2252 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1803, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n245);
   dp_id_stage_regfile_DataPath_Physical_RF_U2251 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3936, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1802
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2250 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1802, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n246);
   dp_id_stage_regfile_DataPath_Physical_RF_U2249 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3936, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1801
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2248 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1801, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n247);
   dp_id_stage_regfile_DataPath_Physical_RF_U2247 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3935, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1800
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2246 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1800, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n248);
   dp_id_stage_regfile_DataPath_Physical_RF_U2245 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3935, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1799
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2244 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1799, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n249);
   dp_id_stage_regfile_DataPath_Physical_RF_U2243 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3935, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1798
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2242 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1798, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n250);
   dp_id_stage_regfile_DataPath_Physical_RF_U2241 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3935, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1797
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2240 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1797, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n251);
   dp_id_stage_regfile_DataPath_Physical_RF_U2239 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3935, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1796
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2238 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1796, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n252);
   dp_id_stage_regfile_DataPath_Physical_RF_U2237 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3934, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1795
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2236 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1795, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n253);
   dp_id_stage_regfile_DataPath_Physical_RF_U2235 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3934, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1794
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2234 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1794, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n254);
   dp_id_stage_regfile_DataPath_Physical_RF_U2233 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3934, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1793
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2232 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1793, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n255);
   dp_id_stage_regfile_DataPath_Physical_RF_U2231 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3934, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1792
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2230 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1792, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n256);
   dp_id_stage_regfile_DataPath_Physical_RF_U2229 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3934, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1790
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2228 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1790, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n257);
   dp_id_stage_regfile_DataPath_Physical_RF_U2227 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4071, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1576
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2226 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1576, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n650);
   dp_id_stage_regfile_DataPath_Physical_RF_U2225 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4071, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1575
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2224 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1575, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n651);
   dp_id_stage_regfile_DataPath_Physical_RF_U2223 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4071, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1574
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2222 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1574, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n652);
   dp_id_stage_regfile_DataPath_Physical_RF_U2221 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4071, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1573
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2220 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1573, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n653);
   dp_id_stage_regfile_DataPath_Physical_RF_U2219 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4070, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1572
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2218 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1572, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n654);
   dp_id_stage_regfile_DataPath_Physical_RF_U2217 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4070, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1571
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2216 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1571, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n655);
   dp_id_stage_regfile_DataPath_Physical_RF_U2215 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4070, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1570
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2214 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1570, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n656);
   dp_id_stage_regfile_DataPath_Physical_RF_U2213 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4070, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1569
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2212 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1569, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n657);
   dp_id_stage_regfile_DataPath_Physical_RF_U2211 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4070, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1568
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2210 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1568, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n658);
   dp_id_stage_regfile_DataPath_Physical_RF_U2209 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4069, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1567
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2208 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1567, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n659);
   dp_id_stage_regfile_DataPath_Physical_RF_U2207 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4069, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1566
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2206 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1566, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n660);
   dp_id_stage_regfile_DataPath_Physical_RF_U2205 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4069, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1565
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2204 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1565, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n661);
   dp_id_stage_regfile_DataPath_Physical_RF_U2203 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4069, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1564
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2202 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1564, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n662);
   dp_id_stage_regfile_DataPath_Physical_RF_U2201 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4069, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1563
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2200 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1563, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n663);
   dp_id_stage_regfile_DataPath_Physical_RF_U2199 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4068, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1562
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2198 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1562, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n664);
   dp_id_stage_regfile_DataPath_Physical_RF_U2197 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4068, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1561
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2196 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1561, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n665);
   dp_id_stage_regfile_DataPath_Physical_RF_U2195 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4068, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1560
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2194 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1560, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n666);
   dp_id_stage_regfile_DataPath_Physical_RF_U2193 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4068, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1559
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2192 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1559, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n667);
   dp_id_stage_regfile_DataPath_Physical_RF_U2191 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4068, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1558
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2190 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1558, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n668);
   dp_id_stage_regfile_DataPath_Physical_RF_U2189 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4067, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1557
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2188 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1557, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n669);
   dp_id_stage_regfile_DataPath_Physical_RF_U2187 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4067, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1556
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2186 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1556, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n670);
   dp_id_stage_regfile_DataPath_Physical_RF_U2185 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4067, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1555
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2184 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1555, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n671);
   dp_id_stage_regfile_DataPath_Physical_RF_U2183 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4067, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1554
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2182 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1554, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n672);
   dp_id_stage_regfile_DataPath_Physical_RF_U2181 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4067, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1552
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2180 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1552, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n673);
   dp_id_stage_regfile_DataPath_Physical_RF_U2179 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4080, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1543
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2178 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1543, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n682);
   dp_id_stage_regfile_DataPath_Physical_RF_U2177 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4080, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1542
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2176 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1542, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n683);
   dp_id_stage_regfile_DataPath_Physical_RF_U2175 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4080, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1541
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2174 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1541, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n684);
   dp_id_stage_regfile_DataPath_Physical_RF_U2173 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4080, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1540
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2172 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1540, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n685);
   dp_id_stage_regfile_DataPath_Physical_RF_U2171 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4079, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1539
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2170 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1539, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n686);
   dp_id_stage_regfile_DataPath_Physical_RF_U2169 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4079, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1538
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2168 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1538, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n687);
   dp_id_stage_regfile_DataPath_Physical_RF_U2167 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4079, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1537
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2166 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1537, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n688);
   dp_id_stage_regfile_DataPath_Physical_RF_U2165 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4079, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1536
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2164 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1536, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n689);
   dp_id_stage_regfile_DataPath_Physical_RF_U2163 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4079, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1535
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2162 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1535, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n690);
   dp_id_stage_regfile_DataPath_Physical_RF_U2161 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4078, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1534
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2160 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1534, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n691);
   dp_id_stage_regfile_DataPath_Physical_RF_U2159 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4078, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1533
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2158 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1533, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n692);
   dp_id_stage_regfile_DataPath_Physical_RF_U2157 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4078, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1532
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2156 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1532, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n693);
   dp_id_stage_regfile_DataPath_Physical_RF_U2155 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4078, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1531
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2154 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1531, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n694);
   dp_id_stage_regfile_DataPath_Physical_RF_U2153 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4078, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1530
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2152 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1530, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n695);
   dp_id_stage_regfile_DataPath_Physical_RF_U2151 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4077, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1529
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2150 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1529, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n696);
   dp_id_stage_regfile_DataPath_Physical_RF_U2149 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4077, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1528
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2148 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1528, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n697);
   dp_id_stage_regfile_DataPath_Physical_RF_U2147 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4077, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1527
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2146 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1527, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n698);
   dp_id_stage_regfile_DataPath_Physical_RF_U2145 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4077, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1526
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2144 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1526, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n699);
   dp_id_stage_regfile_DataPath_Physical_RF_U2143 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4077, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1525
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2142 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1525, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n700);
   dp_id_stage_regfile_DataPath_Physical_RF_U2141 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4076, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1524
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2140 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1524, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n701);
   dp_id_stage_regfile_DataPath_Physical_RF_U2139 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4076, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1523
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2138 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1523, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n702);
   dp_id_stage_regfile_DataPath_Physical_RF_U2137 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4076, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1522
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2136 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1522, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n703);
   dp_id_stage_regfile_DataPath_Physical_RF_U2135 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4076, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1521
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2134 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1521, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n704);
   dp_id_stage_regfile_DataPath_Physical_RF_U2133 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4076, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1519
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2132 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1519, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n705);
   dp_id_stage_regfile_DataPath_Physical_RF_U2131 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3931, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1856
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2130 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1856, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n194);
   dp_id_stage_regfile_DataPath_Physical_RF_U2129 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3931, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1855
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2128 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1855, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n195);
   dp_id_stage_regfile_DataPath_Physical_RF_U2127 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3930, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1854
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2126 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1854, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n196);
   dp_id_stage_regfile_DataPath_Physical_RF_U2125 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3930, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1853
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2124 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1853, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n197);
   dp_id_stage_regfile_DataPath_Physical_RF_U2123 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3930, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1852
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2122 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1852, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n198);
   dp_id_stage_regfile_DataPath_Physical_RF_U2121 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3930, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1851
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2120 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1851, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n199);
   dp_id_stage_regfile_DataPath_Physical_RF_U2119 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3924, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3930, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1850
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2118 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1850, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n200);
   dp_id_stage_regfile_DataPath_Physical_RF_U2117 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3923, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3929, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1849
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2116 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1849, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n201);
   dp_id_stage_regfile_DataPath_Physical_RF_U2115 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3940, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1822
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2114 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1822, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n226);
   dp_id_stage_regfile_DataPath_Physical_RF_U2113 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3940, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1821
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2112 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1821, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n227);
   dp_id_stage_regfile_DataPath_Physical_RF_U2111 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3939, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1820
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2110 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1820, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n228);
   dp_id_stage_regfile_DataPath_Physical_RF_U2109 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3939, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1819
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2108 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1819, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n229);
   dp_id_stage_regfile_DataPath_Physical_RF_U2107 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3939, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1818
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2106 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1818, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n230);
   dp_id_stage_regfile_DataPath_Physical_RF_U2105 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3939, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1817
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2104 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1817, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n231);
   dp_id_stage_regfile_DataPath_Physical_RF_U2103 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3933, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3939, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1816
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2102 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1816, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n232);
   dp_id_stage_regfile_DataPath_Physical_RF_U2101 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3932, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3938, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1815
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2100 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1815, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n233);
   dp_id_stage_regfile_DataPath_Physical_RF_U2099 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4073, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1584
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2098 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1584, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n642);
   dp_id_stage_regfile_DataPath_Physical_RF_U2097 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4073, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1583
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2096 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1583, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n643);
   dp_id_stage_regfile_DataPath_Physical_RF_U2095 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4072, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1582
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2094 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1582, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n644);
   dp_id_stage_regfile_DataPath_Physical_RF_U2093 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4072, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1581
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2092 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1581, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n645);
   dp_id_stage_regfile_DataPath_Physical_RF_U2091 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4072, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1580
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2090 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1580, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n646);
   dp_id_stage_regfile_DataPath_Physical_RF_U2089 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4072, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1579
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2088 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1579, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n647);
   dp_id_stage_regfile_DataPath_Physical_RF_U2087 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4066, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4072, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1578
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2086 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1578, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n648);
   dp_id_stage_regfile_DataPath_Physical_RF_U2085 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4065, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4071, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1577
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2084 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1577, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n649);
   dp_id_stage_regfile_DataPath_Physical_RF_U2083 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4082, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1551
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2082 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1551, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n674);
   dp_id_stage_regfile_DataPath_Physical_RF_U2081 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4082, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1550
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2080 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1550, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n675);
   dp_id_stage_regfile_DataPath_Physical_RF_U2079 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4081, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1549
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2078 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1549, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n676);
   dp_id_stage_regfile_DataPath_Physical_RF_U2077 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4081, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1548
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2076 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1548, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n677);
   dp_id_stage_regfile_DataPath_Physical_RF_U2075 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4081, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1547
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2074 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1547, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n678);
   dp_id_stage_regfile_DataPath_Physical_RF_U2073 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4081, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1546
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2072 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1546, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n679);
   dp_id_stage_regfile_DataPath_Physical_RF_U2071 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4075, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4081, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1545
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2070 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1545, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n680);
   dp_id_stage_regfile_DataPath_Physical_RF_U2069 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4074, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4080, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1544
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2068 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1544, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n681);
   dp_id_stage_regfile_DataPath_Physical_RF_U2067 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3948, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1781
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2066 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1781, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n266);
   dp_id_stage_regfile_DataPath_Physical_RF_U2065 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3948, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1780
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2064 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1780, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n267);
   dp_id_stage_regfile_DataPath_Physical_RF_U2063 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3948, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1779
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2062 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1779, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n268);
   dp_id_stage_regfile_DataPath_Physical_RF_U2061 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3948, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1778
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2060 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1778, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n269);
   dp_id_stage_regfile_DataPath_Physical_RF_U2059 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3947, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1777
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2058 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1777, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n270);
   dp_id_stage_regfile_DataPath_Physical_RF_U2057 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3947, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1776
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2056 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1776, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n271);
   dp_id_stage_regfile_DataPath_Physical_RF_U2055 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3947, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1775
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2054 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1775, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n272);
   dp_id_stage_regfile_DataPath_Physical_RF_U2053 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3947, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1774
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2052 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1774, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n273);
   dp_id_stage_regfile_DataPath_Physical_RF_U2051 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3947, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1773
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2050 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1773, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n274);
   dp_id_stage_regfile_DataPath_Physical_RF_U2049 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3946, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1772
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2048 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1772, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n275);
   dp_id_stage_regfile_DataPath_Physical_RF_U2047 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3946, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1771
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2046 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1771, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n276);
   dp_id_stage_regfile_DataPath_Physical_RF_U2045 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3942, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3946, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1770
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2044 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1770, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n277);
   dp_id_stage_regfile_DataPath_Physical_RF_U2043 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3946, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1769
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2042 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1769, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n278);
   dp_id_stage_regfile_DataPath_Physical_RF_U2041 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3946, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1768
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2040 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1768, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n279);
   dp_id_stage_regfile_DataPath_Physical_RF_U2039 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3945, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1767
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2038 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1767, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n280);
   dp_id_stage_regfile_DataPath_Physical_RF_U2037 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3945, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1766
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2036 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1766, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n281);
   dp_id_stage_regfile_DataPath_Physical_RF_U2035 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3945, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1765
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2034 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1765, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n282);
   dp_id_stage_regfile_DataPath_Physical_RF_U2033 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3945, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1764
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2032 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1764, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n283);
   dp_id_stage_regfile_DataPath_Physical_RF_U2031 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3945, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1763
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2030 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1763, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n284);
   dp_id_stage_regfile_DataPath_Physical_RF_U2029 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3944, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1762
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2028 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1762, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n285);
   dp_id_stage_regfile_DataPath_Physical_RF_U2027 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3944, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1761
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2026 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1761, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n286);
   dp_id_stage_regfile_DataPath_Physical_RF_U2025 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3944, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1760
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2024 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1760, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n287);
   dp_id_stage_regfile_DataPath_Physical_RF_U2023 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3944, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1759
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2022 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1759, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n288);
   dp_id_stage_regfile_DataPath_Physical_RF_U2021 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3941, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3944, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1757
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2020 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1757, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n289);
   dp_id_stage_regfile_DataPath_Physical_RF_U2019 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4030, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1644
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2018 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1644, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n522);
   dp_id_stage_regfile_DataPath_Physical_RF_U2017 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4030, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1643
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2016 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1643, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n523);
   dp_id_stage_regfile_DataPath_Physical_RF_U2015 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4030, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1642
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2014 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1642, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n524);
   dp_id_stage_regfile_DataPath_Physical_RF_U2013 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4030, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1641
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2012 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1641, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n525);
   dp_id_stage_regfile_DataPath_Physical_RF_U2011 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4029, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1640
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2010 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1640, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n526);
   dp_id_stage_regfile_DataPath_Physical_RF_U2009 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4029, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1639
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2008 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1639, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n527);
   dp_id_stage_regfile_DataPath_Physical_RF_U2007 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4029, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1638
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2006 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1638, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n528);
   dp_id_stage_regfile_DataPath_Physical_RF_U2005 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4029, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1637
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2004 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1637, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n529);
   dp_id_stage_regfile_DataPath_Physical_RF_U2003 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4029, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1636
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2002 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1636, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n530);
   dp_id_stage_regfile_DataPath_Physical_RF_U2001 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4028, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1635
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U2000 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1635, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n531);
   dp_id_stage_regfile_DataPath_Physical_RF_U1999 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4028, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1634
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1998 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1634, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n532);
   dp_id_stage_regfile_DataPath_Physical_RF_U1997 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4024, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4028, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1633
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1996 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1633, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n533);
   dp_id_stage_regfile_DataPath_Physical_RF_U1995 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4028, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1632
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1994 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1632, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n534);
   dp_id_stage_regfile_DataPath_Physical_RF_U1993 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4028, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1631
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1992 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1631, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n535);
   dp_id_stage_regfile_DataPath_Physical_RF_U1991 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4027, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1630
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1990 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1630, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n536);
   dp_id_stage_regfile_DataPath_Physical_RF_U1989 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4027, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1629
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1988 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1629, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n537);
   dp_id_stage_regfile_DataPath_Physical_RF_U1987 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4027, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1628
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1986 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1628, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n538);
   dp_id_stage_regfile_DataPath_Physical_RF_U1985 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4027, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1627
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1984 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1627, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n539);
   dp_id_stage_regfile_DataPath_Physical_RF_U1983 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4027, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1626
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1982 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1626, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n540);
   dp_id_stage_regfile_DataPath_Physical_RF_U1981 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4026, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1625
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1980 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1625, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n541);
   dp_id_stage_regfile_DataPath_Physical_RF_U1979 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4026, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1624
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1978 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1624, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n542);
   dp_id_stage_regfile_DataPath_Physical_RF_U1977 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4026, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1623
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1976 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1623, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n543);
   dp_id_stage_regfile_DataPath_Physical_RF_U1975 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4026, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1622
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1974 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1622, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n544);
   dp_id_stage_regfile_DataPath_Physical_RF_U1973 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4023, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4026, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1620
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1972 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1620, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n545);
   dp_id_stage_regfile_DataPath_Physical_RF_U1971 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4112, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1507
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1970 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1507, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n778);
   dp_id_stage_regfile_DataPath_Physical_RF_U1969 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4112, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1506
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1968 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1506, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n779);
   dp_id_stage_regfile_DataPath_Physical_RF_U1967 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4112, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1505
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1966 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1505, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n780);
   dp_id_stage_regfile_DataPath_Physical_RF_U1965 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4112, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1504
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1964 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1504, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n781);
   dp_id_stage_regfile_DataPath_Physical_RF_U1963 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4111, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1503
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1962 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1503, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n782);
   dp_id_stage_regfile_DataPath_Physical_RF_U1961 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4111, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1502
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1960 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1502, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n783);
   dp_id_stage_regfile_DataPath_Physical_RF_U1959 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4111, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1501
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1958 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1501, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n784);
   dp_id_stage_regfile_DataPath_Physical_RF_U1957 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4111, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1500
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1956 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1500, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n785);
   dp_id_stage_regfile_DataPath_Physical_RF_U1955 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4111, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1499
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1954 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1499, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n786);
   dp_id_stage_regfile_DataPath_Physical_RF_U1953 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4110, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1498
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1952 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1498, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n787);
   dp_id_stage_regfile_DataPath_Physical_RF_U1951 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4110, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1497
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1950 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1497, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n788);
   dp_id_stage_regfile_DataPath_Physical_RF_U1949 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4106, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4110, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1496
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1948 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1496, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n789);
   dp_id_stage_regfile_DataPath_Physical_RF_U1947 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4110, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1495
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1946 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1495, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n790);
   dp_id_stage_regfile_DataPath_Physical_RF_U1945 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4110, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1494
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1944 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1494, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n791);
   dp_id_stage_regfile_DataPath_Physical_RF_U1943 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4109, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1493
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1942 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1493, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n792);
   dp_id_stage_regfile_DataPath_Physical_RF_U1941 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4109, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1492
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1940 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1492, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n793);
   dp_id_stage_regfile_DataPath_Physical_RF_U1939 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4109, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1491
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1938 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1491, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n794);
   dp_id_stage_regfile_DataPath_Physical_RF_U1937 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4109, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1490
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1936 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1490, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n795);
   dp_id_stage_regfile_DataPath_Physical_RF_U1935 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4109, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1489
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1934 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1489, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n796);
   dp_id_stage_regfile_DataPath_Physical_RF_U1933 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4108, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1488
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1932 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1488, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n797);
   dp_id_stage_regfile_DataPath_Physical_RF_U1931 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4108, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1487
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1930 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1487, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n798);
   dp_id_stage_regfile_DataPath_Physical_RF_U1929 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4108, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1486
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1928 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1486, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n799);
   dp_id_stage_regfile_DataPath_Physical_RF_U1927 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4108, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1485
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1926 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1485, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n800);
   dp_id_stage_regfile_DataPath_Physical_RF_U1925 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4105, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4108, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1483
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1924 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1483, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n801);
   dp_id_stage_regfile_DataPath_Physical_RF_U1923 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3888, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1916
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1922 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1916, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n74);
   dp_id_stage_regfile_DataPath_Physical_RF_U1921 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3888, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1915
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1920 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1915, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n75);
   dp_id_stage_regfile_DataPath_Physical_RF_U1919 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3888, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1914
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1918 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1914, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n76);
   dp_id_stage_regfile_DataPath_Physical_RF_U1917 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3888, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1913
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1916 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1913, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n77);
   dp_id_stage_regfile_DataPath_Physical_RF_U1915 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3887, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1912
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1914 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1912, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n78);
   dp_id_stage_regfile_DataPath_Physical_RF_U1913 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3887, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1911
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1912 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1911, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n79);
   dp_id_stage_regfile_DataPath_Physical_RF_U1911 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3887, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1910
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1910 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1910, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n80);
   dp_id_stage_regfile_DataPath_Physical_RF_U1909 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3887, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1909
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1908 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1909, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n81);
   dp_id_stage_regfile_DataPath_Physical_RF_U1907 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3887, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1908
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1906 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1908, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n82);
   dp_id_stage_regfile_DataPath_Physical_RF_U1905 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3886, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1907
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1904 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1907, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n83);
   dp_id_stage_regfile_DataPath_Physical_RF_U1903 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3886, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1906
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1902 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1906, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n84);
   dp_id_stage_regfile_DataPath_Physical_RF_U1901 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3882, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3886, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1905
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1900 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1905, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n85);
   dp_id_stage_regfile_DataPath_Physical_RF_U1899 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3886, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1904
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1898 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1904, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n86);
   dp_id_stage_regfile_DataPath_Physical_RF_U1897 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3886, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1903
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1896 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1903, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n87);
   dp_id_stage_regfile_DataPath_Physical_RF_U1895 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3885, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1902
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1894 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1902, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n88);
   dp_id_stage_regfile_DataPath_Physical_RF_U1893 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3885, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1901
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1892 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1901, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n89);
   dp_id_stage_regfile_DataPath_Physical_RF_U1891 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3885, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1900
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1890 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1900, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n90);
   dp_id_stage_regfile_DataPath_Physical_RF_U1889 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3885, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1899
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1888 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1899, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n91);
   dp_id_stage_regfile_DataPath_Physical_RF_U1887 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3885, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1898
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1886 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1898, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n92);
   dp_id_stage_regfile_DataPath_Physical_RF_U1885 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3884, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1897
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1884 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1897, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n93);
   dp_id_stage_regfile_DataPath_Physical_RF_U1883 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3884, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1896
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1882 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1896, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n94);
   dp_id_stage_regfile_DataPath_Physical_RF_U1881 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3884, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1895
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1880 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1895, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n95);
   dp_id_stage_regfile_DataPath_Physical_RF_U1879 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3884, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1894
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1878 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1894, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n96);
   dp_id_stage_regfile_DataPath_Physical_RF_U1877 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3881, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3884, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1892
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1876 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1892, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n97);
   dp_id_stage_regfile_DataPath_Physical_RF_U1875 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3898, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1883
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1874 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1883, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n106);
   dp_id_stage_regfile_DataPath_Physical_RF_U1873 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3898, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1882
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1872 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1882, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n107);
   dp_id_stage_regfile_DataPath_Physical_RF_U1871 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3898, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1881
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1870 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1881, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n108);
   dp_id_stage_regfile_DataPath_Physical_RF_U1869 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3898, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1880
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1868 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1880, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n109);
   dp_id_stage_regfile_DataPath_Physical_RF_U1867 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3897, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1879
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1866 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1879, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n110);
   dp_id_stage_regfile_DataPath_Physical_RF_U1865 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3897, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1878
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1864 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1878, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n111);
   dp_id_stage_regfile_DataPath_Physical_RF_U1863 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3897, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1877
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1862 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1877, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n112);
   dp_id_stage_regfile_DataPath_Physical_RF_U1861 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3897, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1876
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1860 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1876, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n113);
   dp_id_stage_regfile_DataPath_Physical_RF_U1859 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3897, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1875
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1858 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1875, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n114);
   dp_id_stage_regfile_DataPath_Physical_RF_U1857 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3896, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1874
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1856 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1874, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n115);
   dp_id_stage_regfile_DataPath_Physical_RF_U1855 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3896, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1873
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1854 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1873, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n116);
   dp_id_stage_regfile_DataPath_Physical_RF_U1853 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3892, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3896, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1872
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1852 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1872, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n117);
   dp_id_stage_regfile_DataPath_Physical_RF_U1851 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3896, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1871
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1850 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1871, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n118);
   dp_id_stage_regfile_DataPath_Physical_RF_U1849 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3896, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1870
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1848 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1870, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n119);
   dp_id_stage_regfile_DataPath_Physical_RF_U1847 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3895, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1869
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1846 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1869, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n120);
   dp_id_stage_regfile_DataPath_Physical_RF_U1845 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3895, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1868
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1844 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1868, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n121);
   dp_id_stage_regfile_DataPath_Physical_RF_U1843 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3895, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1867
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1842 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1867, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n122);
   dp_id_stage_regfile_DataPath_Physical_RF_U1841 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3895, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1866
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1840 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1866, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n123);
   dp_id_stage_regfile_DataPath_Physical_RF_U1839 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3895, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1865
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1838 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1865, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n124);
   dp_id_stage_regfile_DataPath_Physical_RF_U1837 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3894, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1864
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1836 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1864, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n125);
   dp_id_stage_regfile_DataPath_Physical_RF_U1835 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3894, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1863
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1834 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1863, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n126);
   dp_id_stage_regfile_DataPath_Physical_RF_U1833 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3894, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1862
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1832 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1862, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n127);
   dp_id_stage_regfile_DataPath_Physical_RF_U1831 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3894, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1861
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1830 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1861, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n128);
   dp_id_stage_regfile_DataPath_Physical_RF_U1829 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3891, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3894, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1859
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1828 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1859, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n129);
   dp_id_stage_regfile_DataPath_Physical_RF_U1827 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3980, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1746
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1826 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1746, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n362);
   dp_id_stage_regfile_DataPath_Physical_RF_U1825 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3980, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1745
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1824 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1745, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n363);
   dp_id_stage_regfile_DataPath_Physical_RF_U1823 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3980, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1744
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1822 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1744, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n364);
   dp_id_stage_regfile_DataPath_Physical_RF_U1821 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3980, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1743
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1820 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1743, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n365);
   dp_id_stage_regfile_DataPath_Physical_RF_U1819 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3979, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1742
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1818 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1742, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n366);
   dp_id_stage_regfile_DataPath_Physical_RF_U1817 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3979, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1741
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1816 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1741, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n367);
   dp_id_stage_regfile_DataPath_Physical_RF_U1815 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3979, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1740
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1814 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1740, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n368);
   dp_id_stage_regfile_DataPath_Physical_RF_U1813 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3979, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1739
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1812 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1739, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n369);
   dp_id_stage_regfile_DataPath_Physical_RF_U1811 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3979, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1738
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1810 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1738, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n370);
   dp_id_stage_regfile_DataPath_Physical_RF_U1809 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3978, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1737
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1808 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1737, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n371);
   dp_id_stage_regfile_DataPath_Physical_RF_U1807 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3978, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1736
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1806 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1736, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n372);
   dp_id_stage_regfile_DataPath_Physical_RF_U1805 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3974, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3978, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1735
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1804 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1735, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n373);
   dp_id_stage_regfile_DataPath_Physical_RF_U1803 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3978, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1734
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1802 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1734, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n374);
   dp_id_stage_regfile_DataPath_Physical_RF_U1801 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3978, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1733
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1800 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1733, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n375);
   dp_id_stage_regfile_DataPath_Physical_RF_U1799 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3977, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1732
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1798 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1732, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n376);
   dp_id_stage_regfile_DataPath_Physical_RF_U1797 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3977, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1731
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1796 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1731, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n377);
   dp_id_stage_regfile_DataPath_Physical_RF_U1795 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3977, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1730
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1794 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1730, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n378);
   dp_id_stage_regfile_DataPath_Physical_RF_U1793 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3977, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1729
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1792 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1729, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n379);
   dp_id_stage_regfile_DataPath_Physical_RF_U1791 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3977, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1728
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1790 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1728, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n380);
   dp_id_stage_regfile_DataPath_Physical_RF_U1789 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3976, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1727
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1788 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1727, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n381);
   dp_id_stage_regfile_DataPath_Physical_RF_U1787 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3976, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1726
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1786 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1726, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n382);
   dp_id_stage_regfile_DataPath_Physical_RF_U1785 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3976, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1725
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1784 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1725, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n383);
   dp_id_stage_regfile_DataPath_Physical_RF_U1783 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3976, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1724
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1782 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1724, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n384);
   dp_id_stage_regfile_DataPath_Physical_RF_U1781 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3973, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3976, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1722
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1780 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1722, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n385);
   dp_id_stage_regfile_DataPath_Physical_RF_U1779 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4132, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1441
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1778 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1441, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n842);
   dp_id_stage_regfile_DataPath_Physical_RF_U1777 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4132, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1440
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1776 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1440, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n843);
   dp_id_stage_regfile_DataPath_Physical_RF_U1775 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4132, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1439
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1774 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1439, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n844);
   dp_id_stage_regfile_DataPath_Physical_RF_U1773 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4132, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1438
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1772 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1438, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n845);
   dp_id_stage_regfile_DataPath_Physical_RF_U1771 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4131, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1437
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1770 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1437, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n846);
   dp_id_stage_regfile_DataPath_Physical_RF_U1769 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4131, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1436
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1768 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1436, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n847);
   dp_id_stage_regfile_DataPath_Physical_RF_U1767 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4131, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1435
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1766 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1435, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n848);
   dp_id_stage_regfile_DataPath_Physical_RF_U1765 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4131, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1434
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1764 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1434, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n849);
   dp_id_stage_regfile_DataPath_Physical_RF_U1763 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4131, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1433
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1762 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1433, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n850);
   dp_id_stage_regfile_DataPath_Physical_RF_U1761 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4130, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1432
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1760 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1432, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n851);
   dp_id_stage_regfile_DataPath_Physical_RF_U1759 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4130, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1431
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1758 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1431, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n852);
   dp_id_stage_regfile_DataPath_Physical_RF_U1757 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4126, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4130, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1430
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1756 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1430, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n853);
   dp_id_stage_regfile_DataPath_Physical_RF_U1755 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4130, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1429
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1754 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1429, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n854);
   dp_id_stage_regfile_DataPath_Physical_RF_U1753 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4130, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1428
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1752 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1428, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n855);
   dp_id_stage_regfile_DataPath_Physical_RF_U1751 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4129, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1427
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1750 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1427, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n856);
   dp_id_stage_regfile_DataPath_Physical_RF_U1749 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4129, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1426
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1748 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1426, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n857);
   dp_id_stage_regfile_DataPath_Physical_RF_U1747 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4129, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1425
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1746 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1425, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n858);
   dp_id_stage_regfile_DataPath_Physical_RF_U1745 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4129, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1424
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1744 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1424, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n859);
   dp_id_stage_regfile_DataPath_Physical_RF_U1743 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4129, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1423
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1742 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1423, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n860);
   dp_id_stage_regfile_DataPath_Physical_RF_U1741 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4128, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1422
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1740 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1422, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n861);
   dp_id_stage_regfile_DataPath_Physical_RF_U1739 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4128, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1421
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1738 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1421, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n862);
   dp_id_stage_regfile_DataPath_Physical_RF_U1737 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4128, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1420
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1736 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1420, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n863);
   dp_id_stage_regfile_DataPath_Physical_RF_U1735 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4128, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1419
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1734 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1419, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n864);
   dp_id_stage_regfile_DataPath_Physical_RF_U1733 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4125, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4128, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1417
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1732 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1417, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n865);
   dp_id_stage_regfile_DataPath_Physical_RF_U1731 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4142, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1408
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1730 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1408, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n874);
   dp_id_stage_regfile_DataPath_Physical_RF_U1729 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4142, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1407
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1728 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1407, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n875);
   dp_id_stage_regfile_DataPath_Physical_RF_U1727 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4142, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1406
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1726 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1406, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n876);
   dp_id_stage_regfile_DataPath_Physical_RF_U1725 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4142, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1405
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1724 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1405, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n877);
   dp_id_stage_regfile_DataPath_Physical_RF_U1723 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4141, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1404
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1722 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1404, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n878);
   dp_id_stage_regfile_DataPath_Physical_RF_U1721 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4141, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1403
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1720 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1403, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n879);
   dp_id_stage_regfile_DataPath_Physical_RF_U1719 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4141, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1402
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1718 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1402, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n880);
   dp_id_stage_regfile_DataPath_Physical_RF_U1717 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4141, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1401
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1716 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1401, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n881);
   dp_id_stage_regfile_DataPath_Physical_RF_U1715 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4141, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1400
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1714 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1400, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n882);
   dp_id_stage_regfile_DataPath_Physical_RF_U1713 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4140, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1399
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1712 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1399, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n883);
   dp_id_stage_regfile_DataPath_Physical_RF_U1711 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4140, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1398
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1710 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1398, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n884);
   dp_id_stage_regfile_DataPath_Physical_RF_U1709 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4136, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4140, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1397
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1708 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1397, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n885);
   dp_id_stage_regfile_DataPath_Physical_RF_U1707 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4140, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1396
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1706 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1396, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n886);
   dp_id_stage_regfile_DataPath_Physical_RF_U1705 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4140, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1395
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1704 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1395, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n887);
   dp_id_stage_regfile_DataPath_Physical_RF_U1703 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4139, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1394
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1702 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1394, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n888);
   dp_id_stage_regfile_DataPath_Physical_RF_U1701 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4139, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1393
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1700 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1393, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n889);
   dp_id_stage_regfile_DataPath_Physical_RF_U1699 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4139, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1392
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1698 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1392, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n890);
   dp_id_stage_regfile_DataPath_Physical_RF_U1697 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4139, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1391
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1696 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1391, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n891);
   dp_id_stage_regfile_DataPath_Physical_RF_U1695 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4139, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1390
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1694 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1390, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n892);
   dp_id_stage_regfile_DataPath_Physical_RF_U1693 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4138, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1389
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1692 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1389, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n893);
   dp_id_stage_regfile_DataPath_Physical_RF_U1691 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4138, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1388
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1690 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1388, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n894);
   dp_id_stage_regfile_DataPath_Physical_RF_U1689 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4138, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1387
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1688 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1387, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n895);
   dp_id_stage_regfile_DataPath_Physical_RF_U1687 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4138, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1386
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1686 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1386, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n896);
   dp_id_stage_regfile_DataPath_Physical_RF_U1685 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4135, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4138, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1384
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1684 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1384, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n897);
   dp_id_stage_regfile_DataPath_Physical_RF_U1683 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4040, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1611
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1682 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1611, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n554);
   dp_id_stage_regfile_DataPath_Physical_RF_U1681 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4040, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1610
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1680 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1610, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n555);
   dp_id_stage_regfile_DataPath_Physical_RF_U1679 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4040, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1609
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1678 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1609, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n556);
   dp_id_stage_regfile_DataPath_Physical_RF_U1677 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4040, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1608
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1676 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1608, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n557);
   dp_id_stage_regfile_DataPath_Physical_RF_U1675 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4039, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1607
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1674 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1607, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n558);
   dp_id_stage_regfile_DataPath_Physical_RF_U1673 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4039, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1606
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1672 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1606, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n559);
   dp_id_stage_regfile_DataPath_Physical_RF_U1671 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4039, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1605
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1670 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1605, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n560);
   dp_id_stage_regfile_DataPath_Physical_RF_U1669 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4039, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1604
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1668 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1604, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n561);
   dp_id_stage_regfile_DataPath_Physical_RF_U1667 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4039, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1603
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1666 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1603, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n562);
   dp_id_stage_regfile_DataPath_Physical_RF_U1665 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4038, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1602
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1664 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1602, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n563);
   dp_id_stage_regfile_DataPath_Physical_RF_U1663 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4038, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1601
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1662 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1601, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n564);
   dp_id_stage_regfile_DataPath_Physical_RF_U1661 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4034, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4038, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1600
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1660 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1600, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n565);
   dp_id_stage_regfile_DataPath_Physical_RF_U1659 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4038, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1599
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1658 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1599, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n566);
   dp_id_stage_regfile_DataPath_Physical_RF_U1657 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4038, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1598
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1656 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1598, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n567);
   dp_id_stage_regfile_DataPath_Physical_RF_U1655 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4037, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1597
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1654 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1597, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n568);
   dp_id_stage_regfile_DataPath_Physical_RF_U1653 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4037, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1596
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1652 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1596, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n569);
   dp_id_stage_regfile_DataPath_Physical_RF_U1651 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4037, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1595
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1650 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1595, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n570);
   dp_id_stage_regfile_DataPath_Physical_RF_U1649 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4037, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1594
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1648 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1594, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n571);
   dp_id_stage_regfile_DataPath_Physical_RF_U1647 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4037, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1593
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1646 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1593, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n572);
   dp_id_stage_regfile_DataPath_Physical_RF_U1645 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4036, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1592
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1644 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1592, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n573);
   dp_id_stage_regfile_DataPath_Physical_RF_U1643 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4036, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1591
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1642 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1591, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n574);
   dp_id_stage_regfile_DataPath_Physical_RF_U1641 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4036, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1590
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1640 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1590, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n575);
   dp_id_stage_regfile_DataPath_Physical_RF_U1639 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4036, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1589
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1638 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1589, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n576);
   dp_id_stage_regfile_DataPath_Physical_RF_U1637 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4033, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4036, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1587
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1636 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1587, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n577);
   dp_id_stage_regfile_DataPath_Physical_RF_U1635 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4122, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1474
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1634 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1474, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n810);
   dp_id_stage_regfile_DataPath_Physical_RF_U1633 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4122, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1473
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1632 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1473, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n811);
   dp_id_stage_regfile_DataPath_Physical_RF_U1631 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4122, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1472
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1630 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1472, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n812);
   dp_id_stage_regfile_DataPath_Physical_RF_U1629 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4122, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1471
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1628 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1471, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n813);
   dp_id_stage_regfile_DataPath_Physical_RF_U1627 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4121, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1470
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1626 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1470, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n814);
   dp_id_stage_regfile_DataPath_Physical_RF_U1625 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4121, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1469
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1624 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1469, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n815);
   dp_id_stage_regfile_DataPath_Physical_RF_U1623 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4121, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1468
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1622 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1468, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n816);
   dp_id_stage_regfile_DataPath_Physical_RF_U1621 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4121, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1467
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1620 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1467, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n817);
   dp_id_stage_regfile_DataPath_Physical_RF_U1619 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4121, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1466
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1618 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1466, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n818);
   dp_id_stage_regfile_DataPath_Physical_RF_U1617 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4120, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1465
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1616 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1465, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n819);
   dp_id_stage_regfile_DataPath_Physical_RF_U1615 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4120, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1464
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1614 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1464, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n820);
   dp_id_stage_regfile_DataPath_Physical_RF_U1613 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4116, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4120, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1463
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1612 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1463, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n821);
   dp_id_stage_regfile_DataPath_Physical_RF_U1611 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4120, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1462
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1610 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1462, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n822);
   dp_id_stage_regfile_DataPath_Physical_RF_U1609 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4120, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1461
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1608 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1461, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n823);
   dp_id_stage_regfile_DataPath_Physical_RF_U1607 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4119, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1460
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1606 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1460, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n824);
   dp_id_stage_regfile_DataPath_Physical_RF_U1605 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4119, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1459
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1604 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1459, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n825);
   dp_id_stage_regfile_DataPath_Physical_RF_U1603 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4119, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1458
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1602 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1458, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n826);
   dp_id_stage_regfile_DataPath_Physical_RF_U1601 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4119, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1457
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1600 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1457, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n827);
   dp_id_stage_regfile_DataPath_Physical_RF_U1599 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4119, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1456
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1598 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1456, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n828);
   dp_id_stage_regfile_DataPath_Physical_RF_U1597 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4118, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1455
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1596 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1455, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n829);
   dp_id_stage_regfile_DataPath_Physical_RF_U1595 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4118, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1454
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1594 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1454, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n830);
   dp_id_stage_regfile_DataPath_Physical_RF_U1593 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4118, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1453
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1592 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1453, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n831);
   dp_id_stage_regfile_DataPath_Physical_RF_U1591 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4118, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1452
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1590 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1452, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n832);
   dp_id_stage_regfile_DataPath_Physical_RF_U1589 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4115, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4118, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1450
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1588 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1450, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n833);
   dp_id_stage_regfile_DataPath_Physical_RF_U1587 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4215, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1296
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1586 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1296, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1098);
   dp_id_stage_regfile_DataPath_Physical_RF_U1585 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4215, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1295
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1584 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1295, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1099);
   dp_id_stage_regfile_DataPath_Physical_RF_U1583 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4215, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1294
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1582 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1294, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1100);
   dp_id_stage_regfile_DataPath_Physical_RF_U1581 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4215, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1293
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1580 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1293, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1101);
   dp_id_stage_regfile_DataPath_Physical_RF_U1579 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4214, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1292
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1578 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1292, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1102);
   dp_id_stage_regfile_DataPath_Physical_RF_U1577 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4214, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1291
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1576 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1291, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1103);
   dp_id_stage_regfile_DataPath_Physical_RF_U1575 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4214, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1290
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1574 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1290, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1104);
   dp_id_stage_regfile_DataPath_Physical_RF_U1573 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4214, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1289
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1572 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1289, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1105);
   dp_id_stage_regfile_DataPath_Physical_RF_U1571 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4214, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1288
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1570 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1288, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1106);
   dp_id_stage_regfile_DataPath_Physical_RF_U1569 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4213, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1287
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1568 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1287, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1107);
   dp_id_stage_regfile_DataPath_Physical_RF_U1567 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4213, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1286
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1566 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1286, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1108);
   dp_id_stage_regfile_DataPath_Physical_RF_U1565 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4209, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4213, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1285
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1564 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1285, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1109);
   dp_id_stage_regfile_DataPath_Physical_RF_U1563 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4213, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1284
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1562 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1284, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1110);
   dp_id_stage_regfile_DataPath_Physical_RF_U1561 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4213, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1283
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1560 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1283, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1111);
   dp_id_stage_regfile_DataPath_Physical_RF_U1559 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4212, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1282
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1558 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1282, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1112);
   dp_id_stage_regfile_DataPath_Physical_RF_U1557 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4212, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1281
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1556 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1281, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1113);
   dp_id_stage_regfile_DataPath_Physical_RF_U1555 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4212, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1280
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1554 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1280, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1114);
   dp_id_stage_regfile_DataPath_Physical_RF_U1553 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4212, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1279
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1552 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1279, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1115);
   dp_id_stage_regfile_DataPath_Physical_RF_U1551 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4212, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1278
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1550 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1278, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1116);
   dp_id_stage_regfile_DataPath_Physical_RF_U1549 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4211, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1277
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1548 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1277, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1117);
   dp_id_stage_regfile_DataPath_Physical_RF_U1547 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4211, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1276
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1546 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1276, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1118);
   dp_id_stage_regfile_DataPath_Physical_RF_U1545 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4211, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1275
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1544 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1275, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1119);
   dp_id_stage_regfile_DataPath_Physical_RF_U1543 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4211, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1274
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1542 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1274, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1120);
   dp_id_stage_regfile_DataPath_Physical_RF_U1541 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4208, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4211, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1272
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1540 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1272, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1121);
   dp_id_stage_regfile_DataPath_Physical_RF_U1539 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_23_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4205, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_23_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1330
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1538 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1330, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1066);
   dp_id_stage_regfile_DataPath_Physical_RF_U1537 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_22_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4205, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_22_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1329
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1536 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1329, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1067);
   dp_id_stage_regfile_DataPath_Physical_RF_U1535 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_21_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4205, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_21_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1328
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1534 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1328, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1068);
   dp_id_stage_regfile_DataPath_Physical_RF_U1533 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_20_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4205, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_20_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1327
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1532 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1327, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1069);
   dp_id_stage_regfile_DataPath_Physical_RF_U1531 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_19_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4204, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_19_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1326
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1530 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1326, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1070);
   dp_id_stage_regfile_DataPath_Physical_RF_U1529 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_18_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4204, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_18_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1325
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1528 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1325, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1071);
   dp_id_stage_regfile_DataPath_Physical_RF_U1527 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_17_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4204, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_17_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1324
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1526 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1324, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1072);
   dp_id_stage_regfile_DataPath_Physical_RF_U1525 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_16_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4204, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_16_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1323
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1524 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1323, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1073);
   dp_id_stage_regfile_DataPath_Physical_RF_U1523 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_15_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4204, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_15_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1322
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1522 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1322, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1074);
   dp_id_stage_regfile_DataPath_Physical_RF_U1521 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_14_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4203, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_14_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1321
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1520 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1321, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1075);
   dp_id_stage_regfile_DataPath_Physical_RF_U1519 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_13_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4203, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_13_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1320
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1518 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1320, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1076);
   dp_id_stage_regfile_DataPath_Physical_RF_U1517 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_12_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4199, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4203, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_12_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1319
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1516 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1319, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1077);
   dp_id_stage_regfile_DataPath_Physical_RF_U1515 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_11_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4203, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_11_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1318
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1514 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1318, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1078);
   dp_id_stage_regfile_DataPath_Physical_RF_U1513 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_10_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4203, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_10_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1317
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1512 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1317, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1079);
   dp_id_stage_regfile_DataPath_Physical_RF_U1511 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_9_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4202, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_9_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1316
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1510 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1316, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1080);
   dp_id_stage_regfile_DataPath_Physical_RF_U1509 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_8_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4202, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_8_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1315
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1508 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1315, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1081);
   dp_id_stage_regfile_DataPath_Physical_RF_U1507 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_7_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4202, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_7_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1314
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1506 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1314, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1082);
   dp_id_stage_regfile_DataPath_Physical_RF_U1505 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_6_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4202, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_6_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1313
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1504 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1313, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1083);
   dp_id_stage_regfile_DataPath_Physical_RF_U1503 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_5_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4202, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1312
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1502 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1312, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1084);
   dp_id_stage_regfile_DataPath_Physical_RF_U1501 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_4_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4201, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1311
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1500 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1311, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1085);
   dp_id_stage_regfile_DataPath_Physical_RF_U1499 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_3_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4201, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1310
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1498 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1310, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1086);
   dp_id_stage_regfile_DataPath_Physical_RF_U1497 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_2_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4201, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1309
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1496 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1309, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1087);
   dp_id_stage_regfile_DataPath_Physical_RF_U1495 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_1_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4201, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1308
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1494 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1308, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1088);
   dp_id_stage_regfile_DataPath_Physical_RF_U1493 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_0_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4198, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4201, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1306
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1492 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1306, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1089);
   dp_id_stage_regfile_DataPath_Physical_RF_U1491 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3943, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3950, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1789
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1490 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1789, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n258);
   dp_id_stage_regfile_DataPath_Physical_RF_U1489 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3943, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3950, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1788
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1488 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1788, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n259);
   dp_id_stage_regfile_DataPath_Physical_RF_U1487 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3943, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3949, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1787
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1486 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1787, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n260);
   dp_id_stage_regfile_DataPath_Physical_RF_U1485 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3943, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3949, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1786
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1484 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1786, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n261);
   dp_id_stage_regfile_DataPath_Physical_RF_U1483 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3943, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3949, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1785
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1482 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1785, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n262);
   dp_id_stage_regfile_DataPath_Physical_RF_U1481 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3943, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3949, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1784
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1480 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1784, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n263);
   dp_id_stage_regfile_DataPath_Physical_RF_U1479 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3943, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3949, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1783
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1478 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1783, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n264);
   dp_id_stage_regfile_DataPath_Physical_RF_U1477 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3943, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3948, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1782
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1476 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1782, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n265);
   dp_id_stage_regfile_DataPath_Physical_RF_U1475 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4025, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4032, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1652
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1474 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1652, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n514);
   dp_id_stage_regfile_DataPath_Physical_RF_U1473 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4025, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4032, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1651
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1472 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1651, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n515);
   dp_id_stage_regfile_DataPath_Physical_RF_U1471 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4025, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4031, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1650
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1470 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1650, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n516);
   dp_id_stage_regfile_DataPath_Physical_RF_U1469 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4025, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4031, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1649
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1468 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1649, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n517);
   dp_id_stage_regfile_DataPath_Physical_RF_U1467 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4025, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4031, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1648
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1466 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1648, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n518);
   dp_id_stage_regfile_DataPath_Physical_RF_U1465 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4025, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4031, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1647
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1464 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1647, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n519);
   dp_id_stage_regfile_DataPath_Physical_RF_U1463 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4025, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4031, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1646
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1462 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1646, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n520);
   dp_id_stage_regfile_DataPath_Physical_RF_U1461 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4025, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4030, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1645
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1460 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1645, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n521);
   dp_id_stage_regfile_DataPath_Physical_RF_U1459 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4107, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4114, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1515
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1458 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1515, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n770);
   dp_id_stage_regfile_DataPath_Physical_RF_U1457 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4107, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4114, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1514
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1456 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1514, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n771);
   dp_id_stage_regfile_DataPath_Physical_RF_U1455 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4107, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4113, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1513
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1454 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1513, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n772);
   dp_id_stage_regfile_DataPath_Physical_RF_U1453 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4107, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4113, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1512
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1452 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1512, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n773);
   dp_id_stage_regfile_DataPath_Physical_RF_U1451 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4107, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4113, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1511
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1450 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1511, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n774);
   dp_id_stage_regfile_DataPath_Physical_RF_U1449 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4107, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4113, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1510
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1448 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1510, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n775);
   dp_id_stage_regfile_DataPath_Physical_RF_U1447 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4107, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4113, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1509
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1446 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1509, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n776);
   dp_id_stage_regfile_DataPath_Physical_RF_U1445 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4107, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4112, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1508
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1444 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1508, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n777);
   dp_id_stage_regfile_DataPath_Physical_RF_U1443 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3883, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3890, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1924
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1442 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1924, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n66);
   dp_id_stage_regfile_DataPath_Physical_RF_U1441 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3883, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3890, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1923
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1440 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1923, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n67);
   dp_id_stage_regfile_DataPath_Physical_RF_U1439 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3883, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3889, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1922
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1438 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1922, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n68);
   dp_id_stage_regfile_DataPath_Physical_RF_U1437 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3883, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3889, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1921
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1436 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1921, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n69);
   dp_id_stage_regfile_DataPath_Physical_RF_U1435 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3883, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3889, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1920
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1434 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1920, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n70);
   dp_id_stage_regfile_DataPath_Physical_RF_U1433 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3883, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3889, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1919
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1432 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1919, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n71);
   dp_id_stage_regfile_DataPath_Physical_RF_U1431 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3883, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3889, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1918
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1430 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1918, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n72);
   dp_id_stage_regfile_DataPath_Physical_RF_U1429 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3883, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3888, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1917
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1428 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1917, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n73);
   dp_id_stage_regfile_DataPath_Physical_RF_U1427 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3893, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3900, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1891
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1426 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1891, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n98);
   dp_id_stage_regfile_DataPath_Physical_RF_U1425 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3893, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3900, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1890
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1424 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1890, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n99);
   dp_id_stage_regfile_DataPath_Physical_RF_U1423 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3893, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3899, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1889
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1422 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1889, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n100);
   dp_id_stage_regfile_DataPath_Physical_RF_U1421 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3893, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3899, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1888
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1420 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1888, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n101);
   dp_id_stage_regfile_DataPath_Physical_RF_U1419 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3893, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3899, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1887
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1418 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1887, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n102);
   dp_id_stage_regfile_DataPath_Physical_RF_U1417 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3893, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3899, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1886
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1416 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1886, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n103);
   dp_id_stage_regfile_DataPath_Physical_RF_U1415 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3893, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3899, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1885
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1414 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1885, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n104);
   dp_id_stage_regfile_DataPath_Physical_RF_U1413 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3893, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3898, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1884
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1412 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1884, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n105);
   dp_id_stage_regfile_DataPath_Physical_RF_U1411 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3975, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3982, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1754
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1410 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1754, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n354);
   dp_id_stage_regfile_DataPath_Physical_RF_U1409 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3975, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3982, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1753
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1408 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1753, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n355);
   dp_id_stage_regfile_DataPath_Physical_RF_U1407 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3975, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3981, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1752
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1406 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1752, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n356);
   dp_id_stage_regfile_DataPath_Physical_RF_U1405 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3975, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3981, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1751
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1404 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1751, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n357);
   dp_id_stage_regfile_DataPath_Physical_RF_U1403 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3975, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3981, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1750
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1402 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1750, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n358);
   dp_id_stage_regfile_DataPath_Physical_RF_U1401 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3975, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3981, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1749
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1400 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1749, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n359);
   dp_id_stage_regfile_DataPath_Physical_RF_U1399 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3975, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3981, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1748
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1398 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1748, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n360);
   dp_id_stage_regfile_DataPath_Physical_RF_U1397 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3975, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3980, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1747
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1396 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1747, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n361);
   dp_id_stage_regfile_DataPath_Physical_RF_U1395 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4127, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4134, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1449
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1394 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1449, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n834);
   dp_id_stage_regfile_DataPath_Physical_RF_U1393 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4127, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4134, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1448
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1392 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1448, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n835);
   dp_id_stage_regfile_DataPath_Physical_RF_U1391 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4127, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4133, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1447
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1390 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1447, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n836);
   dp_id_stage_regfile_DataPath_Physical_RF_U1389 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4127, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4133, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1446
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1388 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1446, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n837);
   dp_id_stage_regfile_DataPath_Physical_RF_U1387 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4127, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4133, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1445
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1386 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1445, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n838);
   dp_id_stage_regfile_DataPath_Physical_RF_U1385 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4127, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4133, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1444
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1384 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1444, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n839);
   dp_id_stage_regfile_DataPath_Physical_RF_U1383 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4127, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4133, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1443
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1382 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1443, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n840);
   dp_id_stage_regfile_DataPath_Physical_RF_U1381 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4127, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4132, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1442
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1380 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1442, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n841);
   dp_id_stage_regfile_DataPath_Physical_RF_U1379 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4137, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4144, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1416
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1378 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1416, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n866);
   dp_id_stage_regfile_DataPath_Physical_RF_U1377 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4137, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4144, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1415
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1376 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1415, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n867);
   dp_id_stage_regfile_DataPath_Physical_RF_U1375 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4137, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4143, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1414
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1374 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1414, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n868);
   dp_id_stage_regfile_DataPath_Physical_RF_U1373 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4137, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4143, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1413
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1372 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1413, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n869);
   dp_id_stage_regfile_DataPath_Physical_RF_U1371 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4137, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4143, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1412
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1370 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1412, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n870);
   dp_id_stage_regfile_DataPath_Physical_RF_U1369 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4137, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4143, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1411
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1368 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1411, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n871);
   dp_id_stage_regfile_DataPath_Physical_RF_U1367 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4137, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4143, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1410
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1366 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1410, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n872);
   dp_id_stage_regfile_DataPath_Physical_RF_U1365 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4137, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4142, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1409
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1364 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1409, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n873);
   dp_id_stage_regfile_DataPath_Physical_RF_U1363 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4035, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4042, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1619
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1362 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1619, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n546);
   dp_id_stage_regfile_DataPath_Physical_RF_U1361 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4035, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4042, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1618
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1360 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1618, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n547);
   dp_id_stage_regfile_DataPath_Physical_RF_U1359 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4035, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4041, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1617
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1358 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1617, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n548);
   dp_id_stage_regfile_DataPath_Physical_RF_U1357 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4035, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4041, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1616
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1356 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1616, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n549);
   dp_id_stage_regfile_DataPath_Physical_RF_U1355 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4035, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4041, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1615
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1354 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1615, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n550);
   dp_id_stage_regfile_DataPath_Physical_RF_U1353 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4035, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4041, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1614
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1352 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1614, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n551);
   dp_id_stage_regfile_DataPath_Physical_RF_U1351 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4035, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4041, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1613
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1350 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1613, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n552);
   dp_id_stage_regfile_DataPath_Physical_RF_U1349 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4035, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4040, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1612
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1348 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1612, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n553);
   dp_id_stage_regfile_DataPath_Physical_RF_U1347 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4117, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4124, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1482
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1346 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1482, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n802);
   dp_id_stage_regfile_DataPath_Physical_RF_U1345 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4117, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4124, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1481
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1344 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1481, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n803);
   dp_id_stage_regfile_DataPath_Physical_RF_U1343 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4117, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4123, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1480
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1342 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1480, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n804);
   dp_id_stage_regfile_DataPath_Physical_RF_U1341 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4117, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4123, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1479
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1340 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1479, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n805);
   dp_id_stage_regfile_DataPath_Physical_RF_U1339 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4117, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4123, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1478
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1338 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1478, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n806);
   dp_id_stage_regfile_DataPath_Physical_RF_U1337 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4117, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4123, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1477
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1336 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1477, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n807);
   dp_id_stage_regfile_DataPath_Physical_RF_U1335 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4117, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4123, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1476
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1334 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1476, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n808);
   dp_id_stage_regfile_DataPath_Physical_RF_U1333 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4117, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4122, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1475
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1332 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1475, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n809);
   dp_id_stage_regfile_DataPath_Physical_RF_U1331 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4210, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4217, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1304
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1330 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1304, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1090);
   dp_id_stage_regfile_DataPath_Physical_RF_U1329 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4210, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4217, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1303
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1328 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1303, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1091);
   dp_id_stage_regfile_DataPath_Physical_RF_U1327 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4210, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4216, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1302
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1326 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1302, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1092);
   dp_id_stage_regfile_DataPath_Physical_RF_U1325 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4210, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4216, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1301
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1324 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1301, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1093);
   dp_id_stage_regfile_DataPath_Physical_RF_U1323 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4210, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4216, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1300
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1322 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1300, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1094);
   dp_id_stage_regfile_DataPath_Physical_RF_U1321 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4210, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4216, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1299
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1320 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1299, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1095);
   dp_id_stage_regfile_DataPath_Physical_RF_U1319 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4210, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4216, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1298
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1318 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1298, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1096);
   dp_id_stage_regfile_DataPath_Physical_RF_U1317 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4210, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4215, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1297
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1316 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1297, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1097);
   dp_id_stage_regfile_DataPath_Physical_RF_U1315 : AOI22_X1 port map( A1 => 
                           dp_n12, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4200, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4207, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_31_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1338
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1314 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1338, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1058);
   dp_id_stage_regfile_DataPath_Physical_RF_U1313 : AOI22_X1 port map( A1 => 
                           dp_n10, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4200, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4207, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_30_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1337
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1312 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1337, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1059);
   dp_id_stage_regfile_DataPath_Physical_RF_U1311 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_29_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4200, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4206, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_29_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1336
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1310 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1336, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1060);
   dp_id_stage_regfile_DataPath_Physical_RF_U1309 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_28_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4200, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4206, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_28_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1335
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1308 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1335, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1061);
   dp_id_stage_regfile_DataPath_Physical_RF_U1307 : AOI22_X1 port map( A1 => 
                           dp_n8, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4200, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4206, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_27_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1334
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1306 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1334, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1062);
   dp_id_stage_regfile_DataPath_Physical_RF_U1305 : AOI22_X1 port map( A1 => 
                           dp_n6, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4200, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4206, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_26_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1333
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1304 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1333, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1063);
   dp_id_stage_regfile_DataPath_Physical_RF_U1303 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_25_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4200, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4206, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_25_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1332
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1302 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1332, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1064);
   dp_id_stage_regfile_DataPath_Physical_RF_U1301 : AOI22_X1 port map( A1 => 
                           dp_wr_data_id_i_24_port, A2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4200, B1 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4205, 
                           B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_24_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1331
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U1300 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1331, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1065);
   dp_id_stage_regfile_DataPath_Physical_RF_U1299 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4178
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n994, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3244);
   dp_id_stage_regfile_DataPath_Physical_RF_U1298 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4178
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n995, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3243);
   dp_id_stage_regfile_DataPath_Physical_RF_U1297 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4178
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n996, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3242);
   dp_id_stage_regfile_DataPath_Physical_RF_U1296 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4178
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n997, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3241);
   dp_id_stage_regfile_DataPath_Physical_RF_U1295 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4179
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n998, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3240);
   dp_id_stage_regfile_DataPath_Physical_RF_U1294 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4179
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n999, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3239);
   dp_id_stage_regfile_DataPath_Physical_RF_U1293 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4179
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1000, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3238);
   dp_id_stage_regfile_DataPath_Physical_RF_U1292 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4179
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1001, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3237);
   dp_id_stage_regfile_DataPath_Physical_RF_U1291 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4180
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1002, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3236);
   dp_id_stage_regfile_DataPath_Physical_RF_U1290 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4180
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1003, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3235);
   dp_id_stage_regfile_DataPath_Physical_RF_U1289 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4180
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1004, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3234);
   dp_id_stage_regfile_DataPath_Physical_RF_U1288 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4180
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1005, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3233);
   dp_id_stage_regfile_DataPath_Physical_RF_U1287 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4181
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1006, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3232);
   dp_id_stage_regfile_DataPath_Physical_RF_U1286 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4181
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1007, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3231);
   dp_id_stage_regfile_DataPath_Physical_RF_U1285 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4181
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1008, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3230);
   dp_id_stage_regfile_DataPath_Physical_RF_U1284 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4181
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1009, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3229);
   dp_id_stage_regfile_DataPath_Physical_RF_U1283 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4182
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1010, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3228);
   dp_id_stage_regfile_DataPath_Physical_RF_U1282 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4182
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1011, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3227);
   dp_id_stage_regfile_DataPath_Physical_RF_U1281 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4182
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1012, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3226);
   dp_id_stage_regfile_DataPath_Physical_RF_U1280 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4182
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1013, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3225);
   dp_id_stage_regfile_DataPath_Physical_RF_U1279 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4183
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1014, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3224);
   dp_id_stage_regfile_DataPath_Physical_RF_U1278 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4183
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1015, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3223);
   dp_id_stage_regfile_DataPath_Physical_RF_U1277 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4183
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1016, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3222);
   dp_id_stage_regfile_DataPath_Physical_RF_U1276 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4183
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1017, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3221);
   dp_id_stage_regfile_DataPath_Physical_RF_U1275 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4184
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1018, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3220);
   dp_id_stage_regfile_DataPath_Physical_RF_U1274 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4184
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1019, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3219);
   dp_id_stage_regfile_DataPath_Physical_RF_U1273 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4184
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1020, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3218);
   dp_id_stage_regfile_DataPath_Physical_RF_U1272 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4184
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1021, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3217);
   dp_id_stage_regfile_DataPath_Physical_RF_U1271 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4185
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1022, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3216);
   dp_id_stage_regfile_DataPath_Physical_RF_U1270 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4185
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1023, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3215);
   dp_id_stage_regfile_DataPath_Physical_RF_U1269 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4185
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1024, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3214);
   dp_id_stage_regfile_DataPath_Physical_RF_U1268 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4185
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1025, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3213);
   dp_id_stage_regfile_DataPath_Physical_RF_U1267 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4173
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n986, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3252);
   dp_id_stage_regfile_DataPath_Physical_RF_U1266 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4173
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n987, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3251);
   dp_id_stage_regfile_DataPath_Physical_RF_U1265 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4173
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n988, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3250);
   dp_id_stage_regfile_DataPath_Physical_RF_U1264 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4173
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n989, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3249);
   dp_id_stage_regfile_DataPath_Physical_RF_U1263 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4174
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n990, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3248);
   dp_id_stage_regfile_DataPath_Physical_RF_U1262 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4174
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n991, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3247);
   dp_id_stage_regfile_DataPath_Physical_RF_U1261 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4174
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n992, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3246);
   dp_id_stage_regfile_DataPath_Physical_RF_U1260 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4174
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n993, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3245);
   dp_id_stage_regfile_DataPath_Physical_RF_U1259 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4162
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n954, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3284);
   dp_id_stage_regfile_DataPath_Physical_RF_U1258 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4162
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n955, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3283);
   dp_id_stage_regfile_DataPath_Physical_RF_U1257 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4162
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n956, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3282);
   dp_id_stage_regfile_DataPath_Physical_RF_U1256 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4162
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n957, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3281);
   dp_id_stage_regfile_DataPath_Physical_RF_U1255 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4163
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n958, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3280);
   dp_id_stage_regfile_DataPath_Physical_RF_U1254 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4163
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n959, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3279);
   dp_id_stage_regfile_DataPath_Physical_RF_U1253 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4163
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n960, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3278);
   dp_id_stage_regfile_DataPath_Physical_RF_U1252 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4163
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n961, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3277);
   dp_id_stage_regfile_DataPath_Physical_RF_U1251 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4167
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n962, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3276);
   dp_id_stage_regfile_DataPath_Physical_RF_U1250 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4167
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n963, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3275);
   dp_id_stage_regfile_DataPath_Physical_RF_U1249 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4167
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n964, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3274);
   dp_id_stage_regfile_DataPath_Physical_RF_U1248 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4167
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n965, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3273);
   dp_id_stage_regfile_DataPath_Physical_RF_U1247 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4168
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n966, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3272);
   dp_id_stage_regfile_DataPath_Physical_RF_U1246 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4168
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n967, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3271);
   dp_id_stage_regfile_DataPath_Physical_RF_U1245 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4168
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n968, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3270);
   dp_id_stage_regfile_DataPath_Physical_RF_U1244 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4168
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n969, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3269);
   dp_id_stage_regfile_DataPath_Physical_RF_U1243 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4169
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n970, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3268);
   dp_id_stage_regfile_DataPath_Physical_RF_U1242 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4169
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n971, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3267);
   dp_id_stage_regfile_DataPath_Physical_RF_U1241 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4169
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n972, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3266);
   dp_id_stage_regfile_DataPath_Physical_RF_U1240 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4169
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n973, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3265);
   dp_id_stage_regfile_DataPath_Physical_RF_U1239 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4170
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n974, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3264);
   dp_id_stage_regfile_DataPath_Physical_RF_U1238 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4170
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n975, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3263);
   dp_id_stage_regfile_DataPath_Physical_RF_U1237 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4170
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n976, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3262);
   dp_id_stage_regfile_DataPath_Physical_RF_U1236 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4170
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n977, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3261);
   dp_id_stage_regfile_DataPath_Physical_RF_U1235 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4171
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n978, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3260);
   dp_id_stage_regfile_DataPath_Physical_RF_U1234 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4171
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n979, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3259);
   dp_id_stage_regfile_DataPath_Physical_RF_U1233 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4171
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n980, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3258);
   dp_id_stage_regfile_DataPath_Physical_RF_U1232 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4171
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n981, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3257);
   dp_id_stage_regfile_DataPath_Physical_RF_U1231 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4172
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n982, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3256);
   dp_id_stage_regfile_DataPath_Physical_RF_U1230 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4172
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n983, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3255);
   dp_id_stage_regfile_DataPath_Physical_RF_U1229 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4172
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n984, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3254);
   dp_id_stage_regfile_DataPath_Physical_RF_U1228 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4172
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n985, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3253);
   dp_id_stage_regfile_DataPath_Physical_RF_U1227 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4156
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n930, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3308);
   dp_id_stage_regfile_DataPath_Physical_RF_U1226 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4156
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n931, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3307);
   dp_id_stage_regfile_DataPath_Physical_RF_U1225 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4156
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n932, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3306);
   dp_id_stage_regfile_DataPath_Physical_RF_U1224 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4156
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n933, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3305);
   dp_id_stage_regfile_DataPath_Physical_RF_U1223 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4157
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n934, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3304);
   dp_id_stage_regfile_DataPath_Physical_RF_U1222 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4157
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n935, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3303);
   dp_id_stage_regfile_DataPath_Physical_RF_U1221 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4157
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n936, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3302);
   dp_id_stage_regfile_DataPath_Physical_RF_U1220 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4157
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n937, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3301);
   dp_id_stage_regfile_DataPath_Physical_RF_U1219 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4158
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n938, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3300);
   dp_id_stage_regfile_DataPath_Physical_RF_U1218 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4158
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n939, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3299);
   dp_id_stage_regfile_DataPath_Physical_RF_U1217 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4158
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n940, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3298);
   dp_id_stage_regfile_DataPath_Physical_RF_U1216 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4158
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n941, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3297);
   dp_id_stage_regfile_DataPath_Physical_RF_U1215 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4159
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n942, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3296);
   dp_id_stage_regfile_DataPath_Physical_RF_U1214 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4159
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n943, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3295);
   dp_id_stage_regfile_DataPath_Physical_RF_U1213 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4159
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n944, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3294);
   dp_id_stage_regfile_DataPath_Physical_RF_U1212 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4159
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n945, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3293);
   dp_id_stage_regfile_DataPath_Physical_RF_U1211 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4160
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n946, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3292);
   dp_id_stage_regfile_DataPath_Physical_RF_U1210 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4160
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n947, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3291);
   dp_id_stage_regfile_DataPath_Physical_RF_U1209 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4160
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n948, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3290);
   dp_id_stage_regfile_DataPath_Physical_RF_U1208 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4160
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n949, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3289);
   dp_id_stage_regfile_DataPath_Physical_RF_U1207 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4161
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n950, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3288);
   dp_id_stage_regfile_DataPath_Physical_RF_U1206 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4161
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n951, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3287);
   dp_id_stage_regfile_DataPath_Physical_RF_U1205 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4161
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n952, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3286);
   dp_id_stage_regfile_DataPath_Physical_RF_U1204 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4161
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n953, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3285);
   dp_id_stage_regfile_DataPath_Physical_RF_U1203 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4011
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n474, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3444);
   dp_id_stage_regfile_DataPath_Physical_RF_U1202 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4011
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n475, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3443);
   dp_id_stage_regfile_DataPath_Physical_RF_U1201 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4011
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n476, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3442);
   dp_id_stage_regfile_DataPath_Physical_RF_U1200 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4011
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n477, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3441);
   dp_id_stage_regfile_DataPath_Physical_RF_U1199 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4012
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n478, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3440);
   dp_id_stage_regfile_DataPath_Physical_RF_U1198 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4012
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n479, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3439);
   dp_id_stage_regfile_DataPath_Physical_RF_U1197 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4012
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n480, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3438);
   dp_id_stage_regfile_DataPath_Physical_RF_U1196 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4012
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n481, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3437);
   dp_id_stage_regfile_DataPath_Physical_RF_U1195 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4000
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n442, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3476);
   dp_id_stage_regfile_DataPath_Physical_RF_U1194 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4000
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n443, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3475);
   dp_id_stage_regfile_DataPath_Physical_RF_U1193 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4000
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n444, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3474);
   dp_id_stage_regfile_DataPath_Physical_RF_U1192 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4000
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n445, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3473);
   dp_id_stage_regfile_DataPath_Physical_RF_U1191 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4001
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n446, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3472);
   dp_id_stage_regfile_DataPath_Physical_RF_U1190 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4001
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n447, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3471);
   dp_id_stage_regfile_DataPath_Physical_RF_U1189 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4001
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n448, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3470);
   dp_id_stage_regfile_DataPath_Physical_RF_U1188 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4001
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n449, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3469);
   dp_id_stage_regfile_DataPath_Physical_RF_U1187 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4005
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n450, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3468);
   dp_id_stage_regfile_DataPath_Physical_RF_U1186 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4005
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n451, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3467);
   dp_id_stage_regfile_DataPath_Physical_RF_U1185 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4005
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n452, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3466);
   dp_id_stage_regfile_DataPath_Physical_RF_U1184 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4005
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n453, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3465);
   dp_id_stage_regfile_DataPath_Physical_RF_U1183 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4006
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n454, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3464);
   dp_id_stage_regfile_DataPath_Physical_RF_U1182 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4006
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n455, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3463);
   dp_id_stage_regfile_DataPath_Physical_RF_U1181 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4006
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n456, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3462);
   dp_id_stage_regfile_DataPath_Physical_RF_U1180 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4006
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n457, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3461);
   dp_id_stage_regfile_DataPath_Physical_RF_U1179 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4007
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n458, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3460);
   dp_id_stage_regfile_DataPath_Physical_RF_U1178 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4007
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n459, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3459);
   dp_id_stage_regfile_DataPath_Physical_RF_U1177 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4007
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n460, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3458);
   dp_id_stage_regfile_DataPath_Physical_RF_U1176 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4007
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n461, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3457);
   dp_id_stage_regfile_DataPath_Physical_RF_U1175 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4008
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n462, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3456);
   dp_id_stage_regfile_DataPath_Physical_RF_U1174 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4008
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n463, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3455);
   dp_id_stage_regfile_DataPath_Physical_RF_U1173 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4008
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n464, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3454);
   dp_id_stage_regfile_DataPath_Physical_RF_U1172 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4008
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n465, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3453);
   dp_id_stage_regfile_DataPath_Physical_RF_U1171 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4009
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n466, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3452);
   dp_id_stage_regfile_DataPath_Physical_RF_U1170 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4009
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n467, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3451);
   dp_id_stage_regfile_DataPath_Physical_RF_U1169 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4009
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n468, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3450);
   dp_id_stage_regfile_DataPath_Physical_RF_U1168 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4009
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n469, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3449);
   dp_id_stage_regfile_DataPath_Physical_RF_U1167 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4010
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n470, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3448);
   dp_id_stage_regfile_DataPath_Physical_RF_U1166 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4010
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n471, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3447);
   dp_id_stage_regfile_DataPath_Physical_RF_U1165 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4010
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n472, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3446);
   dp_id_stage_regfile_DataPath_Physical_RF_U1164 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4010
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n473, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3445);
   dp_id_stage_regfile_DataPath_Physical_RF_U1163 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3994
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n418, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3500);
   dp_id_stage_regfile_DataPath_Physical_RF_U1162 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3994
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n419, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3499);
   dp_id_stage_regfile_DataPath_Physical_RF_U1161 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3994
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n420, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3498);
   dp_id_stage_regfile_DataPath_Physical_RF_U1160 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3994
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n421, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3497);
   dp_id_stage_regfile_DataPath_Physical_RF_U1159 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3995
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n422, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3496);
   dp_id_stage_regfile_DataPath_Physical_RF_U1158 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3995
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n423, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3495);
   dp_id_stage_regfile_DataPath_Physical_RF_U1157 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3995
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n424, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3494);
   dp_id_stage_regfile_DataPath_Physical_RF_U1156 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3995
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n425, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3493);
   dp_id_stage_regfile_DataPath_Physical_RF_U1155 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3996
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n426, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3492);
   dp_id_stage_regfile_DataPath_Physical_RF_U1154 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3996
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n427, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3491);
   dp_id_stage_regfile_DataPath_Physical_RF_U1153 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3996
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n428, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3490);
   dp_id_stage_regfile_DataPath_Physical_RF_U1152 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3996
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n429, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3489);
   dp_id_stage_regfile_DataPath_Physical_RF_U1151 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3997
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n430, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3488);
   dp_id_stage_regfile_DataPath_Physical_RF_U1150 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3997
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n431, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3487);
   dp_id_stage_regfile_DataPath_Physical_RF_U1149 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3997
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n432, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3486);
   dp_id_stage_regfile_DataPath_Physical_RF_U1148 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3997
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n433, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3485);
   dp_id_stage_regfile_DataPath_Physical_RF_U1147 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3998
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n434, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3484);
   dp_id_stage_regfile_DataPath_Physical_RF_U1146 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3998
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n435, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3483);
   dp_id_stage_regfile_DataPath_Physical_RF_U1145 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3998
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n436, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3482);
   dp_id_stage_regfile_DataPath_Physical_RF_U1144 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3998
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n437, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3481);
   dp_id_stage_regfile_DataPath_Physical_RF_U1143 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3999
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n438, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3480);
   dp_id_stage_regfile_DataPath_Physical_RF_U1142 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3999
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n439, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3479);
   dp_id_stage_regfile_DataPath_Physical_RF_U1141 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3999
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n440, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3478);
   dp_id_stage_regfile_DataPath_Physical_RF_U1140 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3999
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n441, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3477);
   dp_id_stage_regfile_DataPath_Physical_RF_U1139 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3909
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n154, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3604);
   dp_id_stage_regfile_DataPath_Physical_RF_U1138 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3909
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n155, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3603);
   dp_id_stage_regfile_DataPath_Physical_RF_U1137 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3909
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n156, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3602);
   dp_id_stage_regfile_DataPath_Physical_RF_U1136 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3909
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n157, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3601);
   dp_id_stage_regfile_DataPath_Physical_RF_U1135 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3910
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n158, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3600);
   dp_id_stage_regfile_DataPath_Physical_RF_U1134 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3910
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n159, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3599);
   dp_id_stage_regfile_DataPath_Physical_RF_U1133 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3910
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n160, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3598);
   dp_id_stage_regfile_DataPath_Physical_RF_U1132 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3910
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n161, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3597);
   dp_id_stage_regfile_DataPath_Physical_RF_U1131 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3920
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n186, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3572);
   dp_id_stage_regfile_DataPath_Physical_RF_U1130 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3920
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n187, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3571);
   dp_id_stage_regfile_DataPath_Physical_RF_U1129 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3920
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n188, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3570);
   dp_id_stage_regfile_DataPath_Physical_RF_U1128 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3920
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n189, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3569);
   dp_id_stage_regfile_DataPath_Physical_RF_U1127 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3921
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n190, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3568);
   dp_id_stage_regfile_DataPath_Physical_RF_U1126 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3921
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n191, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3567);
   dp_id_stage_regfile_DataPath_Physical_RF_U1125 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3921
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n192, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3566);
   dp_id_stage_regfile_DataPath_Physical_RF_U1124 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3921
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n193, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3565);
   dp_id_stage_regfile_DataPath_Physical_RF_U1123 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3903
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n130, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3628);
   dp_id_stage_regfile_DataPath_Physical_RF_U1122 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3903
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n131, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3627);
   dp_id_stage_regfile_DataPath_Physical_RF_U1121 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3903
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n132, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3626);
   dp_id_stage_regfile_DataPath_Physical_RF_U1120 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3903
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n133, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3625);
   dp_id_stage_regfile_DataPath_Physical_RF_U1119 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3904
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n134, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3624);
   dp_id_stage_regfile_DataPath_Physical_RF_U1118 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3904
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n135, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3623);
   dp_id_stage_regfile_DataPath_Physical_RF_U1117 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3904
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n136, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3622);
   dp_id_stage_regfile_DataPath_Physical_RF_U1116 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3904
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n137, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3621);
   dp_id_stage_regfile_DataPath_Physical_RF_U1115 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3905
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n138, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3620);
   dp_id_stage_regfile_DataPath_Physical_RF_U1114 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3905
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n139, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3619);
   dp_id_stage_regfile_DataPath_Physical_RF_U1113 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3905
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n140, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3618);
   dp_id_stage_regfile_DataPath_Physical_RF_U1112 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3905
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n141, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3617);
   dp_id_stage_regfile_DataPath_Physical_RF_U1111 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3906
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n142, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3616);
   dp_id_stage_regfile_DataPath_Physical_RF_U1110 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3906
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n143, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3615);
   dp_id_stage_regfile_DataPath_Physical_RF_U1109 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3906
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n144, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3614);
   dp_id_stage_regfile_DataPath_Physical_RF_U1108 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3906
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n145, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3613);
   dp_id_stage_regfile_DataPath_Physical_RF_U1107 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3907
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n146, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3612);
   dp_id_stage_regfile_DataPath_Physical_RF_U1106 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3907
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n147, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3611);
   dp_id_stage_regfile_DataPath_Physical_RF_U1105 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3907
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n148, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3610);
   dp_id_stage_regfile_DataPath_Physical_RF_U1104 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3907
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n149, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3609);
   dp_id_stage_regfile_DataPath_Physical_RF_U1103 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3908
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n150, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3608);
   dp_id_stage_regfile_DataPath_Physical_RF_U1102 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3908
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n151, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3607);
   dp_id_stage_regfile_DataPath_Physical_RF_U1101 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3908
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n152, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3606);
   dp_id_stage_regfile_DataPath_Physical_RF_U1100 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3908
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n153, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3605);
   dp_id_stage_regfile_DataPath_Physical_RF_U1099 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3914
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n162, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3596);
   dp_id_stage_regfile_DataPath_Physical_RF_U1098 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3914
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n163, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3595);
   dp_id_stage_regfile_DataPath_Physical_RF_U1097 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3914
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n164, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3594);
   dp_id_stage_regfile_DataPath_Physical_RF_U1096 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3914
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n165, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3593);
   dp_id_stage_regfile_DataPath_Physical_RF_U1095 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3915
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n166, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3592);
   dp_id_stage_regfile_DataPath_Physical_RF_U1094 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3915
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n167, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3591);
   dp_id_stage_regfile_DataPath_Physical_RF_U1093 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3915
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n168, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3590);
   dp_id_stage_regfile_DataPath_Physical_RF_U1092 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3915
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n169, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3589);
   dp_id_stage_regfile_DataPath_Physical_RF_U1091 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3916
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n170, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3588);
   dp_id_stage_regfile_DataPath_Physical_RF_U1090 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3916
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n171, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3587);
   dp_id_stage_regfile_DataPath_Physical_RF_U1089 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3916
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n172, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3586);
   dp_id_stage_regfile_DataPath_Physical_RF_U1088 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3916
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n173, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3585);
   dp_id_stage_regfile_DataPath_Physical_RF_U1087 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3917
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n174, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3584);
   dp_id_stage_regfile_DataPath_Physical_RF_U1086 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3917
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n175, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3583);
   dp_id_stage_regfile_DataPath_Physical_RF_U1085 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3917
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n176, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3582);
   dp_id_stage_regfile_DataPath_Physical_RF_U1084 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3917
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n177, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3581);
   dp_id_stage_regfile_DataPath_Physical_RF_U1083 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3918
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n178, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3580);
   dp_id_stage_regfile_DataPath_Physical_RF_U1082 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3918
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n179, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3579);
   dp_id_stage_regfile_DataPath_Physical_RF_U1081 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3918
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n180, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3578);
   dp_id_stage_regfile_DataPath_Physical_RF_U1080 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3918
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n181, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3577);
   dp_id_stage_regfile_DataPath_Physical_RF_U1079 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3919
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n182, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3576);
   dp_id_stage_regfile_DataPath_Physical_RF_U1078 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3919
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n183, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3575);
   dp_id_stage_regfile_DataPath_Physical_RF_U1077 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3919
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n184, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3574);
   dp_id_stage_regfile_DataPath_Physical_RF_U1076 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3919
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n185, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3573);
   dp_id_stage_regfile_DataPath_Physical_RF_U1075 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4091
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n730, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3348);
   dp_id_stage_regfile_DataPath_Physical_RF_U1074 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4091
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n731, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3347);
   dp_id_stage_regfile_DataPath_Physical_RF_U1073 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4091
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n732, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3346);
   dp_id_stage_regfile_DataPath_Physical_RF_U1072 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4091
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n733, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3345);
   dp_id_stage_regfile_DataPath_Physical_RF_U1071 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4092
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n734, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3344);
   dp_id_stage_regfile_DataPath_Physical_RF_U1070 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4092
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n735, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3343);
   dp_id_stage_regfile_DataPath_Physical_RF_U1069 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4092
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n736, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3342);
   dp_id_stage_regfile_DataPath_Physical_RF_U1068 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4092
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n737, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3341);
   dp_id_stage_regfile_DataPath_Physical_RF_U1067 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4102
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n762, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3316);
   dp_id_stage_regfile_DataPath_Physical_RF_U1066 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4102
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n763, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3315);
   dp_id_stage_regfile_DataPath_Physical_RF_U1065 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4102
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n764, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3314);
   dp_id_stage_regfile_DataPath_Physical_RF_U1064 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4102
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n765, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3313);
   dp_id_stage_regfile_DataPath_Physical_RF_U1063 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4103
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n766, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3312);
   dp_id_stage_regfile_DataPath_Physical_RF_U1062 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4103
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n767, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3311);
   dp_id_stage_regfile_DataPath_Physical_RF_U1061 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4103
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n768, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3310);
   dp_id_stage_regfile_DataPath_Physical_RF_U1060 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4103
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n769, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3309);
   dp_id_stage_regfile_DataPath_Physical_RF_U1059 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4085
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n706, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3372);
   dp_id_stage_regfile_DataPath_Physical_RF_U1058 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4085
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n707, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3371);
   dp_id_stage_regfile_DataPath_Physical_RF_U1057 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4085
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n708, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3370);
   dp_id_stage_regfile_DataPath_Physical_RF_U1056 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4085
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n709, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3369);
   dp_id_stage_regfile_DataPath_Physical_RF_U1055 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4086
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n710, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3368);
   dp_id_stage_regfile_DataPath_Physical_RF_U1054 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4086
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n711, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3367);
   dp_id_stage_regfile_DataPath_Physical_RF_U1053 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4086
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n712, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3366);
   dp_id_stage_regfile_DataPath_Physical_RF_U1052 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4086
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n713, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3365);
   dp_id_stage_regfile_DataPath_Physical_RF_U1051 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4087
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n714, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3364);
   dp_id_stage_regfile_DataPath_Physical_RF_U1050 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4087
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n715, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3363);
   dp_id_stage_regfile_DataPath_Physical_RF_U1049 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4087
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n716, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3362);
   dp_id_stage_regfile_DataPath_Physical_RF_U1048 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4087
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n717, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3361);
   dp_id_stage_regfile_DataPath_Physical_RF_U1047 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4088
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n718, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3360);
   dp_id_stage_regfile_DataPath_Physical_RF_U1046 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4088
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n719, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3359);
   dp_id_stage_regfile_DataPath_Physical_RF_U1045 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4088
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n720, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3358);
   dp_id_stage_regfile_DataPath_Physical_RF_U1044 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4088
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n721, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3357);
   dp_id_stage_regfile_DataPath_Physical_RF_U1043 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4089
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n722, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3356);
   dp_id_stage_regfile_DataPath_Physical_RF_U1042 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4089
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n723, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3355);
   dp_id_stage_regfile_DataPath_Physical_RF_U1041 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4089
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n724, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3354);
   dp_id_stage_regfile_DataPath_Physical_RF_U1040 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4089
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n725, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3353);
   dp_id_stage_regfile_DataPath_Physical_RF_U1039 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4090
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n726, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3352);
   dp_id_stage_regfile_DataPath_Physical_RF_U1038 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4090
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n727, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3351);
   dp_id_stage_regfile_DataPath_Physical_RF_U1037 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4090
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n728, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3350);
   dp_id_stage_regfile_DataPath_Physical_RF_U1036 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4090
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n729, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3349);
   dp_id_stage_regfile_DataPath_Physical_RF_U1035 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4096
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n738, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3340);
   dp_id_stage_regfile_DataPath_Physical_RF_U1034 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4096
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n739, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3339);
   dp_id_stage_regfile_DataPath_Physical_RF_U1033 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4096
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n740, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3338);
   dp_id_stage_regfile_DataPath_Physical_RF_U1032 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4096
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n741, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3337);
   dp_id_stage_regfile_DataPath_Physical_RF_U1031 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4097
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n742, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3336);
   dp_id_stage_regfile_DataPath_Physical_RF_U1030 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4097
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n743, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3335);
   dp_id_stage_regfile_DataPath_Physical_RF_U1029 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4097
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n744, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3334);
   dp_id_stage_regfile_DataPath_Physical_RF_U1028 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4097
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n745, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3333);
   dp_id_stage_regfile_DataPath_Physical_RF_U1027 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4098
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n746, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3332);
   dp_id_stage_regfile_DataPath_Physical_RF_U1026 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4098
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n747, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3331);
   dp_id_stage_regfile_DataPath_Physical_RF_U1025 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4098
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n748, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3330);
   dp_id_stage_regfile_DataPath_Physical_RF_U1024 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4098
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n749, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3329);
   dp_id_stage_regfile_DataPath_Physical_RF_U1023 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4099
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n750, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3328);
   dp_id_stage_regfile_DataPath_Physical_RF_U1022 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4099
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n751, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3327);
   dp_id_stage_regfile_DataPath_Physical_RF_U1021 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4099
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n752, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3326);
   dp_id_stage_regfile_DataPath_Physical_RF_U1020 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4099
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n753, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3325);
   dp_id_stage_regfile_DataPath_Physical_RF_U1019 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4100
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n754, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3324);
   dp_id_stage_regfile_DataPath_Physical_RF_U1018 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4100
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n755, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3323);
   dp_id_stage_regfile_DataPath_Physical_RF_U1017 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4100
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n756, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3322);
   dp_id_stage_regfile_DataPath_Physical_RF_U1016 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4100
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n757, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3321);
   dp_id_stage_regfile_DataPath_Physical_RF_U1015 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4101
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n758, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3320);
   dp_id_stage_regfile_DataPath_Physical_RF_U1014 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4101
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n759, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3319);
   dp_id_stage_regfile_DataPath_Physical_RF_U1013 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4101
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n760, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3318);
   dp_id_stage_regfile_DataPath_Physical_RF_U1012 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4101
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n761, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3317);
   dp_id_stage_regfile_DataPath_Physical_RF_U1011 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3867
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n26
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3668);
   dp_id_stage_regfile_DataPath_Physical_RF_U1010 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3867
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n27
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3667);
   dp_id_stage_regfile_DataPath_Physical_RF_U1009 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3867
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n28
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3666);
   dp_id_stage_regfile_DataPath_Physical_RF_U1008 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3867
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n29
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3665);
   dp_id_stage_regfile_DataPath_Physical_RF_U1007 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3868
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n30
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3664);
   dp_id_stage_regfile_DataPath_Physical_RF_U1006 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3868
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n31
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3663);
   dp_id_stage_regfile_DataPath_Physical_RF_U1005 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3868
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n32
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3662);
   dp_id_stage_regfile_DataPath_Physical_RF_U1004 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3868
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n33
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3661);
   dp_id_stage_regfile_DataPath_Physical_RF_U1003 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3970
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n346, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3508);
   dp_id_stage_regfile_DataPath_Physical_RF_U1002 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3970
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n347, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3507);
   dp_id_stage_regfile_DataPath_Physical_RF_U1001 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3970
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n348, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3506);
   dp_id_stage_regfile_DataPath_Physical_RF_U1000 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3970
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n349, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3505);
   dp_id_stage_regfile_DataPath_Physical_RF_U999 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3971
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n350, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3504);
   dp_id_stage_regfile_DataPath_Physical_RF_U998 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3971
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n351, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3503);
   dp_id_stage_regfile_DataPath_Physical_RF_U997 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3971
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n352, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3502);
   dp_id_stage_regfile_DataPath_Physical_RF_U996 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3971
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n353, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3501);
   dp_id_stage_regfile_DataPath_Physical_RF_U995 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4051
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n602, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3412);
   dp_id_stage_regfile_DataPath_Physical_RF_U994 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4051
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n603, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3411);
   dp_id_stage_regfile_DataPath_Physical_RF_U993 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4051
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n604, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3410);
   dp_id_stage_regfile_DataPath_Physical_RF_U992 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4051
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n605, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3409);
   dp_id_stage_regfile_DataPath_Physical_RF_U991 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4052
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n606, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3408);
   dp_id_stage_regfile_DataPath_Physical_RF_U990 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4052
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n607, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3407);
   dp_id_stage_regfile_DataPath_Physical_RF_U989 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4052
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n608, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3406);
   dp_id_stage_regfile_DataPath_Physical_RF_U988 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4052
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n609, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3405);
   dp_id_stage_regfile_DataPath_Physical_RF_U987 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4062
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n634, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3380);
   dp_id_stage_regfile_DataPath_Physical_RF_U986 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4062
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n635, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3379);
   dp_id_stage_regfile_DataPath_Physical_RF_U985 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4062
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n636, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3378);
   dp_id_stage_regfile_DataPath_Physical_RF_U984 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4062
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n637, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3377);
   dp_id_stage_regfile_DataPath_Physical_RF_U983 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4063
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n638, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3376);
   dp_id_stage_regfile_DataPath_Physical_RF_U982 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4063
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n639, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3375);
   dp_id_stage_regfile_DataPath_Physical_RF_U981 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4063
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n640, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3374);
   dp_id_stage_regfile_DataPath_Physical_RF_U980 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4063
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n641, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3373);
   dp_id_stage_regfile_DataPath_Physical_RF_U979 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3878
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n58
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3636);
   dp_id_stage_regfile_DataPath_Physical_RF_U978 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3878
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n59
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3635);
   dp_id_stage_regfile_DataPath_Physical_RF_U977 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3878
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n60
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3634);
   dp_id_stage_regfile_DataPath_Physical_RF_U976 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3878
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n61
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3633);
   dp_id_stage_regfile_DataPath_Physical_RF_U975 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3879
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n62
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3632);
   dp_id_stage_regfile_DataPath_Physical_RF_U974 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3879
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n63
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3631);
   dp_id_stage_regfile_DataPath_Physical_RF_U973 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3879
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n64
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3630);
   dp_id_stage_regfile_DataPath_Physical_RF_U972 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3879
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n65
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3629);
   dp_id_stage_regfile_DataPath_Physical_RF_U971 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3959
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n314, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3540);
   dp_id_stage_regfile_DataPath_Physical_RF_U970 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3959
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n315, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3539);
   dp_id_stage_regfile_DataPath_Physical_RF_U969 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3959
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n316, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3538);
   dp_id_stage_regfile_DataPath_Physical_RF_U968 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3959
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n317, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3537);
   dp_id_stage_regfile_DataPath_Physical_RF_U967 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3960
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n318, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3536);
   dp_id_stage_regfile_DataPath_Physical_RF_U966 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3960
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n319, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3535);
   dp_id_stage_regfile_DataPath_Physical_RF_U965 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3960
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n320, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3534);
   dp_id_stage_regfile_DataPath_Physical_RF_U964 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3960
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n321, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3533);
   dp_id_stage_regfile_DataPath_Physical_RF_U963 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4195
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1050, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3188);
   dp_id_stage_regfile_DataPath_Physical_RF_U962 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4195
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1051, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3187);
   dp_id_stage_regfile_DataPath_Physical_RF_U961 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4195
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1052, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3186);
   dp_id_stage_regfile_DataPath_Physical_RF_U960 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4195
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1053, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3185);
   dp_id_stage_regfile_DataPath_Physical_RF_U959 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4196
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1054, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3184);
   dp_id_stage_regfile_DataPath_Physical_RF_U958 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4196
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1055, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3183);
   dp_id_stage_regfile_DataPath_Physical_RF_U957 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4196
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1056, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3182);
   dp_id_stage_regfile_DataPath_Physical_RF_U956 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4196
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1057, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3181);
   dp_id_stage_regfile_DataPath_Physical_RF_U955 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3861
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n2,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3692
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U954 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3861
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n3,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3691
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U953 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3861
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n4,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3690
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U952 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3861
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n5,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3689
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U951 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3862
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n6,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3688
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U950 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3862
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n7,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3687
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U949 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3862
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n8,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3686
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U948 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3862
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n9,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3685
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U947 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3863
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n10
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3684);
   dp_id_stage_regfile_DataPath_Physical_RF_U946 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3863
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n11
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3683);
   dp_id_stage_regfile_DataPath_Physical_RF_U945 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3863
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n12
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3682);
   dp_id_stage_regfile_DataPath_Physical_RF_U944 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3863
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n13
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3681);
   dp_id_stage_regfile_DataPath_Physical_RF_U943 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3864
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n14
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3680);
   dp_id_stage_regfile_DataPath_Physical_RF_U942 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3864
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n15
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3679);
   dp_id_stage_regfile_DataPath_Physical_RF_U941 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3864
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n16
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3678);
   dp_id_stage_regfile_DataPath_Physical_RF_U940 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3864
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n17
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3677);
   dp_id_stage_regfile_DataPath_Physical_RF_U939 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3865
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n18
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3676);
   dp_id_stage_regfile_DataPath_Physical_RF_U938 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3865
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n19
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3675);
   dp_id_stage_regfile_DataPath_Physical_RF_U937 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3865
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n20
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3674);
   dp_id_stage_regfile_DataPath_Physical_RF_U936 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3865
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n21
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3673);
   dp_id_stage_regfile_DataPath_Physical_RF_U935 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3866
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n22
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3672);
   dp_id_stage_regfile_DataPath_Physical_RF_U934 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3866
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n23
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3671);
   dp_id_stage_regfile_DataPath_Physical_RF_U933 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3866
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n24
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3670);
   dp_id_stage_regfile_DataPath_Physical_RF_U932 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3866
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n25
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3669);
   dp_id_stage_regfile_DataPath_Physical_RF_U931 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3964
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n322, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3532);
   dp_id_stage_regfile_DataPath_Physical_RF_U930 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3964
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n323, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3531);
   dp_id_stage_regfile_DataPath_Physical_RF_U929 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3964
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n324, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3530);
   dp_id_stage_regfile_DataPath_Physical_RF_U928 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3964
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n325, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3529);
   dp_id_stage_regfile_DataPath_Physical_RF_U927 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3965
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n326, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3528);
   dp_id_stage_regfile_DataPath_Physical_RF_U926 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3965
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n327, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3527);
   dp_id_stage_regfile_DataPath_Physical_RF_U925 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3965
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n328, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3526);
   dp_id_stage_regfile_DataPath_Physical_RF_U924 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3965
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n329, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3525);
   dp_id_stage_regfile_DataPath_Physical_RF_U923 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3966
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n330, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3524);
   dp_id_stage_regfile_DataPath_Physical_RF_U922 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3966
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n331, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3523);
   dp_id_stage_regfile_DataPath_Physical_RF_U921 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3966
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n332, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3522);
   dp_id_stage_regfile_DataPath_Physical_RF_U920 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3966
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n333, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3521);
   dp_id_stage_regfile_DataPath_Physical_RF_U919 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3967
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n334, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3520);
   dp_id_stage_regfile_DataPath_Physical_RF_U918 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3967
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n335, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3519);
   dp_id_stage_regfile_DataPath_Physical_RF_U917 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3967
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n336, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3518);
   dp_id_stage_regfile_DataPath_Physical_RF_U916 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3967
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n337, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3517);
   dp_id_stage_regfile_DataPath_Physical_RF_U915 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3968
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n338, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3516);
   dp_id_stage_regfile_DataPath_Physical_RF_U914 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3968
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n339, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3515);
   dp_id_stage_regfile_DataPath_Physical_RF_U913 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3968
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n340, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3514);
   dp_id_stage_regfile_DataPath_Physical_RF_U912 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3968
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n341, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3513);
   dp_id_stage_regfile_DataPath_Physical_RF_U911 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3969
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n342, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3512);
   dp_id_stage_regfile_DataPath_Physical_RF_U910 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3969
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n343, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3511);
   dp_id_stage_regfile_DataPath_Physical_RF_U909 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3969
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n344, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3510);
   dp_id_stage_regfile_DataPath_Physical_RF_U908 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3969
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n345, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3509);
   dp_id_stage_regfile_DataPath_Physical_RF_U907 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4045
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n578, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3436);
   dp_id_stage_regfile_DataPath_Physical_RF_U906 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4045
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n579, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3435);
   dp_id_stage_regfile_DataPath_Physical_RF_U905 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4045
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n580, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3434);
   dp_id_stage_regfile_DataPath_Physical_RF_U904 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4045
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n581, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3433);
   dp_id_stage_regfile_DataPath_Physical_RF_U903 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4046
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n582, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3432);
   dp_id_stage_regfile_DataPath_Physical_RF_U902 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4046
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n583, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3431);
   dp_id_stage_regfile_DataPath_Physical_RF_U901 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4046
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n584, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3430);
   dp_id_stage_regfile_DataPath_Physical_RF_U900 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4046
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n585, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3429);
   dp_id_stage_regfile_DataPath_Physical_RF_U899 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4047
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n586, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3428);
   dp_id_stage_regfile_DataPath_Physical_RF_U898 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4047
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n587, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3427);
   dp_id_stage_regfile_DataPath_Physical_RF_U897 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4047
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n588, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3426);
   dp_id_stage_regfile_DataPath_Physical_RF_U896 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4047
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n589, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3425);
   dp_id_stage_regfile_DataPath_Physical_RF_U895 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4048
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n590, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3424);
   dp_id_stage_regfile_DataPath_Physical_RF_U894 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4048
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n591, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3423);
   dp_id_stage_regfile_DataPath_Physical_RF_U893 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4048
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n592, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3422);
   dp_id_stage_regfile_DataPath_Physical_RF_U892 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4048
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n593, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3421);
   dp_id_stage_regfile_DataPath_Physical_RF_U891 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4049
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n594, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3420);
   dp_id_stage_regfile_DataPath_Physical_RF_U890 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4049
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n595, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3419);
   dp_id_stage_regfile_DataPath_Physical_RF_U889 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4049
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n596, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3418);
   dp_id_stage_regfile_DataPath_Physical_RF_U888 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4049
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n597, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3417);
   dp_id_stage_regfile_DataPath_Physical_RF_U887 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4050
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n598, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3416);
   dp_id_stage_regfile_DataPath_Physical_RF_U886 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4050
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n599, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3415);
   dp_id_stage_regfile_DataPath_Physical_RF_U885 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4050
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n600, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3414);
   dp_id_stage_regfile_DataPath_Physical_RF_U884 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4050
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n601, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3413);
   dp_id_stage_regfile_DataPath_Physical_RF_U883 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4056
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n610, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3404);
   dp_id_stage_regfile_DataPath_Physical_RF_U882 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4056
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n611, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3403);
   dp_id_stage_regfile_DataPath_Physical_RF_U881 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4056
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n612, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3402);
   dp_id_stage_regfile_DataPath_Physical_RF_U880 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4056
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n613, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3401);
   dp_id_stage_regfile_DataPath_Physical_RF_U879 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4057
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n614, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3400);
   dp_id_stage_regfile_DataPath_Physical_RF_U878 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4057
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n615, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3399);
   dp_id_stage_regfile_DataPath_Physical_RF_U877 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4057
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n616, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3398);
   dp_id_stage_regfile_DataPath_Physical_RF_U876 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4057
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n617, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3397);
   dp_id_stage_regfile_DataPath_Physical_RF_U875 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4058
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n618, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3396);
   dp_id_stage_regfile_DataPath_Physical_RF_U874 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4058
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n619, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3395);
   dp_id_stage_regfile_DataPath_Physical_RF_U873 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4058
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n620, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3394);
   dp_id_stage_regfile_DataPath_Physical_RF_U872 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4058
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n621, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3393);
   dp_id_stage_regfile_DataPath_Physical_RF_U871 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4059
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n622, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3392);
   dp_id_stage_regfile_DataPath_Physical_RF_U870 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4059
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n623, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3391);
   dp_id_stage_regfile_DataPath_Physical_RF_U869 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4059
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n624, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3390);
   dp_id_stage_regfile_DataPath_Physical_RF_U868 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4059
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n625, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3389);
   dp_id_stage_regfile_DataPath_Physical_RF_U867 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4060
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n626, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3388);
   dp_id_stage_regfile_DataPath_Physical_RF_U866 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4060
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n627, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3387);
   dp_id_stage_regfile_DataPath_Physical_RF_U865 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4060
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n628, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3386);
   dp_id_stage_regfile_DataPath_Physical_RF_U864 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4060
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n629, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3385);
   dp_id_stage_regfile_DataPath_Physical_RF_U863 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4061
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n630, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3384);
   dp_id_stage_regfile_DataPath_Physical_RF_U862 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4061
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n631, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3383);
   dp_id_stage_regfile_DataPath_Physical_RF_U861 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4061
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n632, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3382);
   dp_id_stage_regfile_DataPath_Physical_RF_U860 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4061
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n633, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3381);
   dp_id_stage_regfile_DataPath_Physical_RF_U859 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3872
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n34
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3660);
   dp_id_stage_regfile_DataPath_Physical_RF_U858 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3872
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n35
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3659);
   dp_id_stage_regfile_DataPath_Physical_RF_U857 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3872
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n36
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3658);
   dp_id_stage_regfile_DataPath_Physical_RF_U856 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3872
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n37
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3657);
   dp_id_stage_regfile_DataPath_Physical_RF_U855 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3873
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n38
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3656);
   dp_id_stage_regfile_DataPath_Physical_RF_U854 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3873
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n39
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3655);
   dp_id_stage_regfile_DataPath_Physical_RF_U853 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3873
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n40
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3654);
   dp_id_stage_regfile_DataPath_Physical_RF_U852 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3873
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n41
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3653);
   dp_id_stage_regfile_DataPath_Physical_RF_U851 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3874
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n42
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3652);
   dp_id_stage_regfile_DataPath_Physical_RF_U850 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3874
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n43
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3651);
   dp_id_stage_regfile_DataPath_Physical_RF_U849 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3874
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n44
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3650);
   dp_id_stage_regfile_DataPath_Physical_RF_U848 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3874
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n45
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3649);
   dp_id_stage_regfile_DataPath_Physical_RF_U847 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3875
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n46
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3648);
   dp_id_stage_regfile_DataPath_Physical_RF_U846 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3875
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n47
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3647);
   dp_id_stage_regfile_DataPath_Physical_RF_U845 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3875
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n48
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3646);
   dp_id_stage_regfile_DataPath_Physical_RF_U844 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3875
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n49
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3645);
   dp_id_stage_regfile_DataPath_Physical_RF_U843 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3876
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n50
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3644);
   dp_id_stage_regfile_DataPath_Physical_RF_U842 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3876
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n51
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3643);
   dp_id_stage_regfile_DataPath_Physical_RF_U841 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3876
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n52
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3642);
   dp_id_stage_regfile_DataPath_Physical_RF_U840 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3876
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n53
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3641);
   dp_id_stage_regfile_DataPath_Physical_RF_U839 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3877
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n54
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3640);
   dp_id_stage_regfile_DataPath_Physical_RF_U838 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3877
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n55
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3639);
   dp_id_stage_regfile_DataPath_Physical_RF_U837 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3877
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n56
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3638);
   dp_id_stage_regfile_DataPath_Physical_RF_U836 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3877
                           , B2 => dp_id_stage_regfile_DataPath_Physical_RF_n57
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3637);
   dp_id_stage_regfile_DataPath_Physical_RF_U835 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3953
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n290, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3564);
   dp_id_stage_regfile_DataPath_Physical_RF_U834 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3953
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n291, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3563);
   dp_id_stage_regfile_DataPath_Physical_RF_U833 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3953
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n292, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3562);
   dp_id_stage_regfile_DataPath_Physical_RF_U832 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3953
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n293, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3561);
   dp_id_stage_regfile_DataPath_Physical_RF_U831 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3954
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n294, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3560);
   dp_id_stage_regfile_DataPath_Physical_RF_U830 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3954
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n295, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3559);
   dp_id_stage_regfile_DataPath_Physical_RF_U829 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3954
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n296, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3558);
   dp_id_stage_regfile_DataPath_Physical_RF_U828 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3954
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n297, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3557);
   dp_id_stage_regfile_DataPath_Physical_RF_U827 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3955
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n298, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3556);
   dp_id_stage_regfile_DataPath_Physical_RF_U826 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3955
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n299, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3555);
   dp_id_stage_regfile_DataPath_Physical_RF_U825 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3955
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n300, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3554);
   dp_id_stage_regfile_DataPath_Physical_RF_U824 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3955
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n301, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3553);
   dp_id_stage_regfile_DataPath_Physical_RF_U823 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3956
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n302, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3552);
   dp_id_stage_regfile_DataPath_Physical_RF_U822 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3956
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n303, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3551);
   dp_id_stage_regfile_DataPath_Physical_RF_U821 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3956
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n304, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3550);
   dp_id_stage_regfile_DataPath_Physical_RF_U820 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3956
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n305, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3549);
   dp_id_stage_regfile_DataPath_Physical_RF_U819 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3957
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n306, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3548);
   dp_id_stage_regfile_DataPath_Physical_RF_U818 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3957
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n307, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3547);
   dp_id_stage_regfile_DataPath_Physical_RF_U817 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3957
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n308, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3546);
   dp_id_stage_regfile_DataPath_Physical_RF_U816 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3957
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n309, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3545);
   dp_id_stage_regfile_DataPath_Physical_RF_U815 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3958
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n310, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3544);
   dp_id_stage_regfile_DataPath_Physical_RF_U814 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3958
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n311, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3543);
   dp_id_stage_regfile_DataPath_Physical_RF_U813 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3958
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n312, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3542);
   dp_id_stage_regfile_DataPath_Physical_RF_U812 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n3958
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n313, ZN =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3541);
   dp_id_stage_regfile_DataPath_Physical_RF_U811 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4189
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1026, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3212);
   dp_id_stage_regfile_DataPath_Physical_RF_U810 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4189
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1027, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3211);
   dp_id_stage_regfile_DataPath_Physical_RF_U809 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4189
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1028, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3210);
   dp_id_stage_regfile_DataPath_Physical_RF_U808 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4189
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1029, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3209);
   dp_id_stage_regfile_DataPath_Physical_RF_U807 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4265, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4190
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1030, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3208);
   dp_id_stage_regfile_DataPath_Physical_RF_U806 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4264, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4190
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1031, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3207);
   dp_id_stage_regfile_DataPath_Physical_RF_U805 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4190
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1032, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3206);
   dp_id_stage_regfile_DataPath_Physical_RF_U804 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4190
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1033, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3205);
   dp_id_stage_regfile_DataPath_Physical_RF_U803 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4191
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1034, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3204);
   dp_id_stage_regfile_DataPath_Physical_RF_U802 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4191
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1035, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3203);
   dp_id_stage_regfile_DataPath_Physical_RF_U801 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4191
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1036, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3202);
   dp_id_stage_regfile_DataPath_Physical_RF_U800 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4191
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1037, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3201);
   dp_id_stage_regfile_DataPath_Physical_RF_U799 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4192
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1038, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3200);
   dp_id_stage_regfile_DataPath_Physical_RF_U798 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4192
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1039, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3199);
   dp_id_stage_regfile_DataPath_Physical_RF_U797 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4192
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1040, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3198);
   dp_id_stage_regfile_DataPath_Physical_RF_U796 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4192
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1041, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3197);
   dp_id_stage_regfile_DataPath_Physical_RF_U795 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4193
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1042, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3196);
   dp_id_stage_regfile_DataPath_Physical_RF_U794 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4193
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1043, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3195);
   dp_id_stage_regfile_DataPath_Physical_RF_U793 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4193
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1044, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3194);
   dp_id_stage_regfile_DataPath_Physical_RF_U792 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4193
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1045, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3193);
   dp_id_stage_regfile_DataPath_Physical_RF_U791 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4194
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1046, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3192);
   dp_id_stage_regfile_DataPath_Physical_RF_U790 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4194
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1047, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3191);
   dp_id_stage_regfile_DataPath_Physical_RF_U789 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4194
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1048, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3190);
   dp_id_stage_regfile_DataPath_Physical_RF_U788 : OAI22_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188, 
                           B1 => dp_id_stage_regfile_DataPath_Physical_RF_n4194
                           , B2 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1049, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3189);
   dp_id_stage_regfile_DataPath_Physical_RF_U787 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_3_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1201);
   dp_id_stage_regfile_DataPath_Physical_RF_U786 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N429_port, 
                           Z => dp_id_stage_regfile_DataPath_Physical_RF_n4230)
                           ;
   dp_id_stage_regfile_DataPath_Physical_RF_U785 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N428_port, 
                           Z => dp_id_stage_regfile_DataPath_Physical_RF_n4233)
                           ;
   dp_id_stage_regfile_DataPath_Physical_RF_U784 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N429_port, 
                           Z => dp_id_stage_regfile_DataPath_Physical_RF_n4228)
                           ;
   dp_id_stage_regfile_DataPath_Physical_RF_U783 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N428_port, 
                           Z => dp_id_stage_regfile_DataPath_Physical_RF_n4231)
                           ;
   dp_id_stage_regfile_DataPath_Physical_RF_U782 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N429_port, 
                           Z => dp_id_stage_regfile_DataPath_Physical_RF_n4229)
                           ;
   dp_id_stage_regfile_DataPath_Physical_RF_U781 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N428_port, 
                           Z => dp_id_stage_regfile_DataPath_Physical_RF_n4232)
                           ;
   dp_id_stage_regfile_DataPath_Physical_RF_U780 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4234, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2536
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U779 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_0_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4270);
   dp_id_stage_regfile_DataPath_Physical_RF_U778 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_1_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4236);
   dp_id_stage_regfile_DataPath_Physical_RF_U777 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_0_port, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2529
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U776 : NOR3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_3_port, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_4_port, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n4235
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2548);
   dp_id_stage_regfile_DataPath_Physical_RF_U775 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_3_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1192);
   dp_id_stage_regfile_DataPath_Physical_RF_U774 : AND4_X2 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_3_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1342, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1191
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1190, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1686);
   dp_id_stage_regfile_DataPath_Physical_RF_U773 : AND4_X2 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_4_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1342, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1192
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1190, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1517);
   dp_id_stage_regfile_DataPath_Physical_RF_U772 : AND4_X2 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1342, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1192, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1191
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1190, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1823);
   dp_id_stage_regfile_DataPath_Physical_RF_U771 : AND4_X2 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_4_port, A2 
                           => dp_id_stage_regfile_DataPath_mux_wr_out_3_port, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1342
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1190, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1345);
   dp_id_stage_regfile_DataPath_Physical_RF_U770 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_4_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4234);
   dp_id_stage_regfile_DataPath_Physical_RF_U769 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_4_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1195);
   dp_id_stage_regfile_DataPath_Physical_RF_U768 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_3_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1196);
   dp_id_stage_regfile_DataPath_Physical_RF_U767 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_2_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1197);
   dp_id_stage_regfile_DataPath_Physical_RF_U766 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2531, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1980
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U765 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2551, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1973
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U764 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2549, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1968
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U763 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2539, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1947
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U762 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2535, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1941
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U761 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2528, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1937
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U760 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_5_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1953
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U759 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_5_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2580
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U758 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2531, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1979
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U757 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2535, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1943
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U756 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2535, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1942
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U755 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2528, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1936
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U754 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2532, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1954
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U753 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2530, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1952
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U752 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3159, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2581
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U751 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3157, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2579
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U750 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2548, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1969
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U749 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2548, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1967
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U748 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2546, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1963
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U747 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2546, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1962
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U746 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2551, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1976
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U745 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2549, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1971
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U744 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2539, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1945
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U743 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2551, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1975
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U742 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2549, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1970
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U741 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2539, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1944
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U740 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2528, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1939
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U739 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2531, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2532, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1934
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U738 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2536, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4235, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2531
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U737 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3179, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3178
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U736 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3163, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3155
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U735 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2536, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2528
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U734 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1195, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_3_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3163
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U733 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1196, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3179
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U732 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2529, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1949
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U731 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3156, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_5_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2576
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U730 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1201, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_4_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2552
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U729 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4234, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1201, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2538
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U728 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_2_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3165, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3166
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U727 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_0_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1199);
   dp_id_stage_regfile_DataPath_Physical_RF_U726 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_1_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1198);
   dp_id_stage_regfile_DataPath_Physical_RF_U725 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2548, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1964
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U724 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2548, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1965
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U723 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2546, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2530, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1959
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U722 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2546, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2529, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1960
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U721 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_0_port, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3156
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U720 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4236, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4270, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2533
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U719 : NOR3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_3_port, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_4_port, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1197
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3175);
   dp_id_stage_regfile_DataPath_Physical_RF_U718 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_0_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1194);
   dp_id_stage_regfile_DataPath_Physical_RF_U717 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_4_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1191);
   dp_id_stage_regfile_DataPath_Physical_RF_U716 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_1_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1193);
   dp_id_stage_regfile_DataPath_Physical_RF_U715 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1686, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1344, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1654
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U714 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1686, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1383, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1690
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U713 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1823, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1347, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1825
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U712 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1823, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1344, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1791
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U711 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1517, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1383, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1553
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U710 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1517, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1349, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1520
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U709 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1383, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1345, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1351
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U708 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_5_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1190);
   dp_id_stage_regfile_DataPath_Physical_RF_U707 : AND3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_1_port, A2 
                           => dp_id_stage_regfile_DataPath_mux_wr_out_0_port, 
                           A3 => dp_id_stage_regfile_DataPath_mux_wr_out_2_port
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1344);
   dp_id_stage_regfile_DataPath_Physical_RF_U706 : AND3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1194, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1193, 
                           A3 => dp_id_stage_regfile_DataPath_mux_wr_out_2_port
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1383);
   dp_id_stage_regfile_DataPath_Physical_RF_U705 : AND3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_1_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1194, 
                           A3 => dp_id_stage_regfile_DataPath_mux_wr_out_2_port
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1347);
   dp_id_stage_regfile_DataPath_Physical_RF_U704 : AND3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_0_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1193, 
                           A3 => dp_id_stage_regfile_DataPath_mux_wr_out_2_port
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1349);
   dp_id_stage_regfile_DataPath_Physical_RF_U703 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1686, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1341, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1758
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U702 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1517, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1341, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1621
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U701 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1345, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1341, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1484
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U700 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1823, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1305, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1893
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U699 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1823, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1270, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1860
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U698 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1686, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1270, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1723
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U697 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1345, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1305, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1418
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U696 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1345, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1270, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1385
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U695 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1517, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1339, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1588
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U694 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1345, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1339, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1451
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U693 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1270, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1271, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1238
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U692 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1305, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1271, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1273
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U691 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1339, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1271, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1307
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U690 : INV_X1 port map( A => dp_n12
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4269);
   dp_id_stage_regfile_DataPath_Physical_RF_U689 : INV_X1 port map( A => dp_n10
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4268);
   dp_id_stage_regfile_DataPath_Physical_RF_U688 : INV_X1 port map( A => 
                           dp_wr_data_id_i_29_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4267);
   dp_id_stage_regfile_DataPath_Physical_RF_U687 : INV_X1 port map( A => 
                           dp_wr_data_id_i_28_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4266);
   dp_id_stage_regfile_DataPath_Physical_RF_U686 : INV_X1 port map( A => dp_n8,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n4265
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U685 : INV_X1 port map( A => dp_n6,
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n4264
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U684 : INV_X1 port map( A => 
                           dp_wr_data_id_i_25_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4263);
   dp_id_stage_regfile_DataPath_Physical_RF_U683 : INV_X1 port map( A => 
                           dp_wr_data_id_i_24_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4262);
   dp_id_stage_regfile_DataPath_Physical_RF_U682 : INV_X1 port map( A => 
                           dp_wr_data_id_i_23_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4261);
   dp_id_stage_regfile_DataPath_Physical_RF_U681 : INV_X1 port map( A => 
                           dp_wr_data_id_i_22_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4260);
   dp_id_stage_regfile_DataPath_Physical_RF_U680 : INV_X1 port map( A => 
                           dp_wr_data_id_i_21_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4259);
   dp_id_stage_regfile_DataPath_Physical_RF_U679 : INV_X1 port map( A => 
                           dp_wr_data_id_i_20_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4258);
   dp_id_stage_regfile_DataPath_Physical_RF_U678 : INV_X1 port map( A => 
                           dp_wr_data_id_i_19_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4257);
   dp_id_stage_regfile_DataPath_Physical_RF_U677 : INV_X1 port map( A => 
                           dp_wr_data_id_i_18_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4256);
   dp_id_stage_regfile_DataPath_Physical_RF_U676 : INV_X1 port map( A => 
                           dp_wr_data_id_i_17_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4255);
   dp_id_stage_regfile_DataPath_Physical_RF_U675 : INV_X1 port map( A => 
                           dp_wr_data_id_i_16_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4254);
   dp_id_stage_regfile_DataPath_Physical_RF_U674 : INV_X1 port map( A => 
                           dp_wr_data_id_i_15_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4253);
   dp_id_stage_regfile_DataPath_Physical_RF_U673 : INV_X1 port map( A => 
                           dp_wr_data_id_i_14_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4252);
   dp_id_stage_regfile_DataPath_Physical_RF_U672 : INV_X1 port map( A => 
                           dp_wr_data_id_i_13_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4251);
   dp_id_stage_regfile_DataPath_Physical_RF_U671 : INV_X1 port map( A => 
                           dp_wr_data_id_i_12_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4250);
   dp_id_stage_regfile_DataPath_Physical_RF_U670 : INV_X1 port map( A => 
                           dp_wr_data_id_i_11_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4249);
   dp_id_stage_regfile_DataPath_Physical_RF_U669 : INV_X1 port map( A => 
                           dp_wr_data_id_i_10_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4248);
   dp_id_stage_regfile_DataPath_Physical_RF_U668 : INV_X1 port map( A => 
                           dp_wr_data_id_i_9_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4247);
   dp_id_stage_regfile_DataPath_Physical_RF_U667 : INV_X1 port map( A => 
                           dp_wr_data_id_i_8_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4246);
   dp_id_stage_regfile_DataPath_Physical_RF_U666 : INV_X1 port map( A => 
                           dp_wr_data_id_i_7_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4245);
   dp_id_stage_regfile_DataPath_Physical_RF_U665 : INV_X1 port map( A => 
                           dp_wr_data_id_i_6_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4244);
   dp_id_stage_regfile_DataPath_Physical_RF_U664 : INV_X1 port map( A => 
                           dp_wr_data_id_i_5_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4243);
   dp_id_stage_regfile_DataPath_Physical_RF_U663 : INV_X1 port map( A => 
                           dp_wr_data_id_i_4_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4242);
   dp_id_stage_regfile_DataPath_Physical_RF_U662 : INV_X1 port map( A => 
                           dp_wr_data_id_i_3_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4241);
   dp_id_stage_regfile_DataPath_Physical_RF_U661 : INV_X1 port map( A => 
                           dp_wr_data_id_i_2_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4240);
   dp_id_stage_regfile_DataPath_Physical_RF_U660 : INV_X1 port map( A => 
                           dp_wr_data_id_i_1_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4239);
   dp_id_stage_regfile_DataPath_Physical_RF_U659 : INV_X1 port map( A => 
                           dp_wr_data_id_i_0_port, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4238);
   dp_id_stage_regfile_DataPath_Physical_RF_U658 : NOR3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1194, A2 
                           => dp_id_stage_regfile_DataPath_mux_wr_out_2_port, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1193
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1270);
   dp_id_stage_regfile_DataPath_Physical_RF_U657 : NOR3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_1_port, A2 
                           => dp_id_stage_regfile_DataPath_mux_wr_out_2_port, 
                           A3 => dp_id_stage_regfile_DataPath_mux_wr_out_0_port
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1341);
   dp_id_stage_regfile_DataPath_Physical_RF_U656 : NOR3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_0_port, A2 
                           => dp_id_stage_regfile_DataPath_mux_wr_out_2_port, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1193
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1305);
   dp_id_stage_regfile_DataPath_Physical_RF_U655 : NOR3_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_1_port, A2 
                           => dp_id_stage_regfile_DataPath_mux_wr_out_2_port, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1194
                           , ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1339);
   dp_id_stage_regfile_DataPath_Physical_RF_U654 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1173);
   dp_id_stage_regfile_DataPath_Physical_RF_U653 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1172);
   dp_id_stage_regfile_DataPath_Physical_RF_U652 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2538, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4235, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2535
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U651 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3165, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1197, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3162
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U650 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_2_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4235);
   dp_id_stage_regfile_DataPath_Physical_RF_U649 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3158, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2607
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U648 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3178, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2600
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U647 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3176, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2595
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U646 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3166, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2574
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U645 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3162, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2568
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U644 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3155, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2564
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U643 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2551, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1978
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U642 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2549, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1974
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U641 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2535, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1948
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U640 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3178, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2605
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U639 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3158, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2606
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U638 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3162, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2570
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U637 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3162, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2569
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U636 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3155, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2563
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U635 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3175, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2596
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U634 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3175, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2594
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U633 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3173, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2590
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U632 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3173, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2589
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U631 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2539, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1950
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U630 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2528, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1938
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U629 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2531, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2533, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1933
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U628 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3166, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2577
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U627 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3155, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2565
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U626 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3178, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2603
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U625 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3176, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2598
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U624 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3166, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2572
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U623 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3178, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2602
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U622 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3176, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2597
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U621 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3166, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2571
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U620 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3155, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2566
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U619 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3158, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3159, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2561
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U618 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2552, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4235, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2549
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U617 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3179, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1197, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3176
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U616 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3163, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1197, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3158
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U615 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2552, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_2_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2551
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U614 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1195, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1196, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3165
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U613 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_2_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2538, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2539
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U612 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3175, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2591
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U611 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3175, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2592
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U610 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1980, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3753);
   dp_id_stage_regfile_DataPath_Physical_RF_U609 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1969, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3780);
   dp_id_stage_regfile_DataPath_Physical_RF_U608 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1954, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3807);
   dp_id_stage_regfile_DataPath_Physical_RF_U607 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1943, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3834);
   dp_id_stage_regfile_DataPath_Physical_RF_U606 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2581, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3699);
   dp_id_stage_regfile_DataPath_Physical_RF_U605 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1937, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3849);
   dp_id_stage_regfile_DataPath_Physical_RF_U604 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1963, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3795);
   dp_id_stage_regfile_DataPath_Physical_RF_U603 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1979, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3756);
   dp_id_stage_regfile_DataPath_Physical_RF_U602 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1968, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3783);
   dp_id_stage_regfile_DataPath_Physical_RF_U601 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1953, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3810);
   dp_id_stage_regfile_DataPath_Physical_RF_U600 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1942, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3837);
   dp_id_stage_regfile_DataPath_Physical_RF_U599 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2580, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3702);
   dp_id_stage_regfile_DataPath_Physical_RF_U598 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1975, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3765);
   dp_id_stage_regfile_DataPath_Physical_RF_U597 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1970, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3777);
   dp_id_stage_regfile_DataPath_Physical_RF_U596 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1964, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3792);
   dp_id_stage_regfile_DataPath_Physical_RF_U595 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1959, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3804);
   dp_id_stage_regfile_DataPath_Physical_RF_U594 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1949, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3819);
   dp_id_stage_regfile_DataPath_Physical_RF_U593 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1944, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3831);
   dp_id_stage_regfile_DataPath_Physical_RF_U592 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2576, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3711);
   dp_id_stage_regfile_DataPath_Physical_RF_U591 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1973, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3771);
   dp_id_stage_regfile_DataPath_Physical_RF_U590 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1947, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3825);
   dp_id_stage_regfile_DataPath_Physical_RF_U589 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1936, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3852);
   dp_id_stage_regfile_DataPath_Physical_RF_U588 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1962, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3798);
   dp_id_stage_regfile_DataPath_Physical_RF_U587 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1967, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3786);
   dp_id_stage_regfile_DataPath_Physical_RF_U586 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1952, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3813);
   dp_id_stage_regfile_DataPath_Physical_RF_U585 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1941, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3840);
   dp_id_stage_regfile_DataPath_Physical_RF_U584 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2579, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3705);
   dp_id_stage_regfile_DataPath_Physical_RF_U583 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3173, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3157, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2586
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U582 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3173, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3156, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2587
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U581 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1976, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3762);
   dp_id_stage_regfile_DataPath_Physical_RF_U580 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1971, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3774);
   dp_id_stage_regfile_DataPath_Physical_RF_U579 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1965, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3789);
   dp_id_stage_regfile_DataPath_Physical_RF_U578 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1960, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3801);
   dp_id_stage_regfile_DataPath_Physical_RF_U577 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1945, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3828);
   dp_id_stage_regfile_DataPath_Physical_RF_U576 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1939, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3843);
   dp_id_stage_regfile_DataPath_Physical_RF_U575 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1934, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3855);
   dp_id_stage_regfile_DataPath_Physical_RF_U574 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1980, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3752);
   dp_id_stage_regfile_DataPath_Physical_RF_U573 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1969, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3779);
   dp_id_stage_regfile_DataPath_Physical_RF_U572 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1954, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3806);
   dp_id_stage_regfile_DataPath_Physical_RF_U571 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1943, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3833);
   dp_id_stage_regfile_DataPath_Physical_RF_U570 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2581, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3698);
   dp_id_stage_regfile_DataPath_Physical_RF_U569 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1980, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3751);
   dp_id_stage_regfile_DataPath_Physical_RF_U568 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1969, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3778);
   dp_id_stage_regfile_DataPath_Physical_RF_U567 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1954, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3805);
   dp_id_stage_regfile_DataPath_Physical_RF_U566 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1943, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3832);
   dp_id_stage_regfile_DataPath_Physical_RF_U565 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2581, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3697);
   dp_id_stage_regfile_DataPath_Physical_RF_U564 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1963, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3794);
   dp_id_stage_regfile_DataPath_Physical_RF_U563 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1937, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3848);
   dp_id_stage_regfile_DataPath_Physical_RF_U562 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1963, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3793);
   dp_id_stage_regfile_DataPath_Physical_RF_U561 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1937, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3847);
   dp_id_stage_regfile_DataPath_Physical_RF_U560 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1979, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3755);
   dp_id_stage_regfile_DataPath_Physical_RF_U559 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1968, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3782);
   dp_id_stage_regfile_DataPath_Physical_RF_U558 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1953, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3809);
   dp_id_stage_regfile_DataPath_Physical_RF_U557 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1942, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3836);
   dp_id_stage_regfile_DataPath_Physical_RF_U556 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2580, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3701);
   dp_id_stage_regfile_DataPath_Physical_RF_U555 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1979, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3754);
   dp_id_stage_regfile_DataPath_Physical_RF_U554 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1968, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3781);
   dp_id_stage_regfile_DataPath_Physical_RF_U553 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1953, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3808);
   dp_id_stage_regfile_DataPath_Physical_RF_U552 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1942, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3835);
   dp_id_stage_regfile_DataPath_Physical_RF_U551 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2580, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3700);
   dp_id_stage_regfile_DataPath_Physical_RF_U550 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1975, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3763);
   dp_id_stage_regfile_DataPath_Physical_RF_U549 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1970, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3775);
   dp_id_stage_regfile_DataPath_Physical_RF_U548 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1964, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3790);
   dp_id_stage_regfile_DataPath_Physical_RF_U547 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1959, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3802);
   dp_id_stage_regfile_DataPath_Physical_RF_U546 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1949, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3817);
   dp_id_stage_regfile_DataPath_Physical_RF_U545 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1944, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3829);
   dp_id_stage_regfile_DataPath_Physical_RF_U544 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2576, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3709);
   dp_id_stage_regfile_DataPath_Physical_RF_U543 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1975, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3764);
   dp_id_stage_regfile_DataPath_Physical_RF_U542 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1970, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3776);
   dp_id_stage_regfile_DataPath_Physical_RF_U541 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1964, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3791);
   dp_id_stage_regfile_DataPath_Physical_RF_U540 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1959, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3803);
   dp_id_stage_regfile_DataPath_Physical_RF_U539 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1949, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3818);
   dp_id_stage_regfile_DataPath_Physical_RF_U538 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1944, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3830);
   dp_id_stage_regfile_DataPath_Physical_RF_U537 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2576, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3710);
   dp_id_stage_regfile_DataPath_Physical_RF_U536 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1973, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3769);
   dp_id_stage_regfile_DataPath_Physical_RF_U535 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1962, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3796);
   dp_id_stage_regfile_DataPath_Physical_RF_U534 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1947, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3823);
   dp_id_stage_regfile_DataPath_Physical_RF_U533 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1936, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3850);
   dp_id_stage_regfile_DataPath_Physical_RF_U532 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1973, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3770);
   dp_id_stage_regfile_DataPath_Physical_RF_U531 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1962, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3797);
   dp_id_stage_regfile_DataPath_Physical_RF_U530 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1947, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3824);
   dp_id_stage_regfile_DataPath_Physical_RF_U529 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1936, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3851);
   dp_id_stage_regfile_DataPath_Physical_RF_U528 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1967, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3784);
   dp_id_stage_regfile_DataPath_Physical_RF_U527 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1952, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3811);
   dp_id_stage_regfile_DataPath_Physical_RF_U526 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1941, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3838);
   dp_id_stage_regfile_DataPath_Physical_RF_U525 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2579, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3703);
   dp_id_stage_regfile_DataPath_Physical_RF_U524 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1967, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3785);
   dp_id_stage_regfile_DataPath_Physical_RF_U523 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1952, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3812);
   dp_id_stage_regfile_DataPath_Physical_RF_U522 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1941, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3839);
   dp_id_stage_regfile_DataPath_Physical_RF_U521 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2579, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3704);
   dp_id_stage_regfile_DataPath_Physical_RF_U520 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1976, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3760);
   dp_id_stage_regfile_DataPath_Physical_RF_U519 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1971, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3772);
   dp_id_stage_regfile_DataPath_Physical_RF_U518 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1965, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3787);
   dp_id_stage_regfile_DataPath_Physical_RF_U517 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1960, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3799);
   dp_id_stage_regfile_DataPath_Physical_RF_U516 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1945, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3826);
   dp_id_stage_regfile_DataPath_Physical_RF_U515 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1939, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3841);
   dp_id_stage_regfile_DataPath_Physical_RF_U514 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1934, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3853);
   dp_id_stage_regfile_DataPath_Physical_RF_U513 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1976, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3761);
   dp_id_stage_regfile_DataPath_Physical_RF_U512 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1971, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3773);
   dp_id_stage_regfile_DataPath_Physical_RF_U511 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1965, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3788);
   dp_id_stage_regfile_DataPath_Physical_RF_U510 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1960, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3800);
   dp_id_stage_regfile_DataPath_Physical_RF_U509 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1945, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3827);
   dp_id_stage_regfile_DataPath_Physical_RF_U508 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1939, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3842);
   dp_id_stage_regfile_DataPath_Physical_RF_U507 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1934, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3854);
   dp_id_stage_regfile_DataPath_Physical_RF_U506 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1198, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1199, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3160
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U505 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1654, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4022);
   dp_id_stage_regfile_DataPath_Physical_RF_U504 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1690, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3991);
   dp_id_stage_regfile_DataPath_Physical_RF_U503 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1825, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3931);
   dp_id_stage_regfile_DataPath_Physical_RF_U502 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1791, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3940);
   dp_id_stage_regfile_DataPath_Physical_RF_U501 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1553, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4073);
   dp_id_stage_regfile_DataPath_Physical_RF_U500 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1520, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4082);
   dp_id_stage_regfile_DataPath_Physical_RF_U499 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1238, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4227);
   dp_id_stage_regfile_DataPath_Physical_RF_U498 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1273, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4217);
   dp_id_stage_regfile_DataPath_Physical_RF_U497 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1307, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4207);
   dp_id_stage_regfile_DataPath_Physical_RF_U496 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1351, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4153);
   dp_id_stage_regfile_DataPath_Physical_RF_U495 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1758, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3950);
   dp_id_stage_regfile_DataPath_Physical_RF_U494 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1621, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4032);
   dp_id_stage_regfile_DataPath_Physical_RF_U493 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1484, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4114);
   dp_id_stage_regfile_DataPath_Physical_RF_U492 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1893, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3890);
   dp_id_stage_regfile_DataPath_Physical_RF_U491 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1860, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3900);
   dp_id_stage_regfile_DataPath_Physical_RF_U490 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1723, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3982);
   dp_id_stage_regfile_DataPath_Physical_RF_U489 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1418, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4134);
   dp_id_stage_regfile_DataPath_Physical_RF_U488 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1385, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4144);
   dp_id_stage_regfile_DataPath_Physical_RF_U487 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1588, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4042);
   dp_id_stage_regfile_DataPath_Physical_RF_U486 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1451, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4124);
   dp_id_stage_regfile_DataPath_Physical_RF_U485 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1654, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4021);
   dp_id_stage_regfile_DataPath_Physical_RF_U484 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1654, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4020);
   dp_id_stage_regfile_DataPath_Physical_RF_U483 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1654, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4019);
   dp_id_stage_regfile_DataPath_Physical_RF_U482 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1654, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4018);
   dp_id_stage_regfile_DataPath_Physical_RF_U481 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1654, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4017);
   dp_id_stage_regfile_DataPath_Physical_RF_U480 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1654, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4016);
   dp_id_stage_regfile_DataPath_Physical_RF_U479 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1351, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4152);
   dp_id_stage_regfile_DataPath_Physical_RF_U478 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1351, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4151);
   dp_id_stage_regfile_DataPath_Physical_RF_U477 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1351, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4150);
   dp_id_stage_regfile_DataPath_Physical_RF_U476 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1351, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4149);
   dp_id_stage_regfile_DataPath_Physical_RF_U475 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1351, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4148);
   dp_id_stage_regfile_DataPath_Physical_RF_U474 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1351, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4147);
   dp_id_stage_regfile_DataPath_Physical_RF_U473 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1690, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3990);
   dp_id_stage_regfile_DataPath_Physical_RF_U472 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1690, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3989);
   dp_id_stage_regfile_DataPath_Physical_RF_U471 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1690, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3988);
   dp_id_stage_regfile_DataPath_Physical_RF_U470 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1690, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3987);
   dp_id_stage_regfile_DataPath_Physical_RF_U469 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1690, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3986);
   dp_id_stage_regfile_DataPath_Physical_RF_U468 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1690, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3985);
   dp_id_stage_regfile_DataPath_Physical_RF_U467 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1173, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1169);
   dp_id_stage_regfile_DataPath_Physical_RF_U466 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1172, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1170);
   dp_id_stage_regfile_DataPath_Physical_RF_U465 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1172, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1171);
   dp_id_stage_regfile_DataPath_Physical_RF_U464 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3176, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2601
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U463 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3162, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2575
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U462 : NAND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3158, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3160, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2560
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U461 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2607, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1205);
   dp_id_stage_regfile_DataPath_Physical_RF_U460 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2596, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1232);
   dp_id_stage_regfile_DataPath_Physical_RF_U459 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2570, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3726);
   dp_id_stage_regfile_DataPath_Physical_RF_U458 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1974, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3768);
   dp_id_stage_regfile_DataPath_Physical_RF_U457 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1948, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3822);
   dp_id_stage_regfile_DataPath_Physical_RF_U456 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2564, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3741);
   dp_id_stage_regfile_DataPath_Physical_RF_U455 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2590, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1755);
   dp_id_stage_regfile_DataPath_Physical_RF_U454 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2606, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1208);
   dp_id_stage_regfile_DataPath_Physical_RF_U453 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2595, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1235);
   dp_id_stage_regfile_DataPath_Physical_RF_U452 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2569, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3729);
   dp_id_stage_regfile_DataPath_Physical_RF_U451 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1938, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3846);
   dp_id_stage_regfile_DataPath_Physical_RF_U450 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1933, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3858);
   dp_id_stage_regfile_DataPath_Physical_RF_U449 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2602, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1217);
   dp_id_stage_regfile_DataPath_Physical_RF_U448 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2597, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1229);
   dp_id_stage_regfile_DataPath_Physical_RF_U447 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2591, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1586);
   dp_id_stage_regfile_DataPath_Physical_RF_U446 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2586, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3696);
   dp_id_stage_regfile_DataPath_Physical_RF_U445 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2571, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3723);
   dp_id_stage_regfile_DataPath_Physical_RF_U444 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2565, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3738);
   dp_id_stage_regfile_DataPath_Physical_RF_U443 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2600, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1223);
   dp_id_stage_regfile_DataPath_Physical_RF_U442 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2574, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3717);
   dp_id_stage_regfile_DataPath_Physical_RF_U441 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2563, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3744);
   dp_id_stage_regfile_DataPath_Physical_RF_U440 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2589, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1858);
   dp_id_stage_regfile_DataPath_Physical_RF_U439 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1978, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3759);
   dp_id_stage_regfile_DataPath_Physical_RF_U438 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2605, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1211);
   dp_id_stage_regfile_DataPath_Physical_RF_U437 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2594, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1343);
   dp_id_stage_regfile_DataPath_Physical_RF_U436 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2568, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3732);
   dp_id_stage_regfile_DataPath_Physical_RF_U435 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1950, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3816);
   dp_id_stage_regfile_DataPath_Physical_RF_U434 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2603, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1214);
   dp_id_stage_regfile_DataPath_Physical_RF_U433 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2598, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1226);
   dp_id_stage_regfile_DataPath_Physical_RF_U432 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2592, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1516);
   dp_id_stage_regfile_DataPath_Physical_RF_U431 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2587, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3693);
   dp_id_stage_regfile_DataPath_Physical_RF_U430 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2577, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3708);
   dp_id_stage_regfile_DataPath_Physical_RF_U429 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2572, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3720);
   dp_id_stage_regfile_DataPath_Physical_RF_U428 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2566, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3735);
   dp_id_stage_regfile_DataPath_Physical_RF_U427 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2561, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3747);
   dp_id_stage_regfile_DataPath_Physical_RF_U426 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2607, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1204);
   dp_id_stage_regfile_DataPath_Physical_RF_U425 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2596, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1231);
   dp_id_stage_regfile_DataPath_Physical_RF_U424 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2570, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3725);
   dp_id_stage_regfile_DataPath_Physical_RF_U423 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2607, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1203);
   dp_id_stage_regfile_DataPath_Physical_RF_U422 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2596, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1230);
   dp_id_stage_regfile_DataPath_Physical_RF_U421 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2570, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3724);
   dp_id_stage_regfile_DataPath_Physical_RF_U420 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1974, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3767);
   dp_id_stage_regfile_DataPath_Physical_RF_U419 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1948, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3821);
   dp_id_stage_regfile_DataPath_Physical_RF_U418 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2590, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1688);
   dp_id_stage_regfile_DataPath_Physical_RF_U417 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2564, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3740);
   dp_id_stage_regfile_DataPath_Physical_RF_U416 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1974, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3766);
   dp_id_stage_regfile_DataPath_Physical_RF_U415 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1948, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3820);
   dp_id_stage_regfile_DataPath_Physical_RF_U414 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2590, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1687);
   dp_id_stage_regfile_DataPath_Physical_RF_U413 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2564, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3739);
   dp_id_stage_regfile_DataPath_Physical_RF_U412 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2606, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1207);
   dp_id_stage_regfile_DataPath_Physical_RF_U411 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2595, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1234);
   dp_id_stage_regfile_DataPath_Physical_RF_U410 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2569, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3728);
   dp_id_stage_regfile_DataPath_Physical_RF_U409 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2606, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1206);
   dp_id_stage_regfile_DataPath_Physical_RF_U408 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2595, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1233);
   dp_id_stage_regfile_DataPath_Physical_RF_U407 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2569, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3727);
   dp_id_stage_regfile_DataPath_Physical_RF_U406 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1938, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3844);
   dp_id_stage_regfile_DataPath_Physical_RF_U405 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1933, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3856);
   dp_id_stage_regfile_DataPath_Physical_RF_U404 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2602, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1215);
   dp_id_stage_regfile_DataPath_Physical_RF_U403 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2597, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1227);
   dp_id_stage_regfile_DataPath_Physical_RF_U402 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2591, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1518);
   dp_id_stage_regfile_DataPath_Physical_RF_U401 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2586, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3694);
   dp_id_stage_regfile_DataPath_Physical_RF_U400 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2571, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3721);
   dp_id_stage_regfile_DataPath_Physical_RF_U399 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2565, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3736);
   dp_id_stage_regfile_DataPath_Physical_RF_U398 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1938, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3845);
   dp_id_stage_regfile_DataPath_Physical_RF_U397 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1933, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3857);
   dp_id_stage_regfile_DataPath_Physical_RF_U396 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2602, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1216);
   dp_id_stage_regfile_DataPath_Physical_RF_U395 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2597, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1228);
   dp_id_stage_regfile_DataPath_Physical_RF_U394 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2591, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1585);
   dp_id_stage_regfile_DataPath_Physical_RF_U393 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2586, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3695);
   dp_id_stage_regfile_DataPath_Physical_RF_U392 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2571, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3722);
   dp_id_stage_regfile_DataPath_Physical_RF_U391 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2565, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3737);
   dp_id_stage_regfile_DataPath_Physical_RF_U390 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2600, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1221);
   dp_id_stage_regfile_DataPath_Physical_RF_U389 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2589, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1756);
   dp_id_stage_regfile_DataPath_Physical_RF_U388 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2574, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3715);
   dp_id_stage_regfile_DataPath_Physical_RF_U387 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2563, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3742);
   dp_id_stage_regfile_DataPath_Physical_RF_U386 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2600, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1222);
   dp_id_stage_regfile_DataPath_Physical_RF_U385 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2589, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1857);
   dp_id_stage_regfile_DataPath_Physical_RF_U384 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2574, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3716);
   dp_id_stage_regfile_DataPath_Physical_RF_U383 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2563, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3743);
   dp_id_stage_regfile_DataPath_Physical_RF_U382 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1978, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3757);
   dp_id_stage_regfile_DataPath_Physical_RF_U381 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2605, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1209);
   dp_id_stage_regfile_DataPath_Physical_RF_U380 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2594, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1236);
   dp_id_stage_regfile_DataPath_Physical_RF_U379 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2568, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3730);
   dp_id_stage_regfile_DataPath_Physical_RF_U378 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1978, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3758);
   dp_id_stage_regfile_DataPath_Physical_RF_U377 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2605, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1210);
   dp_id_stage_regfile_DataPath_Physical_RF_U376 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2594, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1340);
   dp_id_stage_regfile_DataPath_Physical_RF_U375 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2568, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3731);
   dp_id_stage_regfile_DataPath_Physical_RF_U374 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1950, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3814);
   dp_id_stage_regfile_DataPath_Physical_RF_U373 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2603, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1212);
   dp_id_stage_regfile_DataPath_Physical_RF_U372 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2598, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1224);
   dp_id_stage_regfile_DataPath_Physical_RF_U371 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2592, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1346);
   dp_id_stage_regfile_DataPath_Physical_RF_U370 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2587, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1925);
   dp_id_stage_regfile_DataPath_Physical_RF_U369 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2577, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3706);
   dp_id_stage_regfile_DataPath_Physical_RF_U368 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2572, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3718);
   dp_id_stage_regfile_DataPath_Physical_RF_U367 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2566, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3733);
   dp_id_stage_regfile_DataPath_Physical_RF_U366 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2561, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3745);
   dp_id_stage_regfile_DataPath_Physical_RF_U365 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1950, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3815);
   dp_id_stage_regfile_DataPath_Physical_RF_U364 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2603, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1213);
   dp_id_stage_regfile_DataPath_Physical_RF_U363 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2598, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1225);
   dp_id_stage_regfile_DataPath_Physical_RF_U362 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2592, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1348);
   dp_id_stage_regfile_DataPath_Physical_RF_U361 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2587, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1926);
   dp_id_stage_regfile_DataPath_Physical_RF_U360 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2577, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3707);
   dp_id_stage_regfile_DataPath_Physical_RF_U359 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2572, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3719);
   dp_id_stage_regfile_DataPath_Physical_RF_U358 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2566, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3734);
   dp_id_stage_regfile_DataPath_Physical_RF_U357 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2561, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3746);
   dp_id_stage_regfile_DataPath_Physical_RF_U356 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1161, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4178);
   dp_id_stage_regfile_DataPath_Physical_RF_U355 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1161, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4179);
   dp_id_stage_regfile_DataPath_Physical_RF_U354 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1161, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4180);
   dp_id_stage_regfile_DataPath_Physical_RF_U353 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1161, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4181);
   dp_id_stage_regfile_DataPath_Physical_RF_U352 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1161, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4182);
   dp_id_stage_regfile_DataPath_Physical_RF_U351 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1161, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4183);
   dp_id_stage_regfile_DataPath_Physical_RF_U350 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4178, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4184);
   dp_id_stage_regfile_DataPath_Physical_RF_U349 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4179, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4185);
   dp_id_stage_regfile_DataPath_Physical_RF_U348 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1160, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4167);
   dp_id_stage_regfile_DataPath_Physical_RF_U347 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1160, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4168);
   dp_id_stage_regfile_DataPath_Physical_RF_U346 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1160, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4169);
   dp_id_stage_regfile_DataPath_Physical_RF_U345 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1160, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4170);
   dp_id_stage_regfile_DataPath_Physical_RF_U344 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1160, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4171);
   dp_id_stage_regfile_DataPath_Physical_RF_U343 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1160, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4172);
   dp_id_stage_regfile_DataPath_Physical_RF_U342 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1159, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4156);
   dp_id_stage_regfile_DataPath_Physical_RF_U341 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1159, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4157);
   dp_id_stage_regfile_DataPath_Physical_RF_U340 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1159, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4158);
   dp_id_stage_regfile_DataPath_Physical_RF_U339 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1159, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4159);
   dp_id_stage_regfile_DataPath_Physical_RF_U338 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1159, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4160);
   dp_id_stage_regfile_DataPath_Physical_RF_U337 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1159, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4161);
   dp_id_stage_regfile_DataPath_Physical_RF_U336 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4167, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4173);
   dp_id_stage_regfile_DataPath_Physical_RF_U335 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4168, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4174);
   dp_id_stage_regfile_DataPath_Physical_RF_U334 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4156, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4162);
   dp_id_stage_regfile_DataPath_Physical_RF_U333 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4157, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4163);
   dp_id_stage_regfile_DataPath_Physical_RF_U332 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1158, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4005);
   dp_id_stage_regfile_DataPath_Physical_RF_U331 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1158, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4006);
   dp_id_stage_regfile_DataPath_Physical_RF_U330 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1158, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4007);
   dp_id_stage_regfile_DataPath_Physical_RF_U329 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1158, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4008);
   dp_id_stage_regfile_DataPath_Physical_RF_U328 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1158, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4009);
   dp_id_stage_regfile_DataPath_Physical_RF_U327 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1158, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4010);
   dp_id_stage_regfile_DataPath_Physical_RF_U326 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1157, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3994);
   dp_id_stage_regfile_DataPath_Physical_RF_U325 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1157, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3995);
   dp_id_stage_regfile_DataPath_Physical_RF_U324 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1157, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3996);
   dp_id_stage_regfile_DataPath_Physical_RF_U323 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1157, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3997);
   dp_id_stage_regfile_DataPath_Physical_RF_U322 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1157, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3998);
   dp_id_stage_regfile_DataPath_Physical_RF_U321 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1157, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3999);
   dp_id_stage_regfile_DataPath_Physical_RF_U320 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4005, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4011);
   dp_id_stage_regfile_DataPath_Physical_RF_U319 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4006, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4012);
   dp_id_stage_regfile_DataPath_Physical_RF_U318 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3994, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4000);
   dp_id_stage_regfile_DataPath_Physical_RF_U317 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3995, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4001);
   dp_id_stage_regfile_DataPath_Physical_RF_U316 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1156, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3903);
   dp_id_stage_regfile_DataPath_Physical_RF_U315 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1156, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3904);
   dp_id_stage_regfile_DataPath_Physical_RF_U314 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1156, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3905);
   dp_id_stage_regfile_DataPath_Physical_RF_U313 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1156, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3906);
   dp_id_stage_regfile_DataPath_Physical_RF_U312 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1156, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3907);
   dp_id_stage_regfile_DataPath_Physical_RF_U311 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1156, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3908);
   dp_id_stage_regfile_DataPath_Physical_RF_U310 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1155, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3914);
   dp_id_stage_regfile_DataPath_Physical_RF_U309 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1155, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3915);
   dp_id_stage_regfile_DataPath_Physical_RF_U308 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1155, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3916);
   dp_id_stage_regfile_DataPath_Physical_RF_U307 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1155, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3917);
   dp_id_stage_regfile_DataPath_Physical_RF_U306 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1155, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3918);
   dp_id_stage_regfile_DataPath_Physical_RF_U305 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1155, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3919);
   dp_id_stage_regfile_DataPath_Physical_RF_U304 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3903, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3909);
   dp_id_stage_regfile_DataPath_Physical_RF_U303 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3904, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3910);
   dp_id_stage_regfile_DataPath_Physical_RF_U302 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3914, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3920);
   dp_id_stage_regfile_DataPath_Physical_RF_U301 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3915, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3921);
   dp_id_stage_regfile_DataPath_Physical_RF_U300 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1154, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4085);
   dp_id_stage_regfile_DataPath_Physical_RF_U299 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1154, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4086);
   dp_id_stage_regfile_DataPath_Physical_RF_U298 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1154, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4087);
   dp_id_stage_regfile_DataPath_Physical_RF_U297 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1154, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4088);
   dp_id_stage_regfile_DataPath_Physical_RF_U296 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1154, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4089);
   dp_id_stage_regfile_DataPath_Physical_RF_U295 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1154, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4090);
   dp_id_stage_regfile_DataPath_Physical_RF_U294 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1, Z => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4096);
   dp_id_stage_regfile_DataPath_Physical_RF_U293 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1, Z => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4097);
   dp_id_stage_regfile_DataPath_Physical_RF_U292 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1, Z => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4098);
   dp_id_stage_regfile_DataPath_Physical_RF_U291 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1, Z => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4099);
   dp_id_stage_regfile_DataPath_Physical_RF_U290 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1, Z => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4100);
   dp_id_stage_regfile_DataPath_Physical_RF_U289 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1, Z => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4101);
   dp_id_stage_regfile_DataPath_Physical_RF_U288 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4085, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4091);
   dp_id_stage_regfile_DataPath_Physical_RF_U287 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4086, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4092);
   dp_id_stage_regfile_DataPath_Physical_RF_U286 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4096, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4102);
   dp_id_stage_regfile_DataPath_Physical_RF_U285 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4097, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4103);
   dp_id_stage_regfile_DataPath_Physical_RF_U284 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3864, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3861);
   dp_id_stage_regfile_DataPath_Physical_RF_U283 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3865, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3862);
   dp_id_stage_regfile_DataPath_Physical_RF_U282 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3866, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3863);
   dp_id_stage_regfile_DataPath_Physical_RF_U281 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1168, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3864);
   dp_id_stage_regfile_DataPath_Physical_RF_U280 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1168, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3865);
   dp_id_stage_regfile_DataPath_Physical_RF_U279 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1168, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3866);
   dp_id_stage_regfile_DataPath_Physical_RF_U278 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3967, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3964);
   dp_id_stage_regfile_DataPath_Physical_RF_U277 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3968, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3965);
   dp_id_stage_regfile_DataPath_Physical_RF_U276 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3969, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3966);
   dp_id_stage_regfile_DataPath_Physical_RF_U275 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1167, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3967);
   dp_id_stage_regfile_DataPath_Physical_RF_U274 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1167, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3968);
   dp_id_stage_regfile_DataPath_Physical_RF_U273 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1167, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3969);
   dp_id_stage_regfile_DataPath_Physical_RF_U272 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4048, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4045);
   dp_id_stage_regfile_DataPath_Physical_RF_U271 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4049, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4046);
   dp_id_stage_regfile_DataPath_Physical_RF_U270 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4050, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4047);
   dp_id_stage_regfile_DataPath_Physical_RF_U269 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1166, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4048);
   dp_id_stage_regfile_DataPath_Physical_RF_U268 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1166, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4049);
   dp_id_stage_regfile_DataPath_Physical_RF_U267 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1166, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4050);
   dp_id_stage_regfile_DataPath_Physical_RF_U266 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4059, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4056);
   dp_id_stage_regfile_DataPath_Physical_RF_U265 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4060, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4057);
   dp_id_stage_regfile_DataPath_Physical_RF_U264 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4061, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4058);
   dp_id_stage_regfile_DataPath_Physical_RF_U263 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1165, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4059);
   dp_id_stage_regfile_DataPath_Physical_RF_U262 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1165, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4060);
   dp_id_stage_regfile_DataPath_Physical_RF_U261 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1165, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4061);
   dp_id_stage_regfile_DataPath_Physical_RF_U260 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3875, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3872);
   dp_id_stage_regfile_DataPath_Physical_RF_U259 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3876, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3873);
   dp_id_stage_regfile_DataPath_Physical_RF_U258 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3877, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3874);
   dp_id_stage_regfile_DataPath_Physical_RF_U257 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1164, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3875);
   dp_id_stage_regfile_DataPath_Physical_RF_U256 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1164, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3876);
   dp_id_stage_regfile_DataPath_Physical_RF_U255 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1164, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3877);
   dp_id_stage_regfile_DataPath_Physical_RF_U254 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3956, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3953);
   dp_id_stage_regfile_DataPath_Physical_RF_U253 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3957, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3954);
   dp_id_stage_regfile_DataPath_Physical_RF_U252 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3958, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3955);
   dp_id_stage_regfile_DataPath_Physical_RF_U251 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1163, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3956);
   dp_id_stage_regfile_DataPath_Physical_RF_U250 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1163, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3957);
   dp_id_stage_regfile_DataPath_Physical_RF_U249 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1163, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3958);
   dp_id_stage_regfile_DataPath_Physical_RF_U248 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4192, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4189);
   dp_id_stage_regfile_DataPath_Physical_RF_U247 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4193, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4190);
   dp_id_stage_regfile_DataPath_Physical_RF_U246 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4194, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4191);
   dp_id_stage_regfile_DataPath_Physical_RF_U245 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1162, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4192);
   dp_id_stage_regfile_DataPath_Physical_RF_U244 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1162, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4193);
   dp_id_stage_regfile_DataPath_Physical_RF_U243 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1162, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4194);
   dp_id_stage_regfile_DataPath_Physical_RF_U242 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1161, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4186);
   dp_id_stage_regfile_DataPath_Physical_RF_U241 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1160, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4175);
   dp_id_stage_regfile_DataPath_Physical_RF_U240 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1159, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4164);
   dp_id_stage_regfile_DataPath_Physical_RF_U239 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1158, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4013);
   dp_id_stage_regfile_DataPath_Physical_RF_U238 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1157, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4002);
   dp_id_stage_regfile_DataPath_Physical_RF_U237 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1156, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3911);
   dp_id_stage_regfile_DataPath_Physical_RF_U236 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1155, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3922);
   dp_id_stage_regfile_DataPath_Physical_RF_U235 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1154, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4093);
   dp_id_stage_regfile_DataPath_Physical_RF_U234 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1, Z => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4104);
   dp_id_stage_regfile_DataPath_Physical_RF_U233 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1168, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3869);
   dp_id_stage_regfile_DataPath_Physical_RF_U232 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1167, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3972);
   dp_id_stage_regfile_DataPath_Physical_RF_U231 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1166, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4053);
   dp_id_stage_regfile_DataPath_Physical_RF_U230 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1165, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4064);
   dp_id_stage_regfile_DataPath_Physical_RF_U229 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1164, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3880);
   dp_id_stage_regfile_DataPath_Physical_RF_U228 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1163, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3961);
   dp_id_stage_regfile_DataPath_Physical_RF_U227 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1162, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4197);
   dp_id_stage_regfile_DataPath_Physical_RF_U226 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4227, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4219);
   dp_id_stage_regfile_DataPath_Physical_RF_U225 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4227, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4218);
   dp_id_stage_regfile_DataPath_Physical_RF_U224 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4022, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4015);
   dp_id_stage_regfile_DataPath_Physical_RF_U223 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4022, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4014);
   dp_id_stage_regfile_DataPath_Physical_RF_U222 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4153, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4146);
   dp_id_stage_regfile_DataPath_Physical_RF_U221 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4153, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4145);
   dp_id_stage_regfile_DataPath_Physical_RF_U220 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3991, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3984);
   dp_id_stage_regfile_DataPath_Physical_RF_U219 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3991, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3983);
   dp_id_stage_regfile_DataPath_Physical_RF_U218 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3931, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3924);
   dp_id_stage_regfile_DataPath_Physical_RF_U217 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3931, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3923);
   dp_id_stage_regfile_DataPath_Physical_RF_U216 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3940, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3933);
   dp_id_stage_regfile_DataPath_Physical_RF_U215 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3940, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3932);
   dp_id_stage_regfile_DataPath_Physical_RF_U214 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4073, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4066);
   dp_id_stage_regfile_DataPath_Physical_RF_U213 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4073, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4065);
   dp_id_stage_regfile_DataPath_Physical_RF_U212 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4082, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4075);
   dp_id_stage_regfile_DataPath_Physical_RF_U211 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4082, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4074);
   dp_id_stage_regfile_DataPath_Physical_RF_U210 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3950, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3942);
   dp_id_stage_regfile_DataPath_Physical_RF_U209 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3950, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3941);
   dp_id_stage_regfile_DataPath_Physical_RF_U208 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4032, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4024);
   dp_id_stage_regfile_DataPath_Physical_RF_U207 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4032, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4023);
   dp_id_stage_regfile_DataPath_Physical_RF_U206 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4114, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4106);
   dp_id_stage_regfile_DataPath_Physical_RF_U205 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4114, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4105);
   dp_id_stage_regfile_DataPath_Physical_RF_U204 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3890, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3882);
   dp_id_stage_regfile_DataPath_Physical_RF_U203 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3890, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3881);
   dp_id_stage_regfile_DataPath_Physical_RF_U202 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3900, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3892);
   dp_id_stage_regfile_DataPath_Physical_RF_U201 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3900, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3891);
   dp_id_stage_regfile_DataPath_Physical_RF_U200 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3982, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3974);
   dp_id_stage_regfile_DataPath_Physical_RF_U199 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3982, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3973);
   dp_id_stage_regfile_DataPath_Physical_RF_U198 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4134, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4126);
   dp_id_stage_regfile_DataPath_Physical_RF_U197 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4134, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4125);
   dp_id_stage_regfile_DataPath_Physical_RF_U196 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4144, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4136);
   dp_id_stage_regfile_DataPath_Physical_RF_U195 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4144, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4135);
   dp_id_stage_regfile_DataPath_Physical_RF_U194 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4042, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4034);
   dp_id_stage_regfile_DataPath_Physical_RF_U193 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4042, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4033);
   dp_id_stage_regfile_DataPath_Physical_RF_U192 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4124, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4116);
   dp_id_stage_regfile_DataPath_Physical_RF_U191 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4124, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4115);
   dp_id_stage_regfile_DataPath_Physical_RF_U190 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4217, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4209);
   dp_id_stage_regfile_DataPath_Physical_RF_U189 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4217, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4208);
   dp_id_stage_regfile_DataPath_Physical_RF_U188 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4207, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4199);
   dp_id_stage_regfile_DataPath_Physical_RF_U187 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4207, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4198);
   dp_id_stage_regfile_DataPath_Physical_RF_U186 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1169, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1189);
   dp_id_stage_regfile_DataPath_Physical_RF_U185 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1170, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1200);
   dp_id_stage_regfile_DataPath_Physical_RF_U184 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1171, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1202);
   dp_id_stage_regfile_DataPath_Physical_RF_U183 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2601, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1220);
   dp_id_stage_regfile_DataPath_Physical_RF_U182 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2575, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3714);
   dp_id_stage_regfile_DataPath_Physical_RF_U181 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2560, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3750);
   dp_id_stage_regfile_DataPath_Physical_RF_U180 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2601, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1219);
   dp_id_stage_regfile_DataPath_Physical_RF_U179 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2575, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3713);
   dp_id_stage_regfile_DataPath_Physical_RF_U178 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2601, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n1218);
   dp_id_stage_regfile_DataPath_Physical_RF_U177 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2575, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3712);
   dp_id_stage_regfile_DataPath_Physical_RF_U176 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2560, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3748);
   dp_id_stage_regfile_DataPath_Physical_RF_U175 : BUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2560, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3749);
   dp_id_stage_regfile_DataPath_Physical_RF_U174 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4186, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4176);
   dp_id_stage_regfile_DataPath_Physical_RF_U173 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4186, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4177);
   dp_id_stage_regfile_DataPath_Physical_RF_U172 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4175, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4165);
   dp_id_stage_regfile_DataPath_Physical_RF_U171 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4175, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4166);
   dp_id_stage_regfile_DataPath_Physical_RF_U170 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4164, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4154);
   dp_id_stage_regfile_DataPath_Physical_RF_U169 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4164, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4155);
   dp_id_stage_regfile_DataPath_Physical_RF_U168 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4013, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4003);
   dp_id_stage_regfile_DataPath_Physical_RF_U167 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4013, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4004);
   dp_id_stage_regfile_DataPath_Physical_RF_U166 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4002, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3992);
   dp_id_stage_regfile_DataPath_Physical_RF_U165 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4002, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3993);
   dp_id_stage_regfile_DataPath_Physical_RF_U164 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3911, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3901);
   dp_id_stage_regfile_DataPath_Physical_RF_U163 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3911, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3902);
   dp_id_stage_regfile_DataPath_Physical_RF_U162 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3922, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3912);
   dp_id_stage_regfile_DataPath_Physical_RF_U161 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3922, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3913);
   dp_id_stage_regfile_DataPath_Physical_RF_U160 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4093, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4083);
   dp_id_stage_regfile_DataPath_Physical_RF_U159 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4093, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4084);
   dp_id_stage_regfile_DataPath_Physical_RF_U158 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4104, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4094);
   dp_id_stage_regfile_DataPath_Physical_RF_U157 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4104, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4095);
   dp_id_stage_regfile_DataPath_Physical_RF_U156 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3869, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3859);
   dp_id_stage_regfile_DataPath_Physical_RF_U155 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3869, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3860);
   dp_id_stage_regfile_DataPath_Physical_RF_U154 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3972, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3962);
   dp_id_stage_regfile_DataPath_Physical_RF_U153 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3972, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3963);
   dp_id_stage_regfile_DataPath_Physical_RF_U152 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4053, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4043);
   dp_id_stage_regfile_DataPath_Physical_RF_U151 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4053, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4044);
   dp_id_stage_regfile_DataPath_Physical_RF_U150 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4064, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4054);
   dp_id_stage_regfile_DataPath_Physical_RF_U149 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4064, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4055);
   dp_id_stage_regfile_DataPath_Physical_RF_U148 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3880, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3870);
   dp_id_stage_regfile_DataPath_Physical_RF_U147 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3880, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3871);
   dp_id_stage_regfile_DataPath_Physical_RF_U146 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3961, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3951);
   dp_id_stage_regfile_DataPath_Physical_RF_U145 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3961, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3952);
   dp_id_stage_regfile_DataPath_Physical_RF_U144 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4197, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4187);
   dp_id_stage_regfile_DataPath_Physical_RF_U143 : INV_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4197, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n4188);
   dp_id_stage_regfile_DataPath_Physical_RF_U142 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4236, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2532
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U141 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4270, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n2530
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U140 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1198, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_0_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3159
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U139 : NOR2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1199, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_1_port, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n3157
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U138 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1825, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3930);
   dp_id_stage_regfile_DataPath_Physical_RF_U137 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1825, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3929);
   dp_id_stage_regfile_DataPath_Physical_RF_U136 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1825, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3928);
   dp_id_stage_regfile_DataPath_Physical_RF_U135 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1825, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3927);
   dp_id_stage_regfile_DataPath_Physical_RF_U134 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1825, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3926);
   dp_id_stage_regfile_DataPath_Physical_RF_U133 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1825, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3925);
   dp_id_stage_regfile_DataPath_Physical_RF_U132 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1791, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3939);
   dp_id_stage_regfile_DataPath_Physical_RF_U131 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1791, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3938);
   dp_id_stage_regfile_DataPath_Physical_RF_U130 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1791, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3937);
   dp_id_stage_regfile_DataPath_Physical_RF_U129 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1791, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3936);
   dp_id_stage_regfile_DataPath_Physical_RF_U128 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1791, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3935);
   dp_id_stage_regfile_DataPath_Physical_RF_U127 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1791, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3934);
   dp_id_stage_regfile_DataPath_Physical_RF_U126 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1553, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4072);
   dp_id_stage_regfile_DataPath_Physical_RF_U125 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1553, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4071);
   dp_id_stage_regfile_DataPath_Physical_RF_U124 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1553, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4070);
   dp_id_stage_regfile_DataPath_Physical_RF_U123 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1553, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4069);
   dp_id_stage_regfile_DataPath_Physical_RF_U122 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1553, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4068);
   dp_id_stage_regfile_DataPath_Physical_RF_U121 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1553, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4067);
   dp_id_stage_regfile_DataPath_Physical_RF_U120 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1520, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4081);
   dp_id_stage_regfile_DataPath_Physical_RF_U119 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1520, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4080);
   dp_id_stage_regfile_DataPath_Physical_RF_U118 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1520, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4079);
   dp_id_stage_regfile_DataPath_Physical_RF_U117 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1520, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4078);
   dp_id_stage_regfile_DataPath_Physical_RF_U116 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1520, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4077);
   dp_id_stage_regfile_DataPath_Physical_RF_U115 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1520, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4076);
   dp_id_stage_regfile_DataPath_Physical_RF_U114 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1758, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3949);
   dp_id_stage_regfile_DataPath_Physical_RF_U113 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1758, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3948);
   dp_id_stage_regfile_DataPath_Physical_RF_U112 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1758, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3947);
   dp_id_stage_regfile_DataPath_Physical_RF_U111 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1758, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3946);
   dp_id_stage_regfile_DataPath_Physical_RF_U110 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1758, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3945);
   dp_id_stage_regfile_DataPath_Physical_RF_U109 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1758, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3944);
   dp_id_stage_regfile_DataPath_Physical_RF_U108 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1621, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4031);
   dp_id_stage_regfile_DataPath_Physical_RF_U107 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1621, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4030);
   dp_id_stage_regfile_DataPath_Physical_RF_U106 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1621, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4029);
   dp_id_stage_regfile_DataPath_Physical_RF_U105 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1621, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4028);
   dp_id_stage_regfile_DataPath_Physical_RF_U104 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1621, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4027);
   dp_id_stage_regfile_DataPath_Physical_RF_U103 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1621, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4026);
   dp_id_stage_regfile_DataPath_Physical_RF_U102 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1484, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4113);
   dp_id_stage_regfile_DataPath_Physical_RF_U101 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1484, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4112);
   dp_id_stage_regfile_DataPath_Physical_RF_U100 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1484, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4111);
   dp_id_stage_regfile_DataPath_Physical_RF_U99 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1484, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4110);
   dp_id_stage_regfile_DataPath_Physical_RF_U98 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1484, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4109);
   dp_id_stage_regfile_DataPath_Physical_RF_U97 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1484, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4108);
   dp_id_stage_regfile_DataPath_Physical_RF_U96 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1893, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3889);
   dp_id_stage_regfile_DataPath_Physical_RF_U95 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1893, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3888);
   dp_id_stage_regfile_DataPath_Physical_RF_U94 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1893, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3887);
   dp_id_stage_regfile_DataPath_Physical_RF_U93 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1893, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3886);
   dp_id_stage_regfile_DataPath_Physical_RF_U92 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1893, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3885);
   dp_id_stage_regfile_DataPath_Physical_RF_U91 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1893, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3884);
   dp_id_stage_regfile_DataPath_Physical_RF_U90 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1860, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3899);
   dp_id_stage_regfile_DataPath_Physical_RF_U89 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1860, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3898);
   dp_id_stage_regfile_DataPath_Physical_RF_U88 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1860, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3897);
   dp_id_stage_regfile_DataPath_Physical_RF_U87 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1860, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3896);
   dp_id_stage_regfile_DataPath_Physical_RF_U86 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1860, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3895);
   dp_id_stage_regfile_DataPath_Physical_RF_U85 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1860, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3894);
   dp_id_stage_regfile_DataPath_Physical_RF_U84 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1723, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3981);
   dp_id_stage_regfile_DataPath_Physical_RF_U83 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1723, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3980);
   dp_id_stage_regfile_DataPath_Physical_RF_U82 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1723, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3979);
   dp_id_stage_regfile_DataPath_Physical_RF_U81 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1723, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3978);
   dp_id_stage_regfile_DataPath_Physical_RF_U80 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1723, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3977);
   dp_id_stage_regfile_DataPath_Physical_RF_U79 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1723, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3976);
   dp_id_stage_regfile_DataPath_Physical_RF_U78 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1418, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4133);
   dp_id_stage_regfile_DataPath_Physical_RF_U77 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1418, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4132);
   dp_id_stage_regfile_DataPath_Physical_RF_U76 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1418, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4131);
   dp_id_stage_regfile_DataPath_Physical_RF_U75 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1418, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4130);
   dp_id_stage_regfile_DataPath_Physical_RF_U74 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1418, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4129);
   dp_id_stage_regfile_DataPath_Physical_RF_U73 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1418, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4128);
   dp_id_stage_regfile_DataPath_Physical_RF_U72 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1385, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4143);
   dp_id_stage_regfile_DataPath_Physical_RF_U71 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1385, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4142);
   dp_id_stage_regfile_DataPath_Physical_RF_U70 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1385, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4141);
   dp_id_stage_regfile_DataPath_Physical_RF_U69 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1385, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4140);
   dp_id_stage_regfile_DataPath_Physical_RF_U68 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1385, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4139);
   dp_id_stage_regfile_DataPath_Physical_RF_U67 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1385, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4138);
   dp_id_stage_regfile_DataPath_Physical_RF_U66 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1588, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4041);
   dp_id_stage_regfile_DataPath_Physical_RF_U65 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1588, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4040);
   dp_id_stage_regfile_DataPath_Physical_RF_U64 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1588, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4039);
   dp_id_stage_regfile_DataPath_Physical_RF_U63 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1588, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4038);
   dp_id_stage_regfile_DataPath_Physical_RF_U62 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1588, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4037);
   dp_id_stage_regfile_DataPath_Physical_RF_U61 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1588, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4036);
   dp_id_stage_regfile_DataPath_Physical_RF_U60 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1451, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4123);
   dp_id_stage_regfile_DataPath_Physical_RF_U59 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1451, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4122);
   dp_id_stage_regfile_DataPath_Physical_RF_U58 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1451, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4121);
   dp_id_stage_regfile_DataPath_Physical_RF_U57 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1451, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4120);
   dp_id_stage_regfile_DataPath_Physical_RF_U56 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1451, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4119);
   dp_id_stage_regfile_DataPath_Physical_RF_U55 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1451, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4118);
   dp_id_stage_regfile_DataPath_Physical_RF_U54 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1273, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4216);
   dp_id_stage_regfile_DataPath_Physical_RF_U53 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1273, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4215);
   dp_id_stage_regfile_DataPath_Physical_RF_U52 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1273, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4214);
   dp_id_stage_regfile_DataPath_Physical_RF_U51 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1273, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4213);
   dp_id_stage_regfile_DataPath_Physical_RF_U50 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1273, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4212);
   dp_id_stage_regfile_DataPath_Physical_RF_U49 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1273, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4211);
   dp_id_stage_regfile_DataPath_Physical_RF_U48 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1307, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4204);
   dp_id_stage_regfile_DataPath_Physical_RF_U47 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1307, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4203);
   dp_id_stage_regfile_DataPath_Physical_RF_U46 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1307, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4202);
   dp_id_stage_regfile_DataPath_Physical_RF_U45 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1307, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4201);
   dp_id_stage_regfile_DataPath_Physical_RF_U44 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1238, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4226);
   dp_id_stage_regfile_DataPath_Physical_RF_U43 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1238, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4225);
   dp_id_stage_regfile_DataPath_Physical_RF_U42 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1238, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4224);
   dp_id_stage_regfile_DataPath_Physical_RF_U41 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1238, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4223);
   dp_id_stage_regfile_DataPath_Physical_RF_U40 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1238, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4222);
   dp_id_stage_regfile_DataPath_Physical_RF_U39 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1238, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4221);
   dp_id_stage_regfile_DataPath_Physical_RF_U38 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1307, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4205);
   dp_id_stage_regfile_DataPath_Physical_RF_U37 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1307, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4206);
   dp_id_stage_regfile_DataPath_Physical_RF_U36 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1168, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3867);
   dp_id_stage_regfile_DataPath_Physical_RF_U35 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1168, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3868);
   dp_id_stage_regfile_DataPath_Physical_RF_U34 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1167, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3970);
   dp_id_stage_regfile_DataPath_Physical_RF_U33 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1167, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3971);
   dp_id_stage_regfile_DataPath_Physical_RF_U32 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1166, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4051);
   dp_id_stage_regfile_DataPath_Physical_RF_U31 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1166, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4052);
   dp_id_stage_regfile_DataPath_Physical_RF_U30 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1165, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4062);
   dp_id_stage_regfile_DataPath_Physical_RF_U29 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1165, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4063);
   dp_id_stage_regfile_DataPath_Physical_RF_U28 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1164, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3878);
   dp_id_stage_regfile_DataPath_Physical_RF_U27 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1164, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3879);
   dp_id_stage_regfile_DataPath_Physical_RF_U26 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1163, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3959);
   dp_id_stage_regfile_DataPath_Physical_RF_U25 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1163, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n3960);
   dp_id_stage_regfile_DataPath_Physical_RF_U24 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1162, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4195);
   dp_id_stage_regfile_DataPath_Physical_RF_U23 : CLKBUF_X1 port map( A => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1162, Z =>
                           dp_id_stage_regfile_DataPath_Physical_RF_n4196);
   dp_id_stage_regfile_DataPath_Physical_RF_U22 : INV_X32 port map( A => 
                           dp_id_stage_regfile_rst_rf, ZN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237);
   dp_id_stage_regfile_DataPath_Physical_RF_U21 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1823, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1341, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1168
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U20 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1686, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1305, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1167
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U19 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1517, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1305, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1166
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U18 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1517, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1270, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1165
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U17 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1823, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1339, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1164
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U16 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1686, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1339, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1163
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U15 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1341, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1271, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1162
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U14 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1344, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1345, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1161
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U13 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1347, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1345, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1160
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U12 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1349, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1345, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1159
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U11 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1686, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1347, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1158
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U10 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1686, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1349, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1157
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U9 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1823, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1383, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1156
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U8 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1823, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1349, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1155
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U7 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1517, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1347, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1154
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_U6 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1517, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1344, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1);
   dp_id_stage_regfile_DataPath_Physical_RF_U5 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_2_port, A2 
                           => dp_id_stage_regfile_DataPath_addr_rd2_p_3_port, 
                           A3 => dp_id_stage_regfile_DataPath_addr_rd2_p_4_port
                           , A4 => 
                           dp_id_stage_regfile_DataPath_addr_rd2_p_5_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n2546);
   dp_id_stage_regfile_DataPath_Physical_RF_U4 : NOR4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_2_port, A2 
                           => dp_id_stage_regfile_DataPath_mux_rd_out_3_port, 
                           A3 => dp_id_stage_regfile_DataPath_mux_rd_out_4_port
                           , A4 => 
                           dp_id_stage_regfile_DataPath_mux_rd_out_5_port, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n3173);
   dp_id_stage_regfile_DataPath_Physical_RF_U3 : AND4_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_out_5_port, A2 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1342, 
                           A3 => dp_id_stage_regfile_DataPath_Physical_RF_n1192
                           , A4 => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1191, ZN 
                           => dp_id_stage_regfile_DataPath_Physical_RF_n1271);
   dp_id_stage_regfile_DataPath_Physical_RF_U2 : AND2_X1 port map( A1 => 
                           dp_id_stage_regfile_DataPath_mux_wr_control_out, A2 
                           => dp_id_stage_regfile_DataPath_mux_en_control_out, 
                           ZN => dp_id_stage_regfile_DataPath_Physical_RF_n1342
                           );
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1089, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_0_port, 
                           QN => n_1161);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1079, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_10_port, 
                           QN => n_1162);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1078, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_11_port, 
                           QN => n_1163);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1077, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_12_port, 
                           QN => n_1164);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1076, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_13_port, 
                           QN => n_1165);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1075, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_14_port, 
                           QN => n_1166);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1074, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_15_port, 
                           QN => n_1167);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1073, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_16_port, 
                           QN => n_1168);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1121, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_0_port, 
                           QN => n_1169);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1111, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_10_port, 
                           QN => n_1170);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1110, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_11_port, 
                           QN => n_1171);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1109, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_12_port, 
                           QN => n_1172);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1108, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_13_port, 
                           QN => n_1173);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1107, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_14_port, 
                           QN => n_1174);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1106, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_15_port, 
                           QN => n_1175);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1105, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_16_port, 
                           QN => n_1176);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1088, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_1_port, 
                           QN => n_1177);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1087, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_2_port, 
                           QN => n_1178);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1086, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_3_port, 
                           QN => n_1179);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1085, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_4_port, 
                           QN => n_1180);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1084, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_5_port, 
                           QN => n_1181);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1083, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_6_port, 
                           QN => n_1182);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1082, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_7_port, 
                           QN => n_1183);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1081, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_8_port, 
                           QN => n_1184);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1080, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_9_port, 
                           QN => n_1185);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1072, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_17_port, 
                           QN => n_1186);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1071, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_18_port, 
                           QN => n_1187);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1070, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_19_port, 
                           QN => n_1188);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1069, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_20_port, 
                           QN => n_1189);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1068, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_21_port, 
                           QN => n_1190);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1067, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_22_port, 
                           QN => n_1191);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1066, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_23_port, 
                           QN => n_1192);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1120, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_1_port, 
                           QN => n_1193);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1119, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_2_port, 
                           QN => n_1194);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1118, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_3_port, 
                           QN => n_1195);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1117, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_4_port, 
                           QN => n_1196);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1116, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_5_port, 
                           QN => n_1197);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1115, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_6_port, 
                           QN => n_1198);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1114, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_7_port, 
                           QN => n_1199);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1113, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_8_port, 
                           QN => n_1200);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1112, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_9_port, 
                           QN => n_1201);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1104, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_17_port, 
                           QN => n_1202);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1103, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_18_port, 
                           QN => n_1203);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1102, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_19_port, 
                           QN => n_1204);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1101, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_20_port, 
                           QN => n_1205);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1100, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_21_port, 
                           QN => n_1206);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1099, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_22_port, 
                           QN => n_1207);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1098, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_23_port, 
                           QN => n_1208);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1153, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_0_port, 
                           QN => n_1209);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1152, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_1_port, 
                           QN => n_1210);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1151, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_2_port, 
                           QN => n_1211);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1150, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_3_port, 
                           QN => n_1212);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1149, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_4_port, 
                           QN => n_1213);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1148, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_5_port, 
                           QN => n_1214);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1147, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_6_port, 
                           QN => n_1215);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1146, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_7_port, 
                           QN => n_1216);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1145, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_8_port, 
                           QN => n_1217);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1144, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_9_port, 
                           QN => n_1218);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1143, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_10_port, 
                           QN => n_1219);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1142, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_11_port, 
                           QN => n_1220);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1141, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_12_port, 
                           QN => n_1221);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1140, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_13_port, 
                           QN => n_1222);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1139, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_14_port, 
                           QN => n_1223);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1138, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_15_port, 
                           QN => n_1224);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1137, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_16_port, 
                           QN => n_1225);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1136, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_17_port, 
                           QN => n_1226);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1135, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_18_port, 
                           QN => n_1227);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1134, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_19_port, 
                           QN => n_1228);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1133, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_20_port, 
                           QN => n_1229);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1132, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_21_port, 
                           QN => n_1230);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1131, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_22_port, 
                           QN => n_1231);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1130, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_23_port, 
                           QN => n_1232);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n577, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_0_port, 
                           QN => n_1233);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n567, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_10_port, 
                           QN => n_1234);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n566, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_11_port, 
                           QN => n_1235);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n565, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_12_port, 
                           QN => n_1236);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n564, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_13_port, 
                           QN => n_1237);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n563, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_14_port, 
                           QN => n_1238);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n562, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_15_port, 
                           QN => n_1239);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n561, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_16_port, 
                           QN => n_1240);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n833, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_0_port, 
                           QN => n_1241);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n823, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_10_port, 
                           QN => n_1242);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n822, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_11_port, 
                           QN => n_1243);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n821, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_12_port, 
                           QN => n_1244);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n820, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_13_port, 
                           QN => n_1245);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n819, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_14_port, 
                           QN => n_1246);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n818, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_15_port, 
                           QN => n_1247);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n817, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_16_port, 
                           QN => n_1248);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n97, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_0_port, 
                           QN => n_1249);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n87, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_10_port, 
                           QN => n_1250);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n86, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_11_port, 
                           QN => n_1251);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n85, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_12_port, 
                           QN => n_1252);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n84, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_13_port, 
                           QN => n_1253);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n83, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_14_port, 
                           QN => n_1254);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n82, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_15_port, 
                           QN => n_1255);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n81, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_16_port, 
                           QN => n_1256);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n129, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_0_port, 
                           QN => n_1257);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n119, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_10_port, 
                           QN => n_1258);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n118, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_11_port, 
                           QN => n_1259);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n117, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_12_port, 
                           QN => n_1260);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n116, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_13_port, 
                           QN => n_1261);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n115, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_14_port, 
                           QN => n_1262);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n114, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_15_port, 
                           QN => n_1263);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n113, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_16_port, 
                           QN => n_1264);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n385, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_0_port, 
                           QN => n_1265);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n375, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_10_port, 
                           QN => n_1266);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n374, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_11_port, 
                           QN => n_1267);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n373, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_12_port, 
                           QN => n_1268);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n372, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_13_port, 
                           QN => n_1269);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n371, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_14_port, 
                           QN => n_1270);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n370, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_15_port, 
                           QN => n_1271);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n369, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_16_port, 
                           QN => n_1272);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n865, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_0_port, 
                           QN => n_1273);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n855, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_10_port, 
                           QN => n_1274);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n854, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_11_port, 
                           QN => n_1275);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n853, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_12_port, 
                           QN => n_1276);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n852, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_13_port, 
                           QN => n_1277);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n851, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_14_port, 
                           QN => n_1278);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n850, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_15_port, 
                           QN => n_1279);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n849, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_16_port, 
                           QN => n_1280);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n897, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_0_port, 
                           QN => n_1281);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n887, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_10_port, 
                           QN => n_1282);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n886, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_11_port, 
                           QN => n_1283);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n885, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_12_port, 
                           QN => n_1284);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n884, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_13_port, 
                           QN => n_1285);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n883, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_14_port, 
                           QN => n_1286);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n882, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_15_port, 
                           QN => n_1287);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n881, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_16_port, 
                           QN => n_1288);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n576, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_1_port, 
                           QN => n_1289);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n575, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_2_port, 
                           QN => n_1290);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n574, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_3_port, 
                           QN => n_1291);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n573, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_4_port, 
                           QN => n_1292);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n572, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_5_port, 
                           QN => n_1293);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n571, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_6_port, 
                           QN => n_1294);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n570, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_7_port, 
                           QN => n_1295);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n569, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_8_port, 
                           QN => n_1296);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n568, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_9_port, 
                           QN => n_1297);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n560, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_17_port, 
                           QN => n_1298);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n559, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_18_port, 
                           QN => n_1299);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n558, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_19_port, 
                           QN => n_1300);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n557, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_20_port, 
                           QN => n_1301);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n556, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_21_port, 
                           QN => n_1302);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n555, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_22_port, 
                           QN => n_1303);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n554, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_23_port, 
                           QN => n_1304);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n832, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_1_port, 
                           QN => n_1305);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n831, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_2_port, 
                           QN => n_1306);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n830, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_3_port, 
                           QN => n_1307);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n829, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_4_port, 
                           QN => n_1308);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n828, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_5_port, 
                           QN => n_1309);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n827, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_6_port, 
                           QN => n_1310);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n826, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_7_port, 
                           QN => n_1311);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n825, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_8_port, 
                           QN => n_1312);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n824, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_9_port, 
                           QN => n_1313);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n816, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_17_port, 
                           QN => n_1314);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n815, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_18_port, 
                           QN => n_1315);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n814, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_19_port, 
                           QN => n_1316);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n813, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_20_port, 
                           QN => n_1317);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n812, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_21_port, 
                           QN => n_1318);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n811, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_22_port, 
                           QN => n_1319);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n810, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_23_port, 
                           QN => n_1320);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n96, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_1_port, 
                           QN => n_1321);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n95, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_2_port, 
                           QN => n_1322);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n94, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_3_port, 
                           QN => n_1323);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n93, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_4_port, 
                           QN => n_1324);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n92, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_5_port, 
                           QN => n_1325);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n91, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_6_port, 
                           QN => n_1326);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n90, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_7_port, 
                           QN => n_1327);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n89, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_8_port, 
                           QN => n_1328);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n88, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_9_port, 
                           QN => n_1329);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n80, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_17_port, 
                           QN => n_1330);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n79, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_18_port, 
                           QN => n_1331);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n78, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_19_port, 
                           QN => n_1332);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n77, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_20_port, 
                           QN => n_1333);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n76, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_21_port, 
                           QN => n_1334);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n75, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_22_port, 
                           QN => n_1335);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n74, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_23_port, 
                           QN => n_1336);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n128, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_1_port, 
                           QN => n_1337);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n127, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_2_port, 
                           QN => n_1338);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n126, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_3_port, 
                           QN => n_1339);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n125, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_4_port, 
                           QN => n_1340);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n124, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_5_port, 
                           QN => n_1341);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n123, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_6_port, 
                           QN => n_1342);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n122, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_7_port, 
                           QN => n_1343);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n121, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_8_port, 
                           QN => n_1344);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n120, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_9_port, 
                           QN => n_1345);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n112, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_17_port, 
                           QN => n_1346);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n111, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_18_port, 
                           QN => n_1347);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n110, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_19_port, 
                           QN => n_1348);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n109, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_20_port, 
                           QN => n_1349);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n108, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_21_port, 
                           QN => n_1350);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n107, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_22_port, 
                           QN => n_1351);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n106, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_23_port, 
                           QN => n_1352);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n384, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_1_port, 
                           QN => n_1353);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n383, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_2_port, 
                           QN => n_1354);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n382, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_3_port, 
                           QN => n_1355);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n381, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_4_port, 
                           QN => n_1356);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n380, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_5_port, 
                           QN => n_1357);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n379, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_6_port, 
                           QN => n_1358);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n378, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_7_port, 
                           QN => n_1359);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n377, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_8_port, 
                           QN => n_1360);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n376, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_9_port, 
                           QN => n_1361);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n368, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_17_port, 
                           QN => n_1362);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n367, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_18_port, 
                           QN => n_1363);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n366, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_19_port, 
                           QN => n_1364);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n365, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_20_port, 
                           QN => n_1365);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n364, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_21_port, 
                           QN => n_1366);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n363, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_22_port, 
                           QN => n_1367);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n362, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_23_port, 
                           QN => n_1368);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n864, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_1_port, 
                           QN => n_1369);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n863, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_2_port, 
                           QN => n_1370);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n862, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_3_port, 
                           QN => n_1371);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n861, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_4_port, 
                           QN => n_1372);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n860, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_5_port, 
                           QN => n_1373);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n859, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_6_port, 
                           QN => n_1374);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n858, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_7_port, 
                           QN => n_1375);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n857, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_8_port, 
                           QN => n_1376);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n856, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_9_port, 
                           QN => n_1377);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n848, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_17_port, 
                           QN => n_1378);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n847, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_18_port, 
                           QN => n_1379);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n846, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_19_port, 
                           QN => n_1380);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n845, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_20_port, 
                           QN => n_1381);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n844, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_21_port, 
                           QN => n_1382);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n843, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_22_port, 
                           QN => n_1383);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n842, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_23_port, 
                           QN => n_1384);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n896, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_1_port, 
                           QN => n_1385);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n895, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_2_port, 
                           QN => n_1386);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n894, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_3_port, 
                           QN => n_1387);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n893, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_4_port, 
                           QN => n_1388);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n892, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_5_port, 
                           QN => n_1389);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n891, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_6_port, 
                           QN => n_1390);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n890, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_7_port, 
                           QN => n_1391);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n889, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_8_port, 
                           QN => n_1392);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n888, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_9_port, 
                           QN => n_1393);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n880, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_17_port, 
                           QN => n_1394);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n879, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_18_port, 
                           QN => n_1395);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n878, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_19_port, 
                           QN => n_1396);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n877, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_20_port, 
                           QN => n_1397);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n876, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_21_port, 
                           QN => n_1398);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n875, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_22_port, 
                           QN => n_1399);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n874, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_23_port, 
                           QN => n_1400);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1063, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_26_port, 
                           QN => n_1401);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1062, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_27_port, 
                           QN => n_1402);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1059, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_30_port, 
                           QN => n_1403);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1058, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_31_port, 
                           QN => n_1404);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1095, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_26_port, 
                           QN => n_1405);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1094, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_27_port, 
                           QN => n_1406);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1091, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_30_port, 
                           QN => n_1407);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1090, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_31_port, 
                           QN => n_1408);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1127, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_26_port, 
                           QN => n_1409);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1126, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_27_port, 
                           QN => n_1410);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1123, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_30_port, 
                           QN => n_1411);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1122, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_31_port, 
                           QN => n_1412);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1065, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_24_port, 
                           QN => n_1413);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1064, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_25_port, 
                           QN => n_1414);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1061, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_28_port, 
                           QN => n_1415);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_33_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1060, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_33_29_port, 
                           QN => n_1416);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1097, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_24_port, 
                           QN => n_1417);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1096, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_25_port, 
                           QN => n_1418);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1093, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_28_port, 
                           QN => n_1419);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_34_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1092, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_34_29_port, 
                           QN => n_1420);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n551, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_26_port, 
                           QN => n_1421);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n550, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_27_port, 
                           QN => n_1422);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n547, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_30_port, 
                           QN => n_1423);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n546, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_31_port, 
                           QN => n_1424);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n807, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_26_port, 
                           QN => n_1425);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n806, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_27_port, 
                           QN => n_1426);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n803, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_30_port, 
                           QN => n_1427);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n802, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_31_port, 
                           QN => n_1428);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n71, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_26_port, 
                           QN => n_1429);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n70, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_27_port, 
                           QN => n_1430);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n67, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_30_port, 
                           QN => n_1431);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n66, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_31_port, 
                           QN => n_1432);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n103, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_26_port, 
                           QN => n_1433);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n102, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_27_port, 
                           QN => n_1434);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n99, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_30_port, 
                           QN => n_1435);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n98, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_31_port, 
                           QN => n_1436);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n359, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_26_port, 
                           QN => n_1437);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n358, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_27_port, 
                           QN => n_1438);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n355, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_30_port, 
                           QN => n_1439);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n354, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_31_port, 
                           QN => n_1440);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n839, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_26_port, 
                           QN => n_1441);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n838, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_27_port, 
                           QN => n_1442);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n835, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_30_port, 
                           QN => n_1443);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n834, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_31_port, 
                           QN => n_1444);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n871, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_26_port, 
                           QN => n_1445);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n870, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_27_port, 
                           QN => n_1446);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n867, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_30_port, 
                           QN => n_1447);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n866, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_31_port, 
                           QN => n_1448);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1129, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_24_port, 
                           QN => n_1449);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1128, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_25_port, 
                           QN => n_1450);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1125, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_28_port, 
                           QN => n_1451);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_35_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1124, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_35_29_port, 
                           QN => n_1452);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n289, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_0_port, 
                           QN => n_1453);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n279, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_10_port, 
                           QN => n_1454);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n278, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_11_port, 
                           QN => n_1455);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n277, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_12_port, 
                           QN => n_1456);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n276, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_13_port, 
                           QN => n_1457);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n275, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_14_port, 
                           QN => n_1458);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n274, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_15_port, 
                           QN => n_1459);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n273, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_16_port, 
                           QN => n_1460);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n545, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_0_port, 
                           QN => n_1461);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n535, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_10_port, 
                           QN => n_1462);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n534, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_11_port, 
                           QN => n_1463);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n533, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_12_port, 
                           QN => n_1464);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n532, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_13_port, 
                           QN => n_1465);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n531, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_14_port, 
                           QN => n_1466);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n530, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_15_port, 
                           QN => n_1467);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n529, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_16_port, 
                           QN => n_1468);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n801, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_0_port, 
                           QN => n_1469);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n791, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_10_port, 
                           QN => n_1470);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n790, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_11_port, 
                           QN => n_1471);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n789, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_12_port, 
                           QN => n_1472);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n788, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_13_port, 
                           QN => n_1473);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n787, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_14_port, 
                           QN => n_1474);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n786, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_15_port, 
                           QN => n_1475);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n785, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_16_port, 
                           QN => n_1476);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n288, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_1_port, 
                           QN => n_1477);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n287, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_2_port, 
                           QN => n_1478);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n286, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_3_port, 
                           QN => n_1479);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n285, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_4_port, 
                           QN => n_1480);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n284, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_5_port, 
                           QN => n_1481);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n283, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_6_port, 
                           QN => n_1482);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n282, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_7_port, 
                           QN => n_1483);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n281, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_8_port, 
                           QN => n_1484);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n280, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_9_port, 
                           QN => n_1485);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n272, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_17_port, 
                           QN => n_1486);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n271, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_18_port, 
                           QN => n_1487);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n270, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_19_port, 
                           QN => n_1488);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n269, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_20_port, 
                           QN => n_1489);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n268, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_21_port, 
                           QN => n_1490);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n267, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_22_port, 
                           QN => n_1491);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n266, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_23_port, 
                           QN => n_1492);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n544, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_1_port, 
                           QN => n_1493);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n543, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_2_port, 
                           QN => n_1494);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n542, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_3_port, 
                           QN => n_1495);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n541, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_4_port, 
                           QN => n_1496);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n540, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_5_port, 
                           QN => n_1497);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n539, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_6_port, 
                           QN => n_1498);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n538, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_7_port, 
                           QN => n_1499);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n537, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_8_port, 
                           QN => n_1500);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n536, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_9_port, 
                           QN => n_1501);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n528, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_17_port, 
                           QN => n_1502);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n527, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_18_port, 
                           QN => n_1503);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n526, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_19_port, 
                           QN => n_1504);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n525, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_20_port, 
                           QN => n_1505);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n524, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_21_port, 
                           QN => n_1506);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n523, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_22_port, 
                           QN => n_1507);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n522, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_23_port, 
                           QN => n_1508);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n800, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_1_port, 
                           QN => n_1509);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n799, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_2_port, 
                           QN => n_1510);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n798, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_3_port, 
                           QN => n_1511);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n797, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_4_port, 
                           QN => n_1512);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n796, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_5_port, 
                           QN => n_1513);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n795, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_6_port, 
                           QN => n_1514);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n794, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_7_port, 
                           QN => n_1515);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n793, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_8_port, 
                           QN => n_1516);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n792, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_9_port, 
                           QN => n_1517);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n784, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_17_port, 
                           QN => n_1518);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n783, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_18_port, 
                           QN => n_1519);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n782, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_19_port, 
                           QN => n_1520);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n781, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_20_port, 
                           QN => n_1521);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n780, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_21_port, 
                           QN => n_1522);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n779, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_22_port, 
                           QN => n_1523);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n778, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_23_port, 
                           QN => n_1524);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n553, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_24_port, 
                           QN => n_1525);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n552, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_25_port, 
                           QN => n_1526);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n549, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_28_port, 
                           QN => n_1527);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_17_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n548, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_17_29_port, 
                           QN => n_1528);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n809, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_24_port, 
                           QN => n_1529);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n808, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_25_port, 
                           QN => n_1530);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n805, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_28_port, 
                           QN => n_1531);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_25_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n804, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_25_29_port, 
                           QN => n_1532);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n73, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_24_port, 
                           QN => n_1533);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n72, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_25_port, 
                           QN => n_1534);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n69, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_28_port, 
                           QN => n_1535);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_2_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n68, CK => 
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_2_29_port, 
                           QN => n_1536);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n105, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_24_port, 
                           QN => n_1537);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n104, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_25_port, 
                           QN => n_1538);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n101, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_28_port, 
                           QN => n_1539);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_3_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n100, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_3_29_port, 
                           QN => n_1540);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n361, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_24_port, 
                           QN => n_1541);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n360, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_25_port, 
                           QN => n_1542);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n357, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_28_port, 
                           QN => n_1543);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_11_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n356, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_11_29_port, 
                           QN => n_1544);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n841, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_24_port, 
                           QN => n_1545);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n840, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_25_port, 
                           QN => n_1546);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n837, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_28_port, 
                           QN => n_1547);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_26_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n836, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_26_29_port, 
                           QN => n_1548);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n873, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_24_port, 
                           QN => n_1549);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n872, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_25_port, 
                           QN => n_1550);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n869, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_28_port, 
                           QN => n_1551);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_27_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n868, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_27_29_port, 
                           QN => n_1552);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n263, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_26_port, 
                           QN => n_1553);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n262, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_27_port, 
                           QN => n_1554);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n259, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_30_port, 
                           QN => n_1555);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n258, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_31_port, 
                           QN => n_1556);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n519, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_26_port, 
                           QN => n_1557);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n518, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_27_port, 
                           QN => n_1558);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n515, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_30_port, 
                           QN => n_1559);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n514, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_31_port, 
                           QN => n_1560);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n775, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_26_port, 
                           QN => n_1561);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n774, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_27_port, 
                           QN => n_1562);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n771, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_30_port, 
                           QN => n_1563);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n770, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_31_port, 
                           QN => n_1564);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n265, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_24_port, 
                           QN => n_1565);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n264, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_25_port, 
                           QN => n_1566);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n261, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_28_port, 
                           QN => n_1567);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_8_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n260, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_8_29_port, 
                           QN => n_1568);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n521, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_24_port, 
                           QN => n_1569);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n520, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_25_port, 
                           QN => n_1570);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n517, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_28_port, 
                           QN => n_1571);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_16_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n516, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_16_29_port, 
                           QN => n_1572);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n777, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_24_port, 
                           QN => n_1573);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n776, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_25_port, 
                           QN => n_1574);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n773, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_28_port, 
                           QN => n_1575);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_24_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n772, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_24_29_port, 
                           QN => n_1576);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n417, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_0_port, 
                           QN => n_1577);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n407, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_10_port, 
                           QN => n_1578);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n406, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_11_port, 
                           QN => n_1579);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n405, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_12_port, 
                           QN => n_1580);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n404, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_13_port, 
                           QN => n_1581);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n403, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_14_port, 
                           QN => n_1582);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n402, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_15_port, 
                           QN => n_1583);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n401, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_16_port, 
                           QN => n_1584);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n416, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_1_port, 
                           QN => n_1585);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n415, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_2_port, 
                           QN => n_1586);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n414, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_3_port, 
                           QN => n_1587);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n413, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_4_port, 
                           QN => n_1588);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n412, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_5_port, 
                           QN => n_1589);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n411, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_6_port, 
                           QN => n_1590);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n410, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_7_port, 
                           QN => n_1591);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n409, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_8_port, 
                           QN => n_1592);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n408, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_9_port, 
                           QN => n_1593);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n400, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_17_port, 
                           QN => n_1594);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n399, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_18_port, 
                           QN => n_1595);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n398, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_19_port, 
                           QN => n_1596);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n397, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_20_port, 
                           QN => n_1597);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n396, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_21_port, 
                           QN => n_1598);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n395, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_22_port, 
                           QN => n_1599);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n394, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_23_port, 
                           QN => n_1600);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n929, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_0_port, 
                           QN => n_1601);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n919, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_10_port, 
                           QN => n_1602);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n918, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_11_port, 
                           QN => n_1603);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n917, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_12_port, 
                           QN => n_1604);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n916, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_13_port, 
                           QN => n_1605);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n915, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_14_port, 
                           QN => n_1606);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n914, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_15_port, 
                           QN => n_1607);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n913, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_16_port, 
                           QN => n_1608);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n928, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_1_port, 
                           QN => n_1609);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n927, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_2_port, 
                           QN => n_1610);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n926, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_3_port, 
                           QN => n_1611);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n925, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_4_port, 
                           QN => n_1612);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n924, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_5_port, 
                           QN => n_1613);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n923, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_6_port, 
                           QN => n_1614);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n922, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_7_port, 
                           QN => n_1615);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n921, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_8_port, 
                           QN => n_1616);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n920, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_9_port, 
                           QN => n_1617);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n912, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_17_port, 
                           QN => n_1618);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n911, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_18_port, 
                           QN => n_1619);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n910, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_19_port, 
                           QN => n_1620);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n909, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_20_port, 
                           QN => n_1621);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n908, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_21_port, 
                           QN => n_1622);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n907, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_22_port, 
                           QN => n_1623);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n906, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_23_port, 
                           QN => n_1624);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n673, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_0_port, 
                           QN => n_1625);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n663, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_10_port, 
                           QN => n_1626);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n662, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_11_port, 
                           QN => n_1627);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n661, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_12_port, 
                           QN => n_1628);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n660, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_13_port, 
                           QN => n_1629);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n659, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_14_port, 
                           QN => n_1630);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n658, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_15_port, 
                           QN => n_1631);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n657, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_16_port, 
                           QN => n_1632);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n705, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_0_port, 
                           QN => n_1633);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n695, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_10_port, 
                           QN => n_1634);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n694, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_11_port, 
                           QN => n_1635);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n693, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_12_port, 
                           QN => n_1636);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n692, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_13_port, 
                           QN => n_1637);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n691, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_14_port, 
                           QN => n_1638);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n690, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_15_port, 
                           QN => n_1639);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n689, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_16_port, 
                           QN => n_1640);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n672, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_1_port, 
                           QN => n_1641);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n671, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_2_port, 
                           QN => n_1642);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n670, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_3_port, 
                           QN => n_1643);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n669, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_4_port, 
                           QN => n_1644);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n668, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_5_port, 
                           QN => n_1645);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n667, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_6_port, 
                           QN => n_1646);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n666, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_7_port, 
                           QN => n_1647);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n665, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_8_port, 
                           QN => n_1648);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n664, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_9_port, 
                           QN => n_1649);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n656, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_17_port, 
                           QN => n_1650);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n655, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_18_port, 
                           QN => n_1651);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n654, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_19_port, 
                           QN => n_1652);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n653, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_20_port, 
                           QN => n_1653);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n652, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_21_port, 
                           QN => n_1654);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n651, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_22_port, 
                           QN => n_1655);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n650, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_23_port, 
                           QN => n_1656);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n704, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_1_port, 
                           QN => n_1657);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n703, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_2_port, 
                           QN => n_1658);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n702, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_3_port, 
                           QN => n_1659);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n701, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_4_port, 
                           QN => n_1660);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n700, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_5_port, 
                           QN => n_1661);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n699, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_6_port, 
                           QN => n_1662);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n698, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_7_port, 
                           QN => n_1663);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n697, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_8_port, 
                           QN => n_1664);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n696, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_9_port, 
                           QN => n_1665);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n688, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_17_port, 
                           QN => n_1666);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n687, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_18_port, 
                           QN => n_1667);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n686, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_19_port, 
                           QN => n_1668);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n685, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_20_port, 
                           QN => n_1669);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n684, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_21_port, 
                           QN => n_1670);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n683, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_22_port, 
                           QN => n_1671);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n682, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_23_port, 
                           QN => n_1672);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n225, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_0_port, 
                           QN => n_1673);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n215, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_10_port, 
                           QN => n_1674);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n214, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_11_port, 
                           QN => n_1675);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n213, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_12_port, 
                           QN => n_1676);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n212, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_13_port, 
                           QN => n_1677);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n211, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_14_port, 
                           QN => n_1678);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n210, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_15_port, 
                           QN => n_1679);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n209, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_16_port, 
                           QN => n_1680);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n224, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_1_port, 
                           QN => n_1681);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n223, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_2_port, 
                           QN => n_1682);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n222, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_3_port, 
                           QN => n_1683);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n221, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_4_port, 
                           QN => n_1684);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n220, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_5_port, 
                           QN => n_1685);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n219, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_6_port, 
                           QN => n_1686);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n218, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_7_port, 
                           QN => n_1687);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n217, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_8_port, 
                           QN => n_1688);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n216, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_9_port, 
                           QN => n_1689);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n208, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_17_port, 
                           QN => n_1690);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n207, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_18_port, 
                           QN => n_1691);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n206, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_19_port, 
                           QN => n_1692);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n205, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_20_port, 
                           QN => n_1693);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n204, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_21_port, 
                           QN => n_1694);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n203, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_22_port, 
                           QN => n_1695);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n202, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_23_port, 
                           QN => n_1696);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n257, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_0_port, 
                           QN => n_1697);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n247, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_10_port, 
                           QN => n_1698);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n246, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_11_port, 
                           QN => n_1699);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n245, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_12_port, 
                           QN => n_1700);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n244, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_13_port, 
                           QN => n_1701);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n243, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_14_port, 
                           QN => n_1702);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n242, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_15_port, 
                           QN => n_1703);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n241, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_16_port, 
                           QN => n_1704);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n256, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_1_port, 
                           QN => n_1705);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n255, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_2_port, 
                           QN => n_1706);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n254, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_3_port, 
                           QN => n_1707);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n253, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_4_port, 
                           QN => n_1708);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n252, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_5_port, 
                           QN => n_1709);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n251, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_6_port, 
                           QN => n_1710);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n250, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_7_port, 
                           QN => n_1711);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n249, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_8_port, 
                           QN => n_1712);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n248, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_9_port, 
                           QN => n_1713);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n240, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_17_port, 
                           QN => n_1714);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n239, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_18_port, 
                           QN => n_1715);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n238, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_19_port, 
                           QN => n_1716);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n237, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_20_port, 
                           QN => n_1717);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n236, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_21_port, 
                           QN => n_1718);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n235, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_22_port, 
                           QN => n_1719);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n234, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_23_port, 
                           QN => n_1720);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n391, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_26_port, 
                           QN => n_1721);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n390, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_27_port, 
                           QN => n_1722);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n387, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_30_port, 
                           QN => n_1723);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n386, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_31_port, 
                           QN => n_1724);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n903, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_26_port, 
                           QN => n_1725);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n902, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_27_port, 
                           QN => n_1726);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n899, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_30_port, 
                           QN => n_1727);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n898, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_31_port, 
                           QN => n_1728);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n647, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_26_port, 
                           QN => n_1729);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n646, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_27_port, 
                           QN => n_1730);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n643, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_30_port, 
                           QN => n_1731);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n642, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_31_port, 
                           QN => n_1732);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n679, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_26_port, 
                           QN => n_1733);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n678, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_27_port, 
                           QN => n_1734);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n675, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_30_port, 
                           QN => n_1735);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n674, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_31_port, 
                           QN => n_1736);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n199, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_26_port, 
                           QN => n_1737);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n198, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_27_port, 
                           QN => n_1738);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n195, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_30_port, 
                           QN => n_1739);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n194, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_31_port, 
                           QN => n_1740);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n231, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_26_port, 
                           QN => n_1741);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n230, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_27_port, 
                           QN => n_1742);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n227, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_30_port, 
                           QN => n_1743);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n226, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_31_port, 
                           QN => n_1744);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n393, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_24_port, 
                           QN => n_1745);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n392, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_25_port, 
                           QN => n_1746);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n389, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_28_port, 
                           QN => n_1747);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_12_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n388, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_12_29_port, 
                           QN => n_1748);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n905, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_24_port, 
                           QN => n_1749);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n904, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_25_port, 
                           QN => n_1750);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n901, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_28_port, 
                           QN => n_1751);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_28_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n900, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_28_29_port, 
                           QN => n_1752);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n649, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_24_port, 
                           QN => n_1753);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n648, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_25_port, 
                           QN => n_1754);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n645, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_28_port, 
                           QN => n_1755);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_20_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n644, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_20_29_port, 
                           QN => n_1756);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n681, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_24_port, 
                           QN => n_1757);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n680, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_25_port, 
                           QN => n_1758);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n677, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_28_port, 
                           QN => n_1759);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_21_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n676, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_21_29_port, 
                           QN => n_1760);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n201, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_24_port, 
                           QN => n_1761);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n200, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_25_port, 
                           QN => n_1762);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n197, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_28_port, 
                           QN => n_1763);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_6_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n196, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_6_29_port, 
                           QN => n_1764);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n233, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_24_port, 
                           QN => n_1765);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n232, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_25_port, 
                           QN => n_1766);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n229, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_28_port, 
                           QN => n_1767);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_7_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n228, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_7_29_port, 
                           QN => n_1768);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n513, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_0_port, 
                           QN => n_1769);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n503, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_10_port, 
                           QN => n_1770);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n502, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_11_port, 
                           QN => n_1771);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n501, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_12_port, 
                           QN => n_1772);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n500, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_13_port, 
                           QN => n_1773);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n499, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_14_port, 
                           QN => n_1774);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n498, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_15_port, 
                           QN => n_1775);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n497, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_16_port, 
                           QN => n_1776);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n512, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_1_port, 
                           QN => n_1777);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n511, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_2_port, 
                           QN => n_1778);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n510, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_3_port, 
                           QN => n_1779);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n509, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_4_port, 
                           QN => n_1780);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n508, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_5_port, 
                           QN => n_1781);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n507, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_6_port, 
                           QN => n_1782);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n506, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_7_port, 
                           QN => n_1783);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n505, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_8_port, 
                           QN => n_1784);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n504, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_9_port, 
                           QN => n_1785);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n496, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_17_port, 
                           QN => n_1786);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n495, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_18_port, 
                           QN => n_1787);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n494, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_19_port, 
                           QN => n_1788);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n493, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_20_port, 
                           QN => n_1789);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n492, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_21_port, 
                           QN => n_1790);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n491, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_22_port, 
                           QN => n_1791);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n490, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_23_port, 
                           QN => n_1792);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n487, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_26_port, 
                           QN => n_1793);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n486, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_27_port, 
                           QN => n_1794);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n483, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_30_port, 
                           QN => n_1795);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n482, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_31_port, 
                           QN => n_1796);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n489, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_24_port, 
                           QN => n_1797);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n488, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_25_port, 
                           QN => n_1798);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n485, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_28_port, 
                           QN => n_1799);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_15_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n484, CK =>
                           CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_15_29_port, 
                           QN => n_1800);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3508, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1801, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n346);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3406, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1802, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n608);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3407, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1803, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n607);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3408, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1804, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n606);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3409, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1805, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n605);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3410, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1806, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n604);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3411, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1807, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n603);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3412, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1808, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n602);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3374, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1809, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n640);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3375, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1810, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n639);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3376, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1811, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n638);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3377, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1812, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n637);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3378, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1813, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n636);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3379, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1814, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n635);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3380, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1815, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n634);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3207, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1816, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1031);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3208, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1817, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1030);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3211, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1818, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1027);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3212, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1819, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1026);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3191, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1820, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1047);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3192, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1821, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1046);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3193, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1822, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1045);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3194, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1823, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1044);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3195, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1824, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1043);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3196, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1825, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1042);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3197, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1826, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1041);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3189, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1827, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1049);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3190, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1828, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1048);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3198, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1829, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1040);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3199, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1830, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1039);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3200, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1831, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1038);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3201, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1832, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1037);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3202, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1833, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1036);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3203, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1834, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1035);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3204, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1835, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1034);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3205, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1836, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1033);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3206, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1837, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1032);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3209, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1838, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1029);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3210, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1839, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1028);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3687, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1840, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n7);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3688, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1841, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n6);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3691, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1842, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3692, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1843, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n2);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3671, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1844, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n23);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3672, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1845, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n22);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3673, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1846, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n21);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3674, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1847, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n20);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3675, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1848, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n19);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3676, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1849, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n18);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3677, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1850, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n17);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3669, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1851, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n25);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3670, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1852, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n24);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3678, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1853, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n16);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3679, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1854, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n15);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3680, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1855, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n14);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3681, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1856, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n13);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3682, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1857, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n12);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3683, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1858, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n11);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3684, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1859, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n10);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3685, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1860, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n9);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3686, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1861, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n8);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3689, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1862, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n5);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3690, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1863, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3181, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1864, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1057);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3182, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1865, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1056);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3183, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1866, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1055);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3184, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1867, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1054);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3185, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1868, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1053);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3186, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1869, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1052);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3187, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1870, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1051);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_32_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3188, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1871, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1050);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3661, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1872, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n33);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3662, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1873, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n32);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3663, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1874, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n31);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3664, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1875, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n30);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3665, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1876, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n29);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3666, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1877, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n28);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3667, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1878, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n27);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_0_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3668, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1879, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n26);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3367, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1880, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n711);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3368, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1881, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n710);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3371, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1882, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n707);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3372, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1883, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n706);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3335, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1884, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n743);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3336, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1885, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n742);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3339, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1886, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n739);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3340, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1887, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n738);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3351, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1888, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n727);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3352, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1889, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n726);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3353, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1890, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n725);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3354, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1891, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n724);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3355, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1892, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n723);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3356, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1893, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n722);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3357, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1894, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n721);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3319, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1895, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n759);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3320, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1896, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n758);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3321, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1897, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n757);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3322, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1898, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n756);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3323, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1899, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n755);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3324, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1900, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n754);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3325, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1901, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n753);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3349, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1902, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n729);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3350, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1903, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n728);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3358, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1904, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n720);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3359, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1905, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n719);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3360, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1906, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n718);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3361, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1907, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n717);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3362, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1908, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n716);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3363, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1909, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n715);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3364, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1910, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n714);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3365, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1911, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n713);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3366, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1912, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n712);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3369, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1913, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n709);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3370, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1914, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n708);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3317, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1915, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n761);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3318, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1916, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n760);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3326, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1917, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n752);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3327, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1918, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n751);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3328, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1919, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n750);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3329, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1920, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n749);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3330, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1921, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n748);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3331, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1922, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n747);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3332, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1923, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n746);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3333, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1924, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n745);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3334, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1925, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n744);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3337, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1926, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n741);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3338, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1927, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n740);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3463, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1928, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n455);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3464, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1929, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n454);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3467, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1930, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n451);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3468, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1931, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n450);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3623, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1932, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n135);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3624, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1933, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n134);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3627, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1934, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n131);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3628, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1935, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n130);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3591, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1936, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n167);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3592, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1937, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n166);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3595, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1938, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n163);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3596, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1939, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n162);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3495, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1940, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n423);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3496, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1941, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n422);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3499, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1942, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n419);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3500, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1943, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n418);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3271, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1944, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n967);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3272, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1945, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n966);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3275, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1946, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n963);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3276, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1947, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n962);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3303, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1948, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n935);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3304, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1949, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n934);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3307, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1950, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n931);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3308, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1951, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n930);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3447, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1952, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n471);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3448, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1953, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n470);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3449, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1954, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n469);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3450, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1955, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n468);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3451, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1956, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n467);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3452, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1957, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n466);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3453, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1958, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n465);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3445, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1959, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n473);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3446, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1960, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n472);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3454, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1961, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n464);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3455, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1962, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n463);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3456, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1963, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n462);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3457, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1964, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n461);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3458, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1965, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n460);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3459, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1966, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n459);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3460, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1967, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n458);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3461, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1968, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n457);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3462, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1969, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n456);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3465, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1970, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n453);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3466, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1971, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n452);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3607, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1972, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n151);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3608, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1973, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n150);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3609, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1974, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n149);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3610, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1975, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n148);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3611, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1976, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n147);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3612, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1977, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n146);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3613, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1978, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n145);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3575, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1979, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n183);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3576, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1980, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n182);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3577, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1981, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n181);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3578, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1982, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n180);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3579, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1983, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n179);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3580, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1984, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n178);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3581, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1985, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n177);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3479, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1986, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n439);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3480, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1987, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n438);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3481, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1988, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n437);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3482, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1989, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n436);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3483, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1990, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n435);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3484, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1991, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n434);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3485, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1992, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n433);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3605, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1993, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n153);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3606, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1994, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n152);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3614, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1995, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n144);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3615, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1996, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n143);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3616, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1997, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n142);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3617, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1998, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n141);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3618, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_1999, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n140);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3619, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2000, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n139);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3620, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2001, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n138);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3621, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2002, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n137);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3622, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2003, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n136);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3625, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2004, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n133);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3626, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2005, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n132);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3573, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2006, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n185);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3574, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2007, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n184);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3582, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2008, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n176);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3583, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2009, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n175);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3584, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2010, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n174);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3585, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2011, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n173);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3586, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2012, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n172);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3587, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2013, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n171);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3588, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2014, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n170);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3589, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2015, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n169);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3590, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2016, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n168);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3593, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2017, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n165);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3594, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2018, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n164);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3477, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2019, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n441);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3478, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2020, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n440);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3486, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2021, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n432);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3487, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2022, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n431);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3488, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2023, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n430);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3489, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2024, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n429);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3490, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2025, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n428);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3491, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2026, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n427);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3492, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2027, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n426);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3493, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2028, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n425);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3494, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2029, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n424);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3497, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2030, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n421);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3498, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2031, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n420);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3255, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2032, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n983);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3256, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2033, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n982);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3257, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2034, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n981);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3258, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2035, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n980);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3259, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2036, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n979);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3260, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2037, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n978);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3261, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2038, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n977);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3253, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2039, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n985);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3254, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2040, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n984);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3262, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2041, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n976);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3263, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2042, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n975);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3264, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2043, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n974);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3265, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2044, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n973);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3266, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2045, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n972);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3267, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2046, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n971);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3268, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2047, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n970);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3269, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2048, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n969);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3270, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2049, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n968);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3273, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2050, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n965);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3274, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2051, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n964);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3287, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2052, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n951);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3288, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2053, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n950);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3289, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2054, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n949);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3290, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2055, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n948);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3291, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2056, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n947);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3292, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2057, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n946);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3293, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2058, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n945);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3285, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2059, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n953);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3286, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2060, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n952);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3294, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2061, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n944);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3295, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2062, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n943);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3296, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2063, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n942);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3297, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2064, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n941);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3298, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2065, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n940);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3299, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2066, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n939);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3300, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2067, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n938);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3301, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2068, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n937);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3302, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2069, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n936);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3305, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2070, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n933);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3306, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2071, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n932);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3341, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2072, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n737);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3309, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2073, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n769);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3342, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2074, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n736);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3343, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2075, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n735);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3344, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2076, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n734);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3345, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2077, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n733);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3346, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2078, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n732);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3347, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2079, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n731);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_22_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3348, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2080, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n730);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3310, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2081, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n768);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3311, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2082, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n767);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3312, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2083, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n766);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3313, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2084, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n765);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3314, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2085, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n764);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3315, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2086, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n763);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_23_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3316, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2087, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n762);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3437, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2088, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n481);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3438, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2089, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n480);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3439, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2090, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n479);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3440, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2091, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n478);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3441, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2092, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n477);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3442, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2093, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n476);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3443, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2094, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n475);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_14_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3444, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2095, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n474);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3597, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2096, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n161);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3565, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2097, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n193);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3469, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2098, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n449);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3598, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2099, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n160);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3599, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2100, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n159);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3600, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2101, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n158);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3601, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2102, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n157);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3602, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2103, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n156);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3603, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2104, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n155);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_4_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3604, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2105, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n154);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3566, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2106, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n192);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3567, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2107, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n191);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3568, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2108, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n190);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3569, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2109, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n189);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3570, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2110, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n188);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3571, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2111, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n187);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_5_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3572, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2112, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n186);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3470, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2113, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n448);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3471, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2114, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n447);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3472, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2115, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n446);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3473, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2116, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n445);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3474, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2117, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n444);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3475, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2118, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n443);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_13_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3476, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2119, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n442);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3245, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2120, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n993);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3246, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2121, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n992);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3247, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2122, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n991);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3248, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2123, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n990);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3249, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2124, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n989);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3250, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2125, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n988);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3251, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2126, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n987);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_30_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3252, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2127, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n986);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3277, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2128, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n961);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3278, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2129, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n960);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3279, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2130, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n959);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3280, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2131, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n958);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3281, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2132, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n957);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3282, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2133, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n956);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3283, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2134, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n955);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_29_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3284, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2135, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n954);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3239, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2136, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n999);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3240, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2137, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n998);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3243, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2138, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n995);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3244, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2139, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n994);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3223, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2140, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1015);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3224, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2141, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1014);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3225, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2142, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1013);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3226, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2143, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1012);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3227, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2144, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1011);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3228, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2145, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1010);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3229, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2146, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1009);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3221, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2147, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1017);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3222, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2148, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1016);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3230, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2149, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1008);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3231, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2150, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1007);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3232, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2151, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1006);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3233, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2152, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1005);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3234, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2153, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1004);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3235, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2154, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1003);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3236, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2155, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1002);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3237, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2156, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1001);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3238, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2157, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1000);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3241, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2158, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n997);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3242, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2159, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n996);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3213, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2160, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1025);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3214, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2161, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1024);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3215, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2162, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1023);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3216, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2163, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1022);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3217, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2164, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1021);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3218, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2165, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1020);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3219, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2166, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1019);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_31_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3220, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n4237, Q =>
                           n_2167, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1018);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_0_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N359_port, 
                           Q => dp_id_stage_out1_i_0_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_0_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N427_port, 
                           Q => dp_id_stage_out2_i_0_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_1_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N358_port, 
                           Q => dp_id_stage_out1_i_1_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_1_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N426_port, 
                           Q => dp_id_stage_out2_i_1_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_2_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N357_port, 
                           Q => dp_id_stage_out1_i_2_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_2_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N425_port, 
                           Q => dp_id_stage_out2_i_2_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_3_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N356_port, 
                           Q => dp_id_stage_out1_i_3_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_3_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N424_port, 
                           Q => dp_id_stage_out2_i_3_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_4_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N355_port, 
                           Q => dp_id_stage_out1_i_4_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_4_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N423_port, 
                           Q => dp_id_stage_out2_i_4_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_5_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N354_port, 
                           Q => dp_id_stage_out1_i_5_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_5_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N422_port, 
                           Q => dp_id_stage_out2_i_5_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_6_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N353_port, 
                           Q => dp_id_stage_out1_i_6_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_6_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N421_port, 
                           Q => dp_id_stage_out2_i_6_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_7_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N352_port, 
                           Q => dp_id_stage_out1_i_7_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_7_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N420_port, 
                           Q => dp_id_stage_out2_i_7_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_8_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N351_port, 
                           Q => dp_id_stage_out1_i_8_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_8_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N419_port, 
                           Q => dp_id_stage_out2_i_8_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_9_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4233,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N350_port, 
                           Q => dp_id_stage_out1_i_9_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_9_inst : DLH_X1 port map( 
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4230,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N418_port, 
                           Q => dp_id_stage_out2_i_9_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_10_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N349_port, 
                           Q => dp_id_stage_out1_i_10_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_10_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N417_port, 
                           Q => dp_id_stage_out2_i_10_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_11_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N348_port, 
                           Q => dp_id_stage_out1_i_11_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_11_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N416_port, 
                           Q => dp_id_stage_out2_i_11_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_12_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N347_port, 
                           Q => dp_id_stage_out1_i_12_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_12_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N415_port, 
                           Q => dp_id_stage_out2_i_12_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_13_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N346_port, 
                           Q => dp_id_stage_out1_i_13_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_13_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N414_port, 
                           Q => dp_id_stage_out2_i_13_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_14_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N345_port, 
                           Q => dp_id_stage_out1_i_14_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_14_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N413_port, 
                           Q => dp_id_stage_out2_i_14_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_15_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N344_port, 
                           Q => dp_id_stage_out1_i_15_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_15_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N412_port, 
                           Q => dp_id_stage_out2_i_15_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_16_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N343_port, 
                           Q => dp_id_stage_out1_i_16_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_16_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N411_port, 
                           Q => dp_id_stage_out2_i_16_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_17_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N342_port, 
                           Q => dp_id_stage_out1_i_17_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_17_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N410_port, 
                           Q => dp_id_stage_out2_i_17_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_18_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N341_port, 
                           Q => dp_id_stage_out1_i_18_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_18_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N409_port, 
                           Q => dp_id_stage_out2_i_18_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_19_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N340_port, 
                           Q => dp_id_stage_out1_i_19_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_19_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N408_port, 
                           Q => dp_id_stage_out2_i_19_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_20_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4232,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N339_port, 
                           Q => dp_id_stage_out1_i_20_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_20_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4229,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N407_port, 
                           Q => dp_id_stage_out2_i_20_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_21_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N338_port, 
                           Q => dp_id_stage_out1_i_21_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_21_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N406_port, 
                           Q => dp_id_stage_out2_i_21_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_22_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N337_port, 
                           Q => dp_id_stage_out1_i_22_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_22_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N405_port, 
                           Q => dp_id_stage_out2_i_22_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_23_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N336_port, 
                           Q => dp_id_stage_out1_i_23_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_23_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N404_port, 
                           Q => dp_id_stage_out2_i_23_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_24_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N335_port, 
                           Q => dp_id_stage_out1_i_24_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_24_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N403_port, 
                           Q => dp_id_stage_out2_i_24_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_25_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N334_port, 
                           Q => dp_id_stage_out1_i_25_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_25_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N402_port, 
                           Q => dp_id_stage_out2_i_25_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_26_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N333_port, 
                           Q => dp_id_stage_out1_i_26_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_26_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N401_port, 
                           Q => dp_id_stage_out2_i_26_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_27_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N332_port, 
                           Q => dp_id_stage_out1_i_27_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_27_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N400_port, 
                           Q => dp_id_stage_out2_i_27_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_28_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N331_port, 
                           Q => dp_id_stage_out1_i_28_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_28_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N399_port, 
                           Q => dp_id_stage_out2_i_28_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_29_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N330_port, 
                           Q => dp_id_stage_out1_i_29_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_29_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N398_port, 
                           Q => dp_id_stage_out2_i_29_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_30_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N329_port, 
                           Q => dp_id_stage_out1_i_30_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_30_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N397_port, 
                           Q => dp_id_stage_out2_i_30_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT1_reg_31_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4231,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N328_port, 
                           Q => dp_id_stage_out1_i_31_port);
   dp_id_stage_regfile_DataPath_Physical_RF_OUT2_reg_31_inst : DLH_X1 port map(
                           G => dp_id_stage_regfile_DataPath_Physical_RF_n4228,
                           D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_N396_port, 
                           Q => dp_id_stage_out2_i_31_port);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3373, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1171, Q =>
                           n_2168, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n641);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3381, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174, Q =>
                           n_2169, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n633);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3382, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174, Q =>
                           n_2170, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n632);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3383, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174, Q =>
                           n_2171, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n631);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3384, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174, Q =>
                           n_2172, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n630);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3385, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174, Q =>
                           n_2173, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n629);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3386, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174, Q =>
                           n_2174, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n628);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3387, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174, Q =>
                           n_2175, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n627);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3388, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1174, Q =>
                           n_2176, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n626);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3389, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2177, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n625);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3390, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2178, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n624);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3391, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2179, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n623);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3392, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2180, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n622);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3393, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2181, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n621);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3394, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2182, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n620);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3395, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2183, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n619);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3396, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2184, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n618);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3397, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2185, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n617);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3398, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2186, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n616);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3399, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2187, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n615);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3400, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1175, Q =>
                           n_2188, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n614);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3401, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1176, Q =>
                           n_2189, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n613);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3402, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1176, Q =>
                           n_2190, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n612);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3403, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1176, Q =>
                           n_2191, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n611);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_19_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3404, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1176, Q =>
                           n_2192, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n610);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3405, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1176, Q =>
                           n_2193, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n609);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3413, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2194, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n601);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3414, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2195, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n600);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3415, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2196, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n599);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3416, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2197, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n598);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3417, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2198, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n597);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3418, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2199, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n596);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3419, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2200, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n595);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3420, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2201, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n594);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3421, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2202, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n593);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3422, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2203, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n592);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3423, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2204, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n591);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3424, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1177, Q =>
                           n_2205, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n590);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3425, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2206, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n589);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3426, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2207, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n588);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3427, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2208, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n587);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3428, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2209, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n586);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3429, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2210, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n585);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3430, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2211, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n584);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3431, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2212, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n583);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3432, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2213, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n582);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3433, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2214, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n581);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3434, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2215, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n580);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3435, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2216, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n579);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_18_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3436, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1178, Q =>
                           n_2217, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n578);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3501, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1179, Q =>
                           n_2218, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n353);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3502, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1179, Q =>
                           n_2219, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n352);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3503, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1179, Q =>
                           n_2220, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n351);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3504, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1179, Q =>
                           n_2221, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n350);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3505, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2222, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n349);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3506, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2223, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n348);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3507, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2224, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n347);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3509, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2225, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n345);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3510, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2226, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n344);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3511, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2227, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n343);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3512, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2228, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n342);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3513, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2229, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n341);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3514, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2230, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n340);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3515, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2231, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n339);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3516, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1180, Q =>
                           n_2232, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n338);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3517, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2233, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n337);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3518, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2234, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n336);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3519, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2235, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n335);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3520, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2236, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n334);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3521, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2237, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n333);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3522, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2238, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n332);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3523, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2239, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n331);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3524, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2240, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n330);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3525, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2241, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n329);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3526, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2242, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n328);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3527, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2243, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n327);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3528, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1181, Q =>
                           n_2244, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n326);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3529, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2245, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n325);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3530, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2246, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n324);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3531, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2247, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n323);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_10_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3532, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2248, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n322);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3533, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2249, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n321);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3534, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2250, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n320);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3535, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2251, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n319);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3536, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2252, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n318);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3537, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2253, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n317);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3538, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2254, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n316);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3539, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2255, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n315);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3540, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1182, Q =>
                           n_2256, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n314);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3541, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2257, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n313);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3542, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2258, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n312);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3543, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2259, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n311);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3544, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2260, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n310);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3545, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2261, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n309);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3546, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2262, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n308);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3547, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2263, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n307);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3548, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2264, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n306);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3549, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2265, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n305);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3550, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2266, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n304);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3551, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2267, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n303);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3552, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1183, Q =>
                           n_2268, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n302);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3553, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2269, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n301);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3554, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2270, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n300);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3555, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2271, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n299);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3556, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2272, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n298);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3557, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2273, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n297);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3558, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2274, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n296);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3559, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2275, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n295);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3560, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2276, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n294);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3561, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2277, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n293);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3562, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2278, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n292);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3563, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2279, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n291);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_9_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3564, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1184, Q =>
                           n_2280, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n290);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_0_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3629, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1185, Q =>
                           n_2281, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n65);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_1_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3630, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1185, Q =>
                           n_2282, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n64);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_2_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3631, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1185, Q =>
                           n_2283, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n63);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_3_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3632, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1185, Q =>
                           n_2284, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n62);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_4_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3633, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2285, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n61);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_5_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3634, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2286, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n60);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_6_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3635, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2287, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n59);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_7_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3636, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2288, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n58);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_8_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3637, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2289, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n57);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_9_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3638, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2290, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n56);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_10_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3639, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2291, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n55);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_11_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3640, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2292, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n54);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_12_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3641, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2293, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n53);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_13_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3642, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2294, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n52);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_14_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3643, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2295, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n51);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_15_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3644, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1186, Q =>
                           n_2296, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n50);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_16_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3645, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2297, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n49);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_17_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3646, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2298, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n48);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_18_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3647, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2299, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n47);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_19_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3648, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2300, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n46);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_20_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3649, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2301, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n45);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_21_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3650, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2302, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n44);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_22_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3651, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2303, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n43);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_23_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3652, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2304, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n42);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_24_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3653, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2305, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n41);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_25_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3654, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2306, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n40);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_26_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3655, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2307, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n39);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_27_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3656, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1187, Q =>
                           n_2308, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n38);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_28_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3657, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1188, Q =>
                           n_2309, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n37);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_29_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3658, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1188, Q =>
                           n_2310, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n36);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_30_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3659, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1188, Q =>
                           n_2311, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n35);
   dp_id_stage_regfile_DataPath_Physical_RF_REGISTERS_reg_1_31_inst : DFFR_X1 
                           port map( D => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n3660, CK 
                           => CLK, RN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n1188, Q =>
                           n_2312, QN => 
                           dp_id_stage_regfile_DataPath_Physical_RF_n34);
   dp_ex_stage_U11 : NOR4_X1 port map( A1 => dp_rf_out1_ex_i_1_port, A2 => 
                           dp_rf_out1_ex_i_19_port, A3 => 
                           dp_rf_out1_ex_i_18_port, A4 => 
                           dp_rf_out1_ex_i_17_port, ZN => dp_ex_stage_n5);
   dp_ex_stage_U10 : NOR4_X1 port map( A1 => dp_rf_out1_ex_i_16_port, A2 => 
                           dp_rf_out1_ex_i_15_port, A3 => 
                           dp_rf_out1_ex_i_14_port, A4 => 
                           dp_rf_out1_ex_i_13_port, ZN => dp_ex_stage_n4);
   dp_ex_stage_U9 : NOR4_X1 port map( A1 => dp_rf_out1_ex_i_12_port, A2 => 
                           dp_rf_out1_ex_i_11_port, A3 => 
                           dp_rf_out1_ex_i_10_port, A4 => 
                           dp_rf_out1_ex_i_0_port, ZN => dp_ex_stage_n3);
   dp_ex_stage_U8 : NAND4_X1 port map( A1 => dp_ex_stage_n3, A2 => 
                           dp_ex_stage_n4, A3 => dp_ex_stage_n5, A4 => 
                           dp_ex_stage_n6, ZN => dp_ex_stage_n2);
   dp_ex_stage_U7 : NAND4_X1 port map( A1 => dp_ex_stage_n7, A2 => 
                           dp_ex_stage_n8, A3 => dp_ex_stage_n9, A4 => 
                           dp_ex_stage_n10, ZN => dp_ex_stage_n1);
   dp_ex_stage_U6 : OR2_X1 port map( A1 => dp_ex_stage_n1, A2 => dp_ex_stage_n2
                           , ZN => dp_branch_t_ex_o);
   dp_ex_stage_U5 : NOR4_X1 port map( A1 => dp_rf_out1_ex_i_27_port, A2 => 
                           dp_rf_out1_ex_i_26_port, A3 => 
                           dp_rf_out1_ex_i_25_port, A4 => 
                           dp_rf_out1_ex_i_24_port, ZN => dp_ex_stage_n7);
   dp_ex_stage_U4 : NOR4_X1 port map( A1 => dp_rf_out1_ex_i_30_port, A2 => 
                           dp_rf_out1_ex_i_2_port, A3 => 
                           dp_rf_out1_ex_i_29_port, A4 => 
                           dp_rf_out1_ex_i_28_port, ZN => dp_ex_stage_n8);
   dp_ex_stage_U3 : NOR4_X1 port map( A1 => dp_rf_out1_ex_i_5_port, A2 => 
                           dp_rf_out1_ex_i_4_port, A3 => dp_rf_out1_ex_i_3_port
                           , A4 => dp_rf_out1_ex_i_31_port, ZN => 
                           dp_ex_stage_n9);
   dp_ex_stage_U2 : NOR4_X1 port map( A1 => dp_rf_out1_ex_i_9_port, A2 => 
                           dp_rf_out1_ex_i_8_port, A3 => dp_rf_out1_ex_i_7_port
                           , A4 => dp_rf_out1_ex_i_6_port, ZN => 
                           dp_ex_stage_n10);
   dp_ex_stage_U1 : NOR4_X1 port map( A1 => dp_rf_out1_ex_i_23_port, A2 => 
                           dp_rf_out1_ex_i_22_port, A3 => 
                           dp_rf_out1_ex_i_21_port, A4 => 
                           dp_rf_out1_ex_i_20_port, ZN => dp_ex_stage_n6);
   dp_ex_stage_muxA_U40 : MUX2_X1 port map( A => dp_rf_out1_ex_i_31_port, B => 
                           dp_npc_ex_i_31_port, S => dp_ex_stage_muxA_n2, Z => 
                           dp_ex_stage_muxA_out_31_port);
   dp_ex_stage_muxA_U39 : MUX2_X1 port map( A => dp_rf_out1_ex_i_30_port, B => 
                           dp_npc_ex_i_30_port, S => dp_ex_stage_muxA_n3, Z => 
                           dp_ex_stage_muxA_out_30_port);
   dp_ex_stage_muxA_U38 : MUX2_X1 port map( A => dp_rf_out1_ex_i_29_port, B => 
                           dp_npc_ex_i_29_port, S => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_out_29_port);
   dp_ex_stage_muxA_U37 : MUX2_X1 port map( A => dp_rf_out1_ex_i_28_port, B => 
                           dp_npc_ex_i_28_port, S => dp_ex_stage_muxA_n2, Z => 
                           dp_ex_stage_muxA_out_28_port);
   dp_ex_stage_muxA_U36 : MUX2_X1 port map( A => dp_rf_out1_ex_i_27_port, B => 
                           dp_npc_ex_i_27_port, S => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_out_27_port);
   dp_ex_stage_muxA_U35 : MUX2_X1 port map( A => dp_rf_out1_ex_i_26_port, B => 
                           dp_npc_ex_i_26_port, S => dp_ex_stage_muxA_n3, Z => 
                           dp_ex_stage_muxA_out_26_port);
   dp_ex_stage_muxA_U34 : MUX2_X1 port map( A => dp_rf_out1_ex_i_25_port, B => 
                           dp_npc_ex_i_25_port, S => dp_ex_stage_muxA_n3, Z => 
                           dp_ex_stage_muxA_out_25_port);
   dp_ex_stage_muxA_U33 : MUX2_X1 port map( A => dp_rf_out1_ex_i_24_port, B => 
                           dp_npc_ex_i_24_port, S => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_out_24_port);
   dp_ex_stage_muxA_U32 : MUX2_X1 port map( A => dp_rf_out1_ex_i_23_port, B => 
                           dp_npc_ex_i_23_port, S => dp_ex_stage_muxA_n6, Z => 
                           dp_ex_stage_muxA_out_23_port);
   dp_ex_stage_muxA_U31 : MUX2_X1 port map( A => dp_rf_out1_ex_i_22_port, B => 
                           dp_npc_ex_i_22_port, S => dp_ex_stage_muxA_n6, Z => 
                           dp_ex_stage_muxA_out_22_port);
   dp_ex_stage_muxA_U30 : MUX2_X1 port map( A => dp_rf_out1_ex_i_21_port, B => 
                           dp_npc_ex_i_21_port, S => dp_ex_stage_muxA_n8, Z => 
                           dp_ex_stage_muxA_out_21_port);
   dp_ex_stage_muxA_U29 : MUX2_X1 port map( A => dp_rf_out1_ex_i_20_port, B => 
                           dp_npc_ex_i_20_port, S => dp_ex_stage_muxA_n6, Z => 
                           dp_ex_stage_muxA_out_20_port);
   dp_ex_stage_muxA_U28 : MUX2_X1 port map( A => dp_rf_out1_ex_i_18_port, B => 
                           dp_npc_ex_i_18_port, S => dp_ex_stage_muxA_n5, Z => 
                           dp_ex_stage_muxA_n27);
   dp_ex_stage_muxA_U27 : MUX2_X1 port map( A => dp_rf_out1_ex_i_17_port, B => 
                           dp_npc_ex_i_17_port, S => dp_ex_stage_muxA_n8, Z => 
                           dp_ex_stage_muxA_out_17_port);
   dp_ex_stage_muxA_U26 : MUX2_X1 port map( A => dp_rf_out1_ex_i_16_port, B => 
                           dp_npc_ex_i_16_port, S => dp_ex_stage_muxA_n4, Z => 
                           dp_ex_stage_muxA_out_16_port);
   dp_ex_stage_muxA_U25 : MUX2_X1 port map( A => dp_rf_out1_ex_i_15_port, B => 
                           dp_npc_ex_i_15_port, S => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_out_15_port);
   dp_ex_stage_muxA_U24 : MUX2_X1 port map( A => dp_rf_out1_ex_i_13_port, B => 
                           dp_npc_ex_i_13_port, S => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_out_13_port);
   dp_ex_stage_muxA_U23 : MUX2_X1 port map( A => dp_rf_out1_ex_i_10_port, B => 
                           dp_npc_ex_i_10_port, S => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_out_10_port);
   dp_ex_stage_muxA_U22 : MUX2_X1 port map( A => dp_rf_out1_ex_i_9_port, B => 
                           dp_npc_ex_i_9_port, S => dp_ex_stage_muxA_n6, Z => 
                           dp_ex_stage_muxA_out_9_port);
   dp_ex_stage_muxA_U21 : MUX2_X1 port map( A => dp_rf_out1_ex_i_8_port, B => 
                           dp_npc_ex_i_8_port, S => dp_ex_stage_muxA_n8, Z => 
                           dp_ex_stage_muxA_out_8_port);
   dp_ex_stage_muxA_U20 : MUX2_X1 port map( A => dp_rf_out1_ex_i_7_port, B => 
                           dp_npc_ex_i_7_port, S => dp_ex_stage_muxA_n6, Z => 
                           dp_ex_stage_muxA_out_7_port);
   dp_ex_stage_muxA_U19 : MUX2_X1 port map( A => dp_rf_out1_ex_i_6_port, B => 
                           dp_npc_ex_i_6_port, S => dp_ex_stage_muxA_n8, Z => 
                           dp_ex_stage_muxA_out_6_port);
   dp_ex_stage_muxA_U18 : MUX2_X1 port map( A => dp_rf_out1_ex_i_5_port, B => 
                           dp_npc_ex_i_5_port, S => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_out_5_port);
   dp_ex_stage_muxA_U17 : MUX2_X1 port map( A => dp_rf_out1_ex_i_4_port, B => 
                           dp_npc_ex_i_4_port, S => dp_ex_stage_muxA_n5, Z => 
                           dp_ex_stage_muxA_out_4_port);
   dp_ex_stage_muxA_U16 : MUX2_X1 port map( A => dp_rf_out1_ex_i_3_port, B => 
                           dp_npc_ex_i_3_port, S => dp_ex_stage_muxA_n8, Z => 
                           dp_ex_stage_muxA_out_3_port);
   dp_ex_stage_muxA_U15 : MUX2_X1 port map( A => dp_rf_out1_ex_i_1_port, B => 
                           dp_npc_ex_i_1_port, S => dp_ex_stage_muxA_n3, Z => 
                           dp_ex_stage_muxA_out_1_port);
   dp_ex_stage_muxA_U14 : MUX2_X1 port map( A => dp_rf_out1_ex_i_0_port, B => 
                           dp_npc_ex_i_0_port, S => dp_ex_stage_muxA_n8, Z => 
                           dp_ex_stage_muxA_out_0_port);
   dp_ex_stage_muxA_U13 : CLKBUF_X3 port map( A => muxA_sel_i, Z => 
                           dp_ex_stage_muxA_n7);
   dp_ex_stage_muxA_U12 : CLKBUF_X1 port map( A => muxA_sel_i, Z => 
                           dp_ex_stage_muxA_n6);
   dp_ex_stage_muxA_U11 : MUX2_X1 port map( A => dp_rf_out1_ex_i_2_port, B => 
                           dp_npc_ex_i_2_port, S => dp_ex_stage_muxA_n8, Z => 
                           dp_ex_stage_muxA_out_2_port);
   dp_ex_stage_muxA_U10 : BUF_X1 port map( A => muxA_sel_i, Z => 
                           dp_ex_stage_muxA_n5);
   dp_ex_stage_muxA_U9 : CLKBUF_X1 port map( A => muxA_sel_i, Z => 
                           dp_ex_stage_muxA_n3);
   dp_ex_stage_muxA_U8 : MUX2_X1 port map( A => dp_rf_out1_ex_i_11_port, B => 
                           dp_npc_ex_i_11_port, S => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_out_11_port);
   dp_ex_stage_muxA_U7 : MUX2_X1 port map( A => dp_rf_out1_ex_i_12_port, B => 
                           dp_npc_ex_i_12_port, S => dp_ex_stage_muxA_n3, Z => 
                           dp_ex_stage_muxA_out_12_port);
   dp_ex_stage_muxA_U6 : BUF_X1 port map( A => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_n2);
   dp_ex_stage_muxA_U5 : CLKBUF_X3 port map( A => muxA_sel_i, Z => 
                           dp_ex_stage_muxA_n8);
   dp_ex_stage_muxA_U4 : BUF_X1 port map( A => dp_ex_stage_muxA_n7, Z => 
                           dp_ex_stage_muxA_n4);
   dp_ex_stage_muxA_U3 : MUX2_X1 port map( A => dp_rf_out1_ex_i_14_port, B => 
                           dp_npc_ex_i_14_port, S => dp_ex_stage_muxA_n5, Z => 
                           dp_ex_stage_muxA_out_14_port);
   dp_ex_stage_muxA_U2 : BUF_X2 port map( A => dp_ex_stage_muxA_n27, Z => 
                           dp_ex_stage_muxA_out_18_port);
   dp_ex_stage_muxA_U1 : MUX2_X1 port map( A => dp_rf_out1_ex_i_19_port, B => 
                           dp_npc_ex_i_19_port, S => dp_ex_stage_muxA_n8, Z => 
                           dp_ex_stage_muxA_out_19_port);
   dp_ex_stage_muxB_U40 : MUX2_X1 port map( A => dp_data_mem_ex_o_31_port, B =>
                           dp_imm_ex_i_31_port, S => dp_ex_stage_muxB_n8, Z => 
                           dp_ex_stage_muxB_out_31_port);
   dp_ex_stage_muxB_U39 : MUX2_X1 port map( A => dp_data_mem_ex_o_30_port, B =>
                           dp_imm_ex_i_30_port, S => dp_ex_stage_muxB_n8, Z => 
                           dp_ex_stage_muxB_out_30_port);
   dp_ex_stage_muxB_U38 : MUX2_X1 port map( A => dp_data_mem_ex_o_29_port, B =>
                           dp_imm_ex_i_29_port, S => dp_ex_stage_muxB_n8, Z => 
                           dp_ex_stage_muxB_out_29_port);
   dp_ex_stage_muxB_U37 : MUX2_X1 port map( A => dp_data_mem_ex_o_28_port, B =>
                           dp_imm_ex_i_28_port, S => dp_ex_stage_muxB_n8, Z => 
                           dp_ex_stage_muxB_out_28_port);
   dp_ex_stage_muxB_U36 : MUX2_X1 port map( A => dp_data_mem_ex_o_27_port, B =>
                           dp_imm_ex_i_27_port, S => dp_ex_stage_muxB_n8, Z => 
                           dp_ex_stage_muxB_out_27_port);
   dp_ex_stage_muxB_U35 : MUX2_X1 port map( A => dp_data_mem_ex_o_26_port, B =>
                           dp_imm_ex_i_26_port, S => dp_ex_stage_muxB_n8, Z => 
                           dp_ex_stage_muxB_out_26_port);
   dp_ex_stage_muxB_U34 : MUX2_X1 port map( A => dp_data_mem_ex_o_25_port, B =>
                           dp_imm_ex_i_25_port, S => dp_ex_stage_muxB_n8, Z => 
                           dp_ex_stage_muxB_out_25_port);
   dp_ex_stage_muxB_U33 : MUX2_X1 port map( A => dp_data_mem_ex_o_24_port, B =>
                           dp_imm_ex_i_24_port, S => dp_ex_stage_muxB_n8, Z => 
                           dp_ex_stage_muxB_out_24_port);
   dp_ex_stage_muxB_U32 : MUX2_X1 port map( A => dp_data_mem_ex_o_23_port, B =>
                           dp_imm_ex_i_23_port, S => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_out_23_port);
   dp_ex_stage_muxB_U31 : MUX2_X1 port map( A => dp_data_mem_ex_o_22_port, B =>
                           dp_imm_ex_i_22_port, S => dp_ex_stage_muxB_n3, Z => 
                           dp_ex_stage_muxB_out_22_port);
   dp_ex_stage_muxB_U30 : MUX2_X1 port map( A => dp_data_mem_ex_o_21_port, B =>
                           dp_imm_ex_i_21_port, S => dp_ex_stage_muxB_n3, Z => 
                           dp_ex_stage_muxB_out_21_port);
   dp_ex_stage_muxB_U29 : MUX2_X1 port map( A => dp_data_mem_ex_o_20_port, B =>
                           dp_imm_ex_i_20_port, S => dp_ex_stage_muxB_n4, Z => 
                           dp_ex_stage_muxB_out_20_port);
   dp_ex_stage_muxB_U28 : MUX2_X1 port map( A => dp_data_mem_ex_o_19_port, B =>
                           dp_imm_ex_i_19_port, S => dp_ex_stage_muxB_n3, Z => 
                           dp_ex_stage_muxB_out_19_port);
   dp_ex_stage_muxB_U27 : MUX2_X1 port map( A => dp_data_mem_ex_o_18_port, B =>
                           dp_imm_ex_i_18_port, S => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_out_18_port);
   dp_ex_stage_muxB_U26 : MUX2_X1 port map( A => dp_data_mem_ex_o_17_port, B =>
                           dp_imm_ex_i_17_port, S => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_out_17_port);
   dp_ex_stage_muxB_U25 : MUX2_X1 port map( A => dp_data_mem_ex_o_16_port, B =>
                           dp_imm_ex_i_16_port, S => dp_ex_stage_muxB_n3, Z => 
                           dp_ex_stage_muxB_out_16_port);
   dp_ex_stage_muxB_U24 : MUX2_X1 port map( A => dp_data_mem_ex_o_15_port, B =>
                           dp_imm_ex_i_15_port, S => dp_ex_stage_muxB_n2, Z => 
                           dp_ex_stage_muxB_out_15_port);
   dp_ex_stage_muxB_U23 : MUX2_X1 port map( A => dp_data_mem_ex_o_14_port, B =>
                           dp_imm_ex_i_14_port, S => dp_ex_stage_muxB_n1, Z => 
                           dp_ex_stage_muxB_out_14_port);
   dp_ex_stage_muxB_U22 : MUX2_X1 port map( A => dp_data_mem_ex_o_13_port, B =>
                           dp_imm_ex_i_13_port, S => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_out_13_port);
   dp_ex_stage_muxB_U21 : MUX2_X1 port map( A => dp_data_mem_ex_o_12_port, B =>
                           dp_imm_ex_i_12_port, S => dp_ex_stage_muxB_n3, Z => 
                           dp_ex_stage_muxB_out_12_port);
   dp_ex_stage_muxB_U20 : MUX2_X1 port map( A => dp_data_mem_ex_o_11_port, B =>
                           dp_imm_ex_i_11_port, S => dp_ex_stage_muxB_n3, Z => 
                           dp_ex_stage_muxB_out_11_port);
   dp_ex_stage_muxB_U19 : MUX2_X1 port map( A => dp_data_mem_ex_o_10_port, B =>
                           dp_imm_ex_i_10_port, S => dp_ex_stage_muxB_n5, Z => 
                           dp_ex_stage_muxB_out_10_port);
   dp_ex_stage_muxB_U18 : MUX2_X1 port map( A => dp_data_mem_ex_o_9_port, B => 
                           dp_imm_ex_i_9_port, S => dp_ex_stage_muxB_n3, Z => 
                           dp_ex_stage_muxB_out_9_port);
   dp_ex_stage_muxB_U17 : MUX2_X1 port map( A => dp_data_mem_ex_o_8_port, B => 
                           dp_imm_ex_i_8_port, S => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_out_8_port);
   dp_ex_stage_muxB_U16 : MUX2_X1 port map( A => dp_data_mem_ex_o_7_port, B => 
                           dp_imm_ex_i_7_port, S => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_out_7_port);
   dp_ex_stage_muxB_U15 : MUX2_X1 port map( A => dp_data_mem_ex_o_6_port, B => 
                           dp_imm_ex_i_6_port, S => dp_ex_stage_muxB_n5, Z => 
                           dp_ex_stage_muxB_out_6_port);
   dp_ex_stage_muxB_U14 : MUX2_X1 port map( A => dp_data_mem_ex_o_5_port, B => 
                           dp_imm_ex_i_5_port, S => dp_ex_stage_muxB_n2, Z => 
                           dp_ex_stage_muxB_out_5_port);
   dp_ex_stage_muxB_U13 : MUX2_X1 port map( A => dp_data_mem_ex_o_4_port, B => 
                           dp_imm_ex_i_4_port, S => dp_ex_stage_muxB_n5, Z => 
                           dp_ex_stage_muxB_out_4_port);
   dp_ex_stage_muxB_U12 : MUX2_X1 port map( A => dp_data_mem_ex_o_3_port, B => 
                           dp_imm_ex_i_3_port, S => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_out_3_port);
   dp_ex_stage_muxB_U11 : MUX2_X1 port map( A => dp_data_mem_ex_o_2_port, B => 
                           dp_imm_ex_i_2_port, S => dp_ex_stage_muxB_n5, Z => 
                           dp_ex_stage_muxB_out_2_port);
   dp_ex_stage_muxB_U10 : MUX2_X1 port map( A => dp_data_mem_ex_o_1_port, B => 
                           dp_imm_ex_i_1_port, S => muxB_sel_i, Z => 
                           dp_ex_stage_muxB_out_1_port);
   dp_ex_stage_muxB_U9 : MUX2_X1 port map( A => dp_data_mem_ex_o_0_port, B => 
                           dp_imm_ex_i_0_port, S => muxB_sel_i, Z => 
                           dp_ex_stage_muxB_out_0_port);
   dp_ex_stage_muxB_U8 : CLKBUF_X1 port map( A => muxB_sel_i, Z => 
                           dp_ex_stage_muxB_n5);
   dp_ex_stage_muxB_U7 : CLKBUF_X1 port map( A => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_n4);
   dp_ex_stage_muxB_U6 : CLKBUF_X3 port map( A => muxB_sel_i, Z => 
                           dp_ex_stage_muxB_n7);
   dp_ex_stage_muxB_U5 : BUF_X1 port map( A => muxB_sel_i, Z => 
                           dp_ex_stage_muxB_n6);
   dp_ex_stage_muxB_U4 : BUF_X2 port map( A => dp_ex_stage_muxB_n6, Z => 
                           dp_ex_stage_muxB_n3);
   dp_ex_stage_muxB_U3 : CLKBUF_X1 port map( A => dp_ex_stage_muxB_n6, Z => 
                           dp_ex_stage_muxB_n2);
   dp_ex_stage_muxB_U2 : CLKBUF_X2 port map( A => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_n8);
   dp_ex_stage_muxB_U1 : CLKBUF_X1 port map( A => dp_ex_stage_muxB_n7, Z => 
                           dp_ex_stage_muxB_n1);
   dp_ex_stage_alu_U347 : OAI211_X1 port map( C1 => dp_ex_stage_alu_n268, C2 =>
                           dp_ex_stage_alu_n267, A => dp_ex_stage_alu_n266, B 
                           => dp_ex_stage_alu_n265, ZN => 
                           dp_alu_out_ex_o_0_port);
   dp_ex_stage_alu_U346 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n263, B2 => 
                           dp_ex_stage_alu_n189, A => dp_ex_stage_alu_n262, ZN 
                           => dp_ex_stage_alu_n264);
   dp_ex_stage_alu_U345 : INV_X1 port map( A => dp_ex_stage_alu_n21, ZN => 
                           dp_ex_stage_alu_n262);
   dp_ex_stage_alu_U344 : MUX2_X1 port map( A => dp_ex_stage_alu_n190, B => 
                           dp_ex_stage_alu_n188, S => dp_ex_stage_alu_n45, Z =>
                           dp_ex_stage_alu_n263);
   dp_ex_stage_alu_U343 : MUX2_X1 port map( A => dp_ex_stage_alu_n258, B => 
                           dp_ex_stage_alu_n257, S => dp_ex_stage_alu_n191, Z 
                           => dp_ex_stage_alu_n259);
   dp_ex_stage_alu_U342 : AND2_X1 port map( A1 => dp_ex_stage_alu_N20_port, A2 
                           => dp_ex_stage_alu_n26, ZN => dp_ex_stage_alu_n255);
   dp_ex_stage_alu_U341 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n254, A2 => 
                           dp_ex_stage_alu_n26, ZN => dp_ex_stage_alu_n258);
   dp_ex_stage_alu_U340 : MUX2_X1 port map( A => dp_ex_stage_alu_N17_port, B =>
                           dp_ex_stage_alu_N18_port, S => dp_ex_stage_alu_n93, 
                           Z => dp_ex_stage_alu_n254);
   dp_ex_stage_alu_U339 : OAI21_X1 port map( B1 => dp_ex_stage_alu_n21, B2 => 
                           dp_ex_stage_alu_n190, A => dp_ex_stage_alu_n189, ZN 
                           => dp_ex_stage_alu_n261);
   dp_ex_stage_alu_U338 : MUX2_X1 port map( A => dp_ex_stage_alu_n253, B => 
                           dp_ex_stage_alu_n252, S => dp_ex_stage_alu_n2, Z => 
                           dp_ex_stage_alu_n268);
   dp_ex_stage_alu_U337 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n251, A2 => 
                           dp_ex_stage_alu_n51, ZN => dp_ex_stage_alu_n252);
   dp_ex_stage_alu_U336 : INV_X1 port map( A => alu_op_i_1_port, ZN => 
                           dp_ex_stage_alu_n271);
   dp_ex_stage_alu_U335 : MUX2_X1 port map( A => dp_ex_stage_alu_N22_port, B =>
                           dp_ex_stage_alu_N21_port, S => alu_op_i_0_port, Z =>
                           dp_ex_stage_alu_n251);
   dp_ex_stage_alu_U334 : NAND2_X1 port map( A1 => dp_ex_stage_alu_N16_port, A2
                           => dp_ex_stage_alu_n24, ZN => dp_ex_stage_alu_n253);
   dp_ex_stage_alu_U333 : NAND3_X1 port map( A1 => dp_ex_stage_alu_n206, A2 => 
                           dp_ex_stage_alu_n40, A3 => dp_ex_stage_alu_n250, ZN 
                           => dp_ex_stage_alu_n97);
   dp_ex_stage_alu_U332 : OAI21_X1 port map( B1 => dp_ex_stage_alu_n24, B2 => 
                           dp_ex_stage_alu_n267, A => alu_op_i_4_port, ZN => 
                           dp_ex_stage_alu_n250);
   dp_ex_stage_alu_U331 : NAND3_X1 port map( A1 => dp_ex_stage_alu_n205, A2 => 
                           dp_ex_stage_alu_n191, A3 => dp_ex_stage_alu_n61, ZN 
                           => dp_ex_stage_alu_n190);
   dp_ex_stage_alu_U330 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n205, A2 => 
                           dp_ex_stage_alu_n54, ZN => dp_ex_stage_alu_n188);
   dp_ex_stage_alu_U329 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n66, A2 => 
                           dp_ex_stage_alu_n269, ZN => dp_ex_stage_alu_n189);
   dp_ex_stage_alu_U328 : INV_X1 port map( A => alu_op_i_4_port, ZN => 
                           dp_ex_stage_alu_n269);
   dp_ex_stage_alu_U327 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n270, A2 => 
                           dp_ex_stage_alu_n311, ZN => dp_ex_stage_alu_n267);
   dp_ex_stage_alu_U326 : INV_X2 port map( A => dp_ex_stage_alu_n241, ZN => 
                           dp_ex_stage_alu_n240);
   dp_ex_stage_alu_U325 : INV_X1 port map( A => dp_ex_stage_alu_n223, ZN => 
                           dp_ex_stage_alu_n222);
   dp_ex_stage_alu_U324 : CLKBUF_X1 port map( A => dp_ex_stage_alu_n310, Z => 
                           dp_ex_stage_alu_n215);
   dp_ex_stage_alu_U323 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_31_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_31_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n118);
   dp_ex_stage_alu_U322 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_20_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_20_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n154);
   dp_ex_stage_alu_U321 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_27_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_27_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n133);
   dp_ex_stage_alu_U320 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_23_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_23_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n145);
   dp_ex_stage_alu_U319 : NAND4_X1 port map( A1 => dp_ex_stage_alu_n272, A2 => 
                           dp_ex_stage_alu_n271, A3 => dp_ex_stage_alu_n270, A4
                           => dp_ex_stage_alu_n27, ZN => dp_ex_stage_alu_n90);
   dp_ex_stage_alu_U318 : NOR3_X1 port map( A1 => dp_ex_stage_alu_n93, A2 => 
                           alu_op_i_4_port, A3 => dp_ex_stage_alu_n272, ZN => 
                           dp_ex_stage_alu_n205);
   dp_ex_stage_alu_U317 : INV_X1 port map( A => alu_op_i_3_port, ZN => 
                           dp_ex_stage_alu_n311);
   dp_ex_stage_alu_U316 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n212, B2 => 
                           dp_ex_stage_alu_n219, A => dp_ex_stage_alu_n201, ZN 
                           => dp_ex_stage_alu_n155);
   dp_ex_stage_alu_U315 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_26_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_26_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n136);
   dp_ex_stage_alu_U314 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_25_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_25_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n139);
   dp_ex_stage_alu_U313 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_21_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_21_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n151);
   dp_ex_stage_alu_U312 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_12_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_12_port, B2 => 
                           dp_ex_stage_alu_n218, ZN => dp_ex_stage_alu_n181);
   dp_ex_stage_alu_U311 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n179, B2 =>
                           dp_ex_stage_alu_n230, C1 => dp_ex_stage_alu_n180, C2
                           => dp_ex_stage_alu_n288, A => dp_ex_stage_alu_n181, 
                           ZN => dp_alu_out_ex_o_12_port);
   dp_ex_stage_alu_U310 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_29_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_29_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n127);
   dp_ex_stage_alu_U309 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_28_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_28_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n130);
   dp_ex_stage_alu_U308 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_22_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_22_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n148);
   dp_ex_stage_alu_U307 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_30_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_30_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n121);
   dp_ex_stage_alu_U306 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_24_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_24_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n142);
   dp_ex_stage_alu_U305 : INV_X1 port map( A => dp_ex_stage_muxB_out_20_port, 
                           ZN => dp_ex_stage_alu_n296);
   dp_ex_stage_alu_U304 : INV_X1 port map( A => dp_ex_stage_muxA_out_20_port, 
                           ZN => dp_ex_stage_alu_n278);
   dp_ex_stage_alu_U303 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n296, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n152);
   dp_ex_stage_alu_U302 : OR2_X1 port map( A1 => dp_ex_stage_alu_n153, A2 => 
                           dp_ex_stage_alu_n296, ZN => dp_ex_stage_alu_n193);
   dp_ex_stage_alu_U301 : OR2_X1 port map( A1 => dp_ex_stage_alu_n152, A2 => 
                           dp_ex_stage_alu_n278, ZN => dp_ex_stage_alu_n192);
   dp_ex_stage_alu_U300 : INV_X1 port map( A => dp_ex_stage_alu_n311, ZN => 
                           dp_ex_stage_alu_n191);
   dp_ex_stage_alu_U299 : CLKBUF_X1 port map( A => alu_op_i_1_port, Z => 
                           dp_ex_stage_alu_n93);
   dp_ex_stage_alu_U298 : INV_X1 port map( A => dp_ex_stage_muxB_out_23_port, 
                           ZN => dp_ex_stage_alu_n299);
   dp_ex_stage_alu_U297 : INV_X1 port map( A => dp_ex_stage_muxA_out_23_port, 
                           ZN => dp_ex_stage_alu_n242);
   dp_ex_stage_alu_U296 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n299, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n143);
   dp_ex_stage_alu_U295 : OR2_X1 port map( A1 => dp_ex_stage_alu_n144, A2 => 
                           dp_ex_stage_alu_n299, ZN => dp_ex_stage_alu_n92);
   dp_ex_stage_alu_U294 : OR2_X1 port map( A1 => dp_ex_stage_alu_n143, A2 => 
                           dp_ex_stage_alu_n242, ZN => dp_ex_stage_alu_n89);
   dp_ex_stage_alu_U293 : INV_X1 port map( A => dp_ex_stage_muxB_out_27_port, 
                           ZN => dp_ex_stage_alu_n303);
   dp_ex_stage_alu_U292 : INV_X1 port map( A => dp_ex_stage_muxA_out_27_port, 
                           ZN => dp_ex_stage_alu_n246);
   dp_ex_stage_alu_U291 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n303, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n131);
   dp_ex_stage_alu_U290 : OR2_X1 port map( A1 => dp_ex_stage_alu_n132, A2 => 
                           dp_ex_stage_alu_n303, ZN => dp_ex_stage_alu_n88);
   dp_ex_stage_alu_U289 : OR2_X1 port map( A1 => dp_ex_stage_alu_n131, A2 => 
                           dp_ex_stage_alu_n246, ZN => dp_ex_stage_alu_n87);
   dp_ex_stage_alu_U288 : INV_X1 port map( A => dp_ex_stage_muxB_out_26_port, 
                           ZN => dp_ex_stage_alu_n302);
   dp_ex_stage_alu_U287 : INV_X1 port map( A => dp_ex_stage_muxA_out_26_port, 
                           ZN => dp_ex_stage_alu_n245);
   dp_ex_stage_alu_U286 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n302, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n134);
   dp_ex_stage_alu_U285 : OR2_X1 port map( A1 => dp_ex_stage_alu_n135, A2 => 
                           dp_ex_stage_alu_n302, ZN => dp_ex_stage_alu_n86);
   dp_ex_stage_alu_U284 : OR2_X1 port map( A1 => dp_ex_stage_alu_n134, A2 => 
                           dp_ex_stage_alu_n245, ZN => dp_ex_stage_alu_n85);
   dp_ex_stage_alu_U283 : INV_X1 port map( A => dp_ex_stage_muxB_out_25_port, 
                           ZN => dp_ex_stage_alu_n301);
   dp_ex_stage_alu_U282 : INV_X1 port map( A => dp_ex_stage_muxA_out_25_port, 
                           ZN => dp_ex_stage_alu_n244);
   dp_ex_stage_alu_U281 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n301, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n137);
   dp_ex_stage_alu_U280 : OR2_X1 port map( A1 => dp_ex_stage_alu_n138, A2 => 
                           dp_ex_stage_alu_n301, ZN => dp_ex_stage_alu_n84);
   dp_ex_stage_alu_U279 : OR2_X1 port map( A1 => dp_ex_stage_alu_n137, A2 => 
                           dp_ex_stage_alu_n244, ZN => dp_ex_stage_alu_n83);
   dp_ex_stage_alu_U278 : INV_X1 port map( A => dp_ex_stage_muxB_out_22_port, 
                           ZN => dp_ex_stage_alu_n298);
   dp_ex_stage_alu_U277 : INV_X1 port map( A => dp_ex_stage_muxA_out_22_port, 
                           ZN => dp_ex_stage_alu_n241);
   dp_ex_stage_alu_U276 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n212, B2 => 
                           dp_ex_stage_alu_n298, A => dp_ex_stage_alu_n201, ZN 
                           => dp_ex_stage_alu_n146);
   dp_ex_stage_alu_U275 : OR2_X1 port map( A1 => dp_ex_stage_alu_n147, A2 => 
                           dp_ex_stage_alu_n298, ZN => dp_ex_stage_alu_n82);
   dp_ex_stage_alu_U274 : OR2_X1 port map( A1 => dp_ex_stage_alu_n146, A2 => 
                           dp_ex_stage_alu_n39, ZN => dp_ex_stage_alu_n81);
   dp_ex_stage_alu_U273 : INV_X1 port map( A => dp_ex_stage_muxB_out_21_port, 
                           ZN => dp_ex_stage_alu_n297);
   dp_ex_stage_alu_U272 : INV_X1 port map( A => dp_ex_stage_muxA_out_21_port, 
                           ZN => dp_ex_stage_alu_n239);
   dp_ex_stage_alu_U271 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n212, B2 => 
                           dp_ex_stage_alu_n297, A => dp_ex_stage_alu_n201, ZN 
                           => dp_ex_stage_alu_n149);
   dp_ex_stage_alu_U270 : OR2_X1 port map( A1 => dp_ex_stage_alu_n150, A2 => 
                           dp_ex_stage_alu_n297, ZN => dp_ex_stage_alu_n80);
   dp_ex_stage_alu_U269 : OR2_X1 port map( A1 => dp_ex_stage_alu_n149, A2 => 
                           dp_ex_stage_alu_n239, ZN => dp_ex_stage_alu_n79);
   dp_ex_stage_alu_U268 : INV_X1 port map( A => dp_ex_stage_alu_n71, ZN => 
                           dp_ex_stage_alu_n226);
   dp_ex_stage_alu_U267 : INV_X1 port map( A => dp_ex_stage_alu_n34, ZN => 
                           dp_ex_stage_alu_n225);
   dp_ex_stage_alu_U266 : INV_X1 port map( A => dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_n221);
   dp_ex_stage_alu_U265 : INV_X1 port map( A => dp_ex_stage_alu_n52, ZN => 
                           dp_ex_stage_alu_n274);
   dp_ex_stage_alu_U264 : INV_X1 port map( A => dp_ex_stage_alu_n74, ZN => 
                           dp_ex_stage_alu_n228);
   dp_ex_stage_alu_U263 : INV_X1 port map( A => dp_ex_stage_alu_n69, ZN => 
                           dp_ex_stage_alu_n224);
   dp_ex_stage_alu_U262 : INV_X1 port map( A => dp_ex_stage_alu_n72, ZN => 
                           dp_ex_stage_alu_n227);
   dp_ex_stage_alu_U261 : INV_X1 port map( A => dp_ex_stage_alu_n50, ZN => 
                           dp_ex_stage_alu_n220);
   dp_ex_stage_alu_U260 : INV_X1 port map( A => dp_ex_stage_alu_n29, ZN => 
                           dp_ex_stage_alu_n234);
   dp_ex_stage_alu_U259 : INV_X1 port map( A => dp_ex_stage_muxA_out_16_port, 
                           ZN => dp_ex_stage_alu_n235);
   dp_ex_stage_alu_U258 : INV_X1 port map( A => dp_ex_stage_muxB_out_1_port, ZN
                           => dp_ex_stage_alu_n219);
   dp_ex_stage_alu_U257 : INV_X1 port map( A => dp_ex_stage_alu_n33, ZN => 
                           dp_ex_stage_alu_n229);
   dp_ex_stage_alu_U256 : INV_X1 port map( A => dp_ex_stage_muxA_out_14_port, 
                           ZN => dp_ex_stage_alu_n233);
   dp_ex_stage_alu_U255 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n110, B2 =>
                           dp_ex_stage_alu_n274, C1 => dp_ex_stage_alu_n111, C2
                           => dp_ex_stage_alu_n223, A => dp_ex_stage_alu_n112, 
                           ZN => dp_alu_out_ex_o_4_port);
   dp_ex_stage_alu_U254 : INV_X1 port map( A => dp_ex_stage_muxA_out_18_port, 
                           ZN => dp_ex_stage_alu_n237);
   dp_ex_stage_alu_U253 : INV_X1 port map( A => dp_ex_stage_alu_n78, ZN => 
                           dp_ex_stage_alu_n276);
   dp_ex_stage_alu_U252 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n104, B2 =>
                           dp_ex_stage_alu_n276, C1 => dp_ex_stage_alu_n105, C2
                           => dp_ex_stage_alu_n282, A => dp_ex_stage_alu_n106, 
                           ZN => dp_alu_out_ex_o_6_port);
   dp_ex_stage_alu_U251 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n107, B2 =>
                           dp_ex_stage_alu_n275, C1 => dp_ex_stage_alu_n108, C2
                           => dp_ex_stage_alu_n281, A => dp_ex_stage_alu_n109, 
                           ZN => dp_alu_out_ex_o_5_port);
   dp_ex_stage_alu_U250 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n113, B2 =>
                           dp_ex_stage_alu_n224, C1 => dp_ex_stage_alu_n114, C2
                           => dp_ex_stage_alu_n221, A => dp_ex_stage_alu_n115, 
                           ZN => dp_alu_out_ex_o_3_port);
   dp_ex_stage_alu_U249 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n164, B2 =>
                           dp_ex_stage_alu_n236, C1 => dp_ex_stage_alu_n165, C2
                           => dp_ex_stage_alu_n293, A => dp_ex_stage_alu_n166, 
                           ZN => dp_alu_out_ex_o_17_port);
   dp_ex_stage_alu_U248 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n212, B2 => 
                           dp_ex_stage_alu_n300, A => dp_ex_stage_alu_n201, ZN 
                           => dp_ex_stage_alu_n140);
   dp_ex_stage_alu_U247 : NAND2_X1 port map( A1 => alu_op_i_4_port, A2 => 
                           dp_ex_stage_alu_n66, ZN => 
                           dp_ex_stage_alu_shift_arith_i);
   dp_ex_stage_alu_U246 : INV_X1 port map( A => dp_ex_stage_muxB_out_4_port, ZN
                           => dp_ex_stage_alu_n223);
   dp_ex_stage_alu_U245 : INV_X1 port map( A => dp_ex_stage_muxA_out_17_port, 
                           ZN => dp_ex_stage_alu_n236);
   dp_ex_stage_alu_U244 : INV_X1 port map( A => dp_ex_stage_alu_n32, ZN => 
                           dp_ex_stage_alu_n230);
   dp_ex_stage_alu_U243 : INV_X1 port map( A => dp_ex_stage_muxA_out_24_port, 
                           ZN => dp_ex_stage_alu_n243);
   dp_ex_stage_alu_U242 : INV_X1 port map( A => dp_ex_stage_muxA_out_31_port, 
                           ZN => dp_ex_stage_alu_n249);
   dp_ex_stage_alu_U241 : INV_X1 port map( A => dp_ex_stage_muxA_out_28_port, 
                           ZN => dp_ex_stage_alu_n248);
   dp_ex_stage_alu_U240 : INV_X1 port map( A => alu_op_i_2_port, ZN => 
                           dp_ex_stage_alu_n270);
   dp_ex_stage_alu_U239 : INV_X1 port map( A => dp_ex_stage_muxA_out_13_port, 
                           ZN => dp_ex_stage_alu_n232);
   dp_ex_stage_alu_U238 : AND4_X1 port map( A1 => alu_op_i_2_port, A2 => 
                           alu_op_i_0_port, A3 => dp_ex_stage_alu_n311, A4 => 
                           dp_ex_stage_alu_n269, ZN => dp_ex_stage_alu_n68);
   dp_ex_stage_alu_U237 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n295, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n158);
   dp_ex_stage_alu_U236 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n283, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n101);
   dp_ex_stage_alu_U234 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n101, B2 =>
                           dp_ex_stage_alu_n225, C1 => dp_ex_stage_alu_n102, C2
                           => dp_ex_stage_alu_n283, A => dp_ex_stage_alu_n103, 
                           ZN => dp_alu_out_ex_o_7_port);
   dp_ex_stage_alu_U233 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n212, B2 => 
                           dp_ex_stage_alu_n294, A => dp_ex_stage_alu_n201, ZN 
                           => dp_ex_stage_alu_n161);
   dp_ex_stage_alu_U232 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n289, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n176);
   dp_ex_stage_alu_U231 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n176, B2 =>
                           dp_ex_stage_alu_n232, C1 => dp_ex_stage_alu_n177, C2
                           => dp_ex_stage_alu_n289, A => dp_ex_stage_alu_n178, 
                           ZN => dp_alu_out_ex_o_13_port);
   dp_ex_stage_alu_U229 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n290, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n173);
   dp_ex_stage_alu_U228 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n173, B2 =>
                           dp_ex_stage_alu_n233, C1 => dp_ex_stage_alu_n174, C2
                           => dp_ex_stage_alu_n290, A => dp_ex_stage_alu_n175, 
                           ZN => dp_alu_out_ex_o_14_port);
   dp_ex_stage_alu_U227 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n291, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n170);
   dp_ex_stage_alu_U226 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n170, B2 =>
                           dp_ex_stage_alu_n234, C1 => dp_ex_stage_alu_n171, C2
                           => dp_ex_stage_alu_n291, A => dp_ex_stage_alu_n172, 
                           ZN => dp_alu_out_ex_o_15_port);
   dp_ex_stage_alu_U225 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n215, B2 => 
                           dp_ex_stage_alu_n285, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n94);
   dp_ex_stage_alu_U224 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n94, B2 => 
                           dp_ex_stage_alu_n227, C1 => dp_ex_stage_alu_n95, C2 
                           => dp_ex_stage_alu_n285, A => dp_ex_stage_alu_n96, 
                           ZN => dp_alu_out_ex_o_9_port);
   dp_ex_stage_alu_U223 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n284, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n98);
   dp_ex_stage_alu_U222 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n98, B2 => 
                           dp_ex_stage_alu_n226, C1 => dp_ex_stage_alu_n99, C2 
                           => dp_ex_stage_alu_n284, A => dp_ex_stage_alu_n100, 
                           ZN => dp_alu_out_ex_o_8_port);
   dp_ex_stage_alu_U221 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n215, B2 => 
                           dp_ex_stage_alu_n286, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n185);
   dp_ex_stage_alu_U220 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n185, B2 =>
                           dp_ex_stage_alu_n228, C1 => dp_ex_stage_alu_n186, C2
                           => dp_ex_stage_alu_n286, A => dp_ex_stage_alu_n187, 
                           ZN => dp_alu_out_ex_o_10_port);
   dp_ex_stage_alu_U219 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n293, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n164);
   dp_ex_stage_alu_U218 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n287, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n182);
   dp_ex_stage_alu_U217 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n182, B2 =>
                           dp_ex_stage_alu_n229, C1 => dp_ex_stage_alu_n183, C2
                           => dp_ex_stage_alu_n287, A => dp_ex_stage_alu_n184, 
                           ZN => dp_alu_out_ex_o_11_port);
   dp_ex_stage_alu_U216 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n288, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n179);
   dp_ex_stage_alu_U215 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n292, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n167);
   dp_ex_stage_alu_U214 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n167, B2 =>
                           dp_ex_stage_alu_n235, C1 => dp_ex_stage_alu_n168, C2
                           => dp_ex_stage_alu_n292, A => dp_ex_stage_alu_n169, 
                           ZN => dp_alu_out_ex_o_16_port);
   dp_ex_stage_alu_U213 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n281, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n107);
   dp_ex_stage_alu_U212 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n221, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n113);
   dp_ex_stage_alu_U211 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n220, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n122);
   dp_ex_stage_alu_U210 : OAI221_X1 port map( B1 => dp_ex_stage_alu_n122, B2 =>
                           dp_ex_stage_alu_n43, C1 => dp_ex_stage_alu_n123, C2 
                           => dp_ex_stage_alu_n220, A => dp_ex_stage_alu_n124, 
                           ZN => dp_alu_out_ex_o_2_port);
   dp_ex_stage_alu_U209 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n223, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n110);
   dp_ex_stage_alu_U208 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n306, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n119);
   dp_ex_stage_alu_U207 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n307, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n116);
   dp_ex_stage_alu_U206 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n304, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n128);
   dp_ex_stage_alu_U205 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n213, B2 => 
                           dp_ex_stage_alu_n305, A => dp_ex_stage_alu_n202, ZN 
                           => dp_ex_stage_alu_n125);
   dp_ex_stage_alu_U204 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_muxA_out_23_port, B2 => 
                           dp_ex_stage_alu_n207, C1 => dp_ex_stage_alu_n211, C2
                           => dp_ex_stage_alu_n242, A => dp_ex_stage_alu_n200, 
                           ZN => dp_ex_stage_alu_n144);
   dp_ex_stage_alu_U203 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_muxA_out_26_port, B2 => 
                           dp_ex_stage_alu_n207, C1 => dp_ex_stage_alu_n211, C2
                           => dp_ex_stage_alu_n245, A => dp_ex_stage_alu_n200, 
                           ZN => dp_ex_stage_alu_n135);
   dp_ex_stage_alu_U202 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n74, B2 => 
                           dp_ex_stage_alu_n209, C1 => dp_ex_stage_alu_n212, C2
                           => dp_ex_stage_alu_n228, A => dp_ex_stage_alu_n201, 
                           ZN => dp_ex_stage_alu_n186);
   dp_ex_stage_alu_U201 : INV_X1 port map( A => dp_ex_stage_alu_n70, ZN => 
                           dp_ex_stage_alu_n275);
   dp_ex_stage_alu_U200 : INV_X1 port map( A => dp_ex_stage_alu_n76, ZN => 
                           dp_ex_stage_alu_n273);
   dp_ex_stage_alu_U199 : INV_X1 port map( A => dp_ex_stage_muxB_out_5_port, ZN
                           => dp_ex_stage_alu_n281);
   dp_ex_stage_alu_U198 : INV_X1 port map( A => dp_ex_stage_muxB_out_6_port, ZN
                           => dp_ex_stage_alu_n282);
   dp_ex_stage_alu_U197 : INV_X1 port map( A => dp_ex_stage_muxB_out_12_port, 
                           ZN => dp_ex_stage_alu_n288);
   dp_ex_stage_alu_U196 : INV_X1 port map( A => dp_ex_stage_muxB_out_17_port, 
                           ZN => dp_ex_stage_alu_n293);
   dp_ex_stage_alu_U195 : INV_X1 port map( A => dp_ex_stage_muxB_out_24_port, 
                           ZN => dp_ex_stage_alu_n300);
   dp_ex_stage_alu_U194 : INV_X1 port map( A => dp_ex_stage_muxB_out_28_port, 
                           ZN => dp_ex_stage_alu_n304);
   dp_ex_stage_alu_U193 : INV_X1 port map( A => dp_ex_stage_muxB_out_29_port, 
                           ZN => dp_ex_stage_alu_n305);
   dp_ex_stage_alu_U192 : INV_X1 port map( A => dp_ex_stage_muxB_out_7_port, ZN
                           => dp_ex_stage_alu_n283);
   dp_ex_stage_alu_U191 : INV_X1 port map( A => dp_ex_stage_muxB_out_8_port, ZN
                           => dp_ex_stage_alu_n284);
   dp_ex_stage_alu_U190 : INV_X1 port map( A => dp_ex_stage_alu_n35, ZN => 
                           dp_ex_stage_alu_n286);
   dp_ex_stage_alu_U189 : INV_X1 port map( A => dp_ex_stage_muxB_out_11_port, 
                           ZN => dp_ex_stage_alu_n287);
   dp_ex_stage_alu_U188 : INV_X1 port map( A => dp_ex_stage_muxB_out_13_port, 
                           ZN => dp_ex_stage_alu_n289);
   dp_ex_stage_alu_U187 : INV_X1 port map( A => dp_ex_stage_muxB_out_14_port, 
                           ZN => dp_ex_stage_alu_n290);
   dp_ex_stage_alu_U186 : INV_X1 port map( A => dp_ex_stage_muxB_out_16_port, 
                           ZN => dp_ex_stage_alu_n292);
   dp_ex_stage_alu_U185 : INV_X1 port map( A => dp_ex_stage_muxB_out_18_port, 
                           ZN => dp_ex_stage_alu_n294);
   dp_ex_stage_alu_U184 : INV_X1 port map( A => dp_ex_stage_muxB_out_19_port, 
                           ZN => dp_ex_stage_alu_n295);
   dp_ex_stage_alu_U183 : INV_X1 port map( A => dp_ex_stage_muxB_out_9_port, ZN
                           => dp_ex_stage_alu_n285);
   dp_ex_stage_alu_U182 : INV_X1 port map( A => dp_ex_stage_muxB_out_15_port, 
                           ZN => dp_ex_stage_alu_n291);
   dp_ex_stage_alu_U181 : AND3_X1 port map( A1 => dp_ex_stage_alu_n93, A2 => 
                           dp_ex_stage_alu_n272, A3 => dp_ex_stage_alu_n54, ZN 
                           => dp_ex_stage_alu_n66);
   dp_ex_stage_alu_U180 : INV_X1 port map( A => dp_ex_stage_muxB_out_30_port, 
                           ZN => dp_ex_stage_alu_n306);
   dp_ex_stage_alu_U179 : INV_X1 port map( A => dp_ex_stage_muxB_out_31_port, 
                           ZN => dp_ex_stage_alu_n307);
   dp_ex_stage_alu_U178 : AND2_X1 port map( A1 => dp_ex_stage_alu_n271, A2 => 
                           dp_ex_stage_alu_n196, ZN => dp_ex_stage_alu_n208);
   dp_ex_stage_alu_U177 : BUF_X1 port map( A => dp_ex_stage_alu_n97, Z => 
                           dp_ex_stage_alu_n217);
   dp_ex_stage_alu_U176 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_4_port, A2 => 
                           dp_ex_stage_alu_n196, B1 => 
                           dp_ex_stage_alu_adder_out_4_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n112);
   dp_ex_stage_alu_U175 : BUF_X1 port map( A => dp_ex_stage_alu_n68, Z => 
                           dp_ex_stage_alu_n195);
   dp_ex_stage_alu_U174 : BUF_X1 port map( A => dp_ex_stage_alu_n97, Z => 
                           dp_ex_stage_alu_n218);
   dp_ex_stage_alu_U173 : BUF_X1 port map( A => dp_ex_stage_alu_n97, Z => 
                           dp_ex_stage_alu_n216);
   dp_ex_stage_alu_U172 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_8_port, A2 => 
                           dp_ex_stage_alu_n196, B1 => 
                           dp_ex_stage_alu_adder_out_8_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n100);
   dp_ex_stage_alu_U171 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_16_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_16_port, B2 => 
                           dp_ex_stage_alu_n218, ZN => dp_ex_stage_alu_n169);
   dp_ex_stage_alu_U170 : INV_X1 port map( A => dp_ex_stage_muxA_out_30_port, 
                           ZN => dp_ex_stage_alu_n280);
   dp_ex_stage_alu_U169 : BUF_X1 port map( A => dp_ex_stage_alu_n68, Z => 
                           dp_ex_stage_alu_n196);
   dp_ex_stage_alu_U168 : INV_X1 port map( A => dp_ex_stage_muxA_out_29_port, 
                           ZN => dp_ex_stage_alu_n279);
   dp_ex_stage_alu_U167 : INV_X1 port map( A => dp_ex_stage_muxA_out_19_port, 
                           ZN => dp_ex_stage_alu_n277);
   dp_ex_stage_alu_U166 : BUF_X1 port map( A => dp_ex_stage_alu_n68, Z => 
                           dp_ex_stage_alu_n194);
   dp_ex_stage_alu_U165 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_muxA_out_30_port, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n280, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n120);
   dp_ex_stage_alu_U164 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_muxA_out_29_port, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n279, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n126);
   dp_ex_stage_alu_U163 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n204, B2 =>
                           dp_ex_stage_alu_n72, C1 => dp_ex_stage_alu_n210, C2 
                           => dp_ex_stage_alu_n227, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n95);
   dp_ex_stage_alu_U162 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n33, B2 => 
                           dp_ex_stage_alu_n209, C1 => dp_ex_stage_alu_n212, C2
                           => dp_ex_stage_alu_n229, A => dp_ex_stage_alu_n201, 
                           ZN => dp_ex_stage_alu_n183);
   dp_ex_stage_alu_U161 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_muxA_out_19_port, B2 => 
                           dp_ex_stage_alu_n207, C1 => dp_ex_stage_alu_n211, C2
                           => dp_ex_stage_alu_n277, A => dp_ex_stage_alu_n200, 
                           ZN => dp_ex_stage_alu_n159);
   dp_ex_stage_alu_U160 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_15_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_15_port, B2 => 
                           dp_ex_stage_alu_n218, ZN => dp_ex_stage_alu_n172);
   dp_ex_stage_alu_U159 : INV_X1 port map( A => dp_ex_stage_alu_n189, ZN => 
                           dp_ex_stage_alu_n308);
   dp_ex_stage_alu_U158 : INV_X1 port map( A => dp_ex_stage_alu_n188, ZN => 
                           dp_ex_stage_alu_n309);
   dp_ex_stage_alu_U157 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_11_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_11_port, B2 => 
                           dp_ex_stage_alu_n218, ZN => dp_ex_stage_alu_n184);
   dp_ex_stage_alu_U156 : INV_X1 port map( A => dp_ex_stage_alu_n190, ZN => 
                           dp_ex_stage_alu_n310);
   dp_ex_stage_alu_U155 : AOI21_X1 port map( B1 => dp_ex_stage_alu_n214, B2 => 
                           dp_ex_stage_alu_n282, A => dp_ex_stage_alu_n203, ZN 
                           => dp_ex_stage_alu_n104);
   dp_ex_stage_alu_U154 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_5_port, A2 => 
                           dp_ex_stage_alu_n196, B1 => 
                           dp_ex_stage_alu_adder_out_5_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n109);
   dp_ex_stage_alu_U153 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_3_port, A2 => 
                           dp_ex_stage_alu_n196, B1 => 
                           dp_ex_stage_alu_adder_out_3_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n115);
   dp_ex_stage_alu_U152 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_6_port, A2 => 
                           dp_ex_stage_alu_n196, B1 => 
                           dp_ex_stage_alu_adder_out_6_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n106);
   dp_ex_stage_alu_U151 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_17_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_17_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n166);
   dp_ex_stage_alu_U150 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_1_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_1_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n157);
   dp_ex_stage_alu_U149 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_2_port, A2 => 
                           dp_ex_stage_alu_n195, B1 => 
                           dp_ex_stage_alu_adder_out_2_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n124);
   dp_ex_stage_alu_U148 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_7_port, A2 => 
                           dp_ex_stage_alu_n196, B1 => 
                           dp_ex_stage_alu_adder_out_7_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n103);
   dp_ex_stage_alu_U147 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_9_port, A2 => 
                           dp_ex_stage_alu_n196, B1 => 
                           dp_ex_stage_alu_adder_out_9_port, B2 => 
                           dp_ex_stage_alu_n216, ZN => dp_ex_stage_alu_n96);
   dp_ex_stage_alu_U146 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_18_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_18_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n163);
   dp_ex_stage_alu_U145 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_13_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_13_port, B2 => 
                           dp_ex_stage_alu_n218, ZN => dp_ex_stage_alu_n178);
   dp_ex_stage_alu_U144 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_14_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_14_port, B2 => 
                           dp_ex_stage_alu_n218, ZN => dp_ex_stage_alu_n175);
   dp_ex_stage_alu_U143 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_10_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_10_port, B2 => 
                           dp_ex_stage_alu_n218, ZN => dp_ex_stage_alu_n187);
   dp_ex_stage_alu_U142 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_19_port, A2 => 
                           dp_ex_stage_alu_n194, B1 => 
                           dp_ex_stage_alu_adder_out_19_port, B2 => 
                           dp_ex_stage_alu_n217, ZN => dp_ex_stage_alu_n160);
   dp_ex_stage_alu_U141 : BUF_X1 port map( A => dp_ex_stage_alu_n308, Z => 
                           dp_ex_stage_alu_n198);
   dp_ex_stage_alu_U140 : BUF_X1 port map( A => dp_ex_stage_alu_n308, Z => 
                           dp_ex_stage_alu_n197);
   dp_ex_stage_alu_U139 : BUF_X1 port map( A => dp_ex_stage_alu_n309, Z => 
                           dp_ex_stage_alu_n209);
   dp_ex_stage_alu_U138 : BUF_X1 port map( A => dp_ex_stage_alu_n309, Z => 
                           dp_ex_stage_alu_n207);
   dp_ex_stage_alu_U137 : BUF_X1 port map( A => dp_ex_stage_alu_n309, Z => 
                           dp_ex_stage_alu_n204);
   dp_ex_stage_alu_U136 : BUF_X1 port map( A => dp_ex_stage_alu_n310, Z => 
                           dp_ex_stage_alu_n211);
   dp_ex_stage_alu_U135 : BUF_X1 port map( A => dp_ex_stage_alu_n310, Z => 
                           dp_ex_stage_alu_n213);
   dp_ex_stage_alu_U134 : BUF_X1 port map( A => dp_ex_stage_alu_n310, Z => 
                           dp_ex_stage_alu_n212);
   dp_ex_stage_alu_U133 : BUF_X1 port map( A => dp_ex_stage_alu_n310, Z => 
                           dp_ex_stage_alu_n210);
   dp_ex_stage_alu_U132 : BUF_X1 port map( A => dp_ex_stage_alu_n310, Z => 
                           dp_ex_stage_alu_n214);
   dp_ex_stage_alu_U131 : BUF_X1 port map( A => dp_ex_stage_alu_n197, Z => 
                           dp_ex_stage_alu_n200);
   dp_ex_stage_alu_U130 : BUF_X1 port map( A => dp_ex_stage_alu_n197, Z => 
                           dp_ex_stage_alu_n201);
   dp_ex_stage_alu_U129 : BUF_X1 port map( A => dp_ex_stage_alu_n198, Z => 
                           dp_ex_stage_alu_n202);
   dp_ex_stage_alu_U128 : BUF_X1 port map( A => dp_ex_stage_alu_n197, Z => 
                           dp_ex_stage_alu_n199);
   dp_ex_stage_alu_U127 : BUF_X1 port map( A => dp_ex_stage_alu_n198, Z => 
                           dp_ex_stage_alu_n203);
   dp_ex_stage_alu_U126 : INV_X2 port map( A => dp_ex_stage_alu_n232, ZN => 
                           dp_ex_stage_alu_n231);
   dp_ex_stage_alu_U125 : OR2_X1 port map( A1 => dp_ex_stage_alu_n141, A2 => 
                           dp_ex_stage_alu_n300, ZN => dp_ex_stage_alu_n65);
   dp_ex_stage_alu_U124 : OR2_X1 port map( A1 => dp_ex_stage_alu_n140, A2 => 
                           dp_ex_stage_alu_n243, ZN => dp_ex_stage_alu_n64);
   dp_ex_stage_alu_U123 : OR2_X1 port map( A1 => dp_ex_stage_alu_n117, A2 => 
                           dp_ex_stage_alu_n307, ZN => dp_ex_stage_alu_n63);
   dp_ex_stage_alu_U122 : OR2_X1 port map( A1 => dp_ex_stage_alu_n116, A2 => 
                           dp_ex_stage_alu_n249, ZN => dp_ex_stage_alu_n62);
   dp_ex_stage_alu_U121 : INV_X1 port map( A => alu_op_i_2_port, ZN => 
                           dp_ex_stage_alu_n61);
   dp_ex_stage_alu_U120 : OR2_X1 port map( A1 => dp_ex_stage_alu_n126, A2 => 
                           dp_ex_stage_alu_n305, ZN => dp_ex_stage_alu_n60);
   dp_ex_stage_alu_U119 : OR2_X1 port map( A1 => dp_ex_stage_alu_n125, A2 => 
                           dp_ex_stage_alu_n279, ZN => dp_ex_stage_alu_n59);
   dp_ex_stage_alu_U118 : OR2_X1 port map( A1 => dp_ex_stage_alu_n120, A2 => 
                           dp_ex_stage_alu_n306, ZN => dp_ex_stage_alu_n58);
   dp_ex_stage_alu_U117 : OR2_X1 port map( A1 => dp_ex_stage_alu_n119, A2 => 
                           dp_ex_stage_alu_n280, ZN => dp_ex_stage_alu_n57);
   dp_ex_stage_alu_U116 : OR2_X1 port map( A1 => dp_ex_stage_alu_n129, A2 => 
                           dp_ex_stage_alu_n304, ZN => dp_ex_stage_alu_n56);
   dp_ex_stage_alu_U115 : OR2_X1 port map( A1 => dp_ex_stage_alu_n128, A2 => 
                           dp_ex_stage_alu_n248, ZN => dp_ex_stage_alu_n55);
   dp_ex_stage_alu_U114 : AOI221_X4 port map( B1 => dp_ex_stage_alu_n247, B2 =>
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n248, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n129);
   dp_ex_stage_alu_U113 : NOR2_X1 port map( A1 => dp_ex_stage_alu_n259, A2 => 
                           dp_ex_stage_alu_n17, ZN => dp_ex_stage_alu_n260);
   dp_ex_stage_alu_U112 : NOR2_X1 port map( A1 => dp_ex_stage_alu_n260, A2 => 
                           dp_ex_stage_alu_n53, ZN => dp_ex_stage_alu_n266);
   dp_ex_stage_alu_U111 : AND2_X1 port map( A1 => dp_ex_stage_alu_n45, A2 => 
                           dp_ex_stage_alu_n261, ZN => dp_ex_stage_alu_n53);
   dp_ex_stage_alu_U110 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n130, A2 => 
                           dp_ex_stage_alu_n16, ZN => dp_alu_out_ex_o_28_port);
   dp_ex_stage_alu_U109 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n133, A2 => 
                           dp_ex_stage_alu_n15, ZN => dp_alu_out_ex_o_27_port);
   dp_ex_stage_alu_U108 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n139, A2 => 
                           dp_ex_stage_alu_n14, ZN => dp_alu_out_ex_o_25_port);
   dp_ex_stage_alu_U107 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n142, A2 => 
                           dp_ex_stage_alu_n11, ZN => dp_alu_out_ex_o_24_port);
   dp_ex_stage_alu_U106 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n145, A2 => 
                           dp_ex_stage_alu_n6, ZN => dp_alu_out_ex_o_23_port);
   dp_ex_stage_alu_U105 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n151, A2 => 
                           dp_ex_stage_alu_n10, ZN => dp_alu_out_ex_o_21_port);
   dp_ex_stage_alu_U104 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n154, A2 => 
                           dp_ex_stage_alu_n9, ZN => dp_alu_out_ex_o_20_port);
   dp_ex_stage_alu_U103 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n118, A2 => 
                           dp_ex_stage_alu_n7, ZN => dp_alu_out_ex_o_31_port);
   dp_ex_stage_alu_U102 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n121, A2 => 
                           dp_ex_stage_alu_n5, ZN => dp_alu_out_ex_o_30_port);
   dp_ex_stage_alu_U101 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n127, A2 => 
                           dp_ex_stage_alu_n4, ZN => dp_alu_out_ex_o_29_port);
   dp_ex_stage_alu_U100 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n136, A2 => 
                           dp_ex_stage_alu_n3, ZN => dp_alu_out_ex_o_26_port);
   dp_ex_stage_alu_U99 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n148, A2 => 
                           dp_ex_stage_alu_n8, ZN => dp_alu_out_ex_o_22_port);
   dp_ex_stage_alu_U98 : AOI221_X4 port map( B1 => dp_ex_stage_alu_n231, B2 => 
                           dp_ex_stage_alu_n209, C1 => dp_ex_stage_alu_n212, C2
                           => dp_ex_stage_alu_n232, A => dp_ex_stage_alu_n201, 
                           ZN => dp_ex_stage_alu_n177);
   dp_ex_stage_alu_U97 : OAI21_X2 port map( B1 => dp_ex_stage_alu_n90, B2 => 
                           dp_ex_stage_alu_n311, A => dp_ex_stage_alu_n91, ZN 
                           => dp_ex_stage_alu_N23_port);
   dp_ex_stage_alu_U96 : AOI221_X4 port map( B1 => dp_ex_stage_alu_n71, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n226, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n99);
   dp_ex_stage_alu_U95 : BUF_X2 port map( A => dp_ex_stage_muxA_out_9_port, Z 
                           => dp_ex_stage_alu_n72);
   dp_ex_stage_alu_U94 : NAND3_X1 port map( A1 => dp_ex_stage_alu_n47, A2 => 
                           dp_ex_stage_alu_n48, A3 => dp_ex_stage_alu_n157, ZN 
                           => dp_alu_out_ex_o_1_port);
   dp_ex_stage_alu_U93 : OR2_X1 port map( A1 => dp_ex_stage_alu_n156, A2 => 
                           dp_ex_stage_alu_n219, ZN => dp_ex_stage_alu_n48);
   dp_ex_stage_alu_U92 : OR2_X1 port map( A1 => dp_ex_stage_alu_n155, A2 => 
                           dp_ex_stage_alu_n273, ZN => dp_ex_stage_alu_n47);
   dp_ex_stage_alu_U91 : BUF_X1 port map( A => dp_ex_stage_alu_n30, Z => 
                           dp_ex_stage_alu_n74);
   dp_ex_stage_alu_U90 : BUF_X4 port map( A => dp_ex_stage_muxB_out_0_port, Z 
                           => dp_ex_stage_alu_n45);
   dp_ex_stage_alu_U89 : BUF_X2 port map( A => dp_ex_stage_muxA_out_1_port, Z 
                           => dp_ex_stage_alu_n76);
   dp_ex_stage_alu_U88 : INV_X2 port map( A => dp_ex_stage_alu_n43, ZN => 
                           dp_ex_stage_alu_n44);
   dp_ex_stage_alu_U87 : INV_X1 port map( A => dp_ex_stage_muxA_out_2_port, ZN 
                           => dp_ex_stage_alu_n43);
   dp_ex_stage_alu_U86 : AOI221_X4 port map( B1 => dp_ex_stage_muxA_out_18_port
                           , B2 => dp_ex_stage_alu_n207, C1 => 
                           dp_ex_stage_alu_n212, C2 => dp_ex_stage_alu_n237, A 
                           => dp_ex_stage_alu_n201, ZN => dp_ex_stage_alu_n162)
                           ;
   dp_ex_stage_alu_U85 : NAND3_X1 port map( A1 => dp_ex_stage_alu_n41, A2 => 
                           dp_ex_stage_alu_n42, A3 => dp_ex_stage_alu_n163, ZN 
                           => dp_alu_out_ex_o_18_port);
   dp_ex_stage_alu_U84 : OR2_X1 port map( A1 => dp_ex_stage_alu_n162, A2 => 
                           dp_ex_stage_alu_n294, ZN => dp_ex_stage_alu_n42);
   dp_ex_stage_alu_U83 : OR2_X1 port map( A1 => dp_ex_stage_alu_n161, A2 => 
                           dp_ex_stage_alu_n237, ZN => dp_ex_stage_alu_n41);
   dp_ex_stage_alu_U82 : NAND4_X1 port map( A1 => dp_ex_stage_alu_n26, A2 => 
                           dp_ex_stage_alu_n271, A3 => dp_ex_stage_alu_n61, A4 
                           => dp_ex_stage_alu_n269, ZN => dp_ex_stage_alu_n40);
   dp_ex_stage_alu_U81 : CLKBUF_X1 port map( A => dp_ex_stage_alu_n241, Z => 
                           dp_ex_stage_alu_n39);
   dp_ex_stage_alu_U80 : INV_X2 port map( A => dp_ex_stage_alu_n235, ZN => 
                           dp_ex_stage_alu_n38);
   dp_ex_stage_alu_U79 : BUF_X2 port map( A => dp_ex_stage_muxA_out_8_port, Z 
                           => dp_ex_stage_alu_n71);
   dp_ex_stage_alu_U78 : NOR3_X1 port map( A1 => dp_ex_stage_alu_n36, A2 => 
                           dp_ex_stage_alu_n37, A3 => dp_ex_stage_alu_n264, ZN 
                           => dp_ex_stage_alu_n265);
   dp_ex_stage_alu_U77 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_out_0_port, A2 => 
                           dp_ex_stage_alu_n218, ZN => dp_ex_stage_alu_n37);
   dp_ex_stage_alu_U76 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_out_0_port, A2 => 
                           dp_ex_stage_alu_n196, ZN => dp_ex_stage_alu_n36);
   dp_ex_stage_alu_U75 : AOI221_X4 port map( B1 => dp_ex_stage_alu_n238, B2 => 
                           dp_ex_stage_alu_n207, C1 => dp_ex_stage_alu_n211, C2
                           => dp_ex_stage_alu_n239, A => dp_ex_stage_alu_n200, 
                           ZN => dp_ex_stage_alu_n150);
   dp_ex_stage_alu_U74 : INV_X1 port map( A => dp_ex_stage_alu_n248, ZN => 
                           dp_ex_stage_alu_n247);
   dp_ex_stage_alu_U73 : BUF_X1 port map( A => dp_ex_stage_muxB_out_2_port, Z 
                           => dp_ex_stage_alu_n73);
   dp_ex_stage_alu_U72 : CLKBUF_X1 port map( A => dp_ex_stage_muxB_out_10_port,
                           Z => dp_ex_stage_alu_n35);
   dp_ex_stage_alu_U71 : BUF_X2 port map( A => dp_ex_stage_muxA_out_11_port, Z 
                           => dp_ex_stage_alu_n33);
   dp_ex_stage_alu_U70 : CLKBUF_X1 port map( A => dp_ex_stage_muxA_out_12_port,
                           Z => dp_ex_stage_alu_n32);
   dp_ex_stage_alu_U69 : CLKBUF_X1 port map( A => dp_ex_stage_muxA_out_5_port, 
                           Z => dp_ex_stage_alu_n70);
   dp_ex_stage_alu_U68 : BUF_X4 port map( A => dp_ex_stage_muxB_out_3_port, Z 
                           => dp_ex_stage_alu_n31);
   dp_ex_stage_alu_U67 : INV_X1 port map( A => dp_ex_stage_alu_n239, ZN => 
                           dp_ex_stage_alu_n238);
   dp_ex_stage_alu_U66 : CLKBUF_X1 port map( A => dp_ex_stage_muxA_out_10_port,
                           Z => dp_ex_stage_alu_n30);
   dp_ex_stage_alu_U65 : BUF_X2 port map( A => dp_ex_stage_muxA_out_6_port, Z 
                           => dp_ex_stage_alu_n78);
   dp_ex_stage_alu_U64 : BUF_X2 port map( A => dp_ex_stage_muxA_out_3_port, Z 
                           => dp_ex_stage_alu_n69);
   dp_ex_stage_alu_U63 : BUF_X2 port map( A => dp_ex_stage_muxA_out_15_port, Z 
                           => dp_ex_stage_alu_n29);
   dp_ex_stage_alu_U62 : AOI221_X4 port map( B1 => dp_ex_stage_muxA_out_17_port
                           , B2 => dp_ex_stage_alu_n207, C1 => 
                           dp_ex_stage_alu_n211, C2 => dp_ex_stage_alu_n236, A 
                           => dp_ex_stage_alu_n200, ZN => dp_ex_stage_alu_n165)
                           ;
   dp_ex_stage_alu_U61 : NOR2_X1 port map( A1 => dp_ex_stage_alu_n256, A2 => 
                           dp_ex_stage_alu_n28, ZN => dp_ex_stage_alu_n257);
   dp_ex_stage_alu_U60 : AND2_X1 port map( A1 => dp_ex_stage_alu_N21_port, A2 
                           => dp_ex_stage_alu_n24, ZN => dp_ex_stage_alu_n28);
   dp_ex_stage_alu_U59 : CLKBUF_X3 port map( A => dp_ex_stage_muxB_out_1_port, 
                           Z => dp_ex_stage_alu_n46);
   dp_ex_stage_alu_U58 : NOR2_X1 port map( A1 => alu_op_i_2_port, A2 => 
                           alu_op_i_3_port, ZN => dp_ex_stage_alu_n54);
   dp_ex_stage_alu_U57 : INV_X1 port map( A => alu_op_i_4_port, ZN => 
                           dp_ex_stage_alu_n27);
   dp_ex_stage_alu_U56 : INV_X1 port map( A => alu_op_i_0_port, ZN => 
                           dp_ex_stage_alu_n272);
   dp_ex_stage_alu_U55 : CLKBUF_X1 port map( A => dp_ex_stage_alu_n272, Z => 
                           dp_ex_stage_alu_n26);
   dp_ex_stage_alu_U54 : INV_X1 port map( A => dp_ex_stage_alu_n278, ZN => 
                           dp_ex_stage_alu_n25);
   dp_ex_stage_alu_U53 : AND2_X1 port map( A1 => alu_op_i_0_port, A2 => 
                           alu_op_i_1_port, ZN => dp_ex_stage_alu_n67);
   dp_ex_stage_alu_U52 : CLKBUF_X1 port map( A => dp_ex_stage_alu_n67, Z => 
                           dp_ex_stage_alu_n24);
   dp_ex_stage_alu_U51 : BUF_X1 port map( A => dp_ex_stage_alu_n23, Z => 
                           dp_ex_stage_alu_n52);
   dp_ex_stage_alu_U50 : BUF_X1 port map( A => dp_ex_stage_muxA_out_4_port, Z 
                           => dp_ex_stage_alu_n23);
   dp_ex_stage_alu_U49 : BUF_X2 port map( A => dp_ex_stage_muxB_out_3_port, Z 
                           => dp_ex_stage_alu_n77);
   dp_ex_stage_alu_U48 : INV_X1 port map( A => dp_ex_stage_alu_n93, ZN => 
                           dp_ex_stage_alu_n51);
   dp_ex_stage_alu_U47 : CLKBUF_X1 port map( A => dp_ex_stage_muxB_out_4_port, 
                           Z => dp_ex_stage_alu_n22);
   dp_ex_stage_alu_U46 : BUF_X2 port map( A => dp_ex_stage_muxA_out_0_port, Z 
                           => dp_ex_stage_alu_shifter_N202);
   dp_ex_stage_alu_U45 : CLKBUF_X1 port map( A => dp_ex_stage_alu_N23_port, Z 
                           => dp_ex_stage_alu_n20);
   dp_ex_stage_alu_U44 : NAND3_X1 port map( A1 => dp_ex_stage_alu_n18, A2 => 
                           dp_ex_stage_alu_n19, A3 => dp_ex_stage_alu_n160, ZN 
                           => dp_alu_out_ex_o_19_port);
   dp_ex_stage_alu_U43 : OR2_X1 port map( A1 => dp_ex_stage_alu_n159, A2 => 
                           dp_ex_stage_alu_n295, ZN => dp_ex_stage_alu_n19);
   dp_ex_stage_alu_U42 : OR2_X1 port map( A1 => dp_ex_stage_alu_n158, A2 => 
                           dp_ex_stage_alu_n277, ZN => dp_ex_stage_alu_n18);
   dp_ex_stage_alu_U41 : CLKBUF_X1 port map( A => dp_ex_stage_muxB_out_2_port, 
                           Z => dp_ex_stage_alu_n50);
   dp_ex_stage_alu_U40 : BUF_X1 port map( A => dp_ex_stage_muxA_out_0_port, Z 
                           => dp_ex_stage_alu_n21);
   dp_ex_stage_alu_U39 : OR2_X1 port map( A1 => dp_ex_stage_alu_n2, A2 => 
                           dp_ex_stage_alu_n61, ZN => dp_ex_stage_alu_n17);
   dp_ex_stage_alu_U38 : AND2_X1 port map( A1 => dp_ex_stage_alu_n56, A2 => 
                           dp_ex_stage_alu_n55, ZN => dp_ex_stage_alu_n16);
   dp_ex_stage_alu_U37 : AND2_X1 port map( A1 => dp_ex_stage_alu_n88, A2 => 
                           dp_ex_stage_alu_n87, ZN => dp_ex_stage_alu_n15);
   dp_ex_stage_alu_U36 : AND2_X1 port map( A1 => dp_ex_stage_alu_n84, A2 => 
                           dp_ex_stage_alu_n83, ZN => dp_ex_stage_alu_n14);
   dp_ex_stage_alu_U35 : AND2_X1 port map( A1 => dp_ex_stage_alu_n65, A2 => 
                           dp_ex_stage_alu_n64, ZN => dp_ex_stage_alu_n11);
   dp_ex_stage_alu_U34 : AND2_X1 port map( A1 => dp_ex_stage_alu_n80, A2 => 
                           dp_ex_stage_alu_n79, ZN => dp_ex_stage_alu_n10);
   dp_ex_stage_alu_U33 : AND2_X1 port map( A1 => dp_ex_stage_alu_n193, A2 => 
                           dp_ex_stage_alu_n192, ZN => dp_ex_stage_alu_n9);
   dp_ex_stage_alu_U32 : AND2_X1 port map( A1 => dp_ex_stage_alu_n82, A2 => 
                           dp_ex_stage_alu_n81, ZN => dp_ex_stage_alu_n8);
   dp_ex_stage_alu_U31 : AND2_X1 port map( A1 => dp_ex_stage_alu_n63, A2 => 
                           dp_ex_stage_alu_n62, ZN => dp_ex_stage_alu_n7);
   dp_ex_stage_alu_U30 : AND2_X1 port map( A1 => dp_ex_stage_alu_n92, A2 => 
                           dp_ex_stage_alu_n89, ZN => dp_ex_stage_alu_n6);
   dp_ex_stage_alu_U29 : AND2_X1 port map( A1 => dp_ex_stage_alu_n58, A2 => 
                           dp_ex_stage_alu_n57, ZN => dp_ex_stage_alu_n5);
   dp_ex_stage_alu_U28 : AND2_X1 port map( A1 => dp_ex_stage_alu_n60, A2 => 
                           dp_ex_stage_alu_n59, ZN => dp_ex_stage_alu_n4);
   dp_ex_stage_alu_U27 : AND2_X1 port map( A1 => dp_ex_stage_alu_n86, A2 => 
                           dp_ex_stage_alu_n85, ZN => dp_ex_stage_alu_n3);
   dp_ex_stage_alu_U26 : CLKBUF_X2 port map( A => dp_ex_stage_muxB_out_2_port, 
                           Z => dp_ex_stage_alu_n49);
   dp_ex_stage_alu_U25 : INV_X1 port map( A => dp_ex_stage_alu_n269, ZN => 
                           dp_ex_stage_alu_n2);
   dp_ex_stage_alu_U24 : INV_X1 port map( A => dp_ex_stage_alu_n248, ZN => 
                           dp_ex_stage_alu_n1);
   dp_ex_stage_alu_U23 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n76, B2 => 
                           dp_ex_stage_alu_n207, C1 => dp_ex_stage_alu_n211, C2
                           => dp_ex_stage_alu_n273, A => dp_ex_stage_alu_n200, 
                           ZN => dp_ex_stage_alu_n156);
   dp_ex_stage_alu_U22 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n44, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n43, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n123);
   dp_ex_stage_alu_U21 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n69, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n224, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n114);
   dp_ex_stage_alu_U20 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n52, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n274, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n111);
   dp_ex_stage_alu_U19 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n70, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n275, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n108);
   dp_ex_stage_alu_U18 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n78, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n276, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n105);
   dp_ex_stage_alu_U17 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n34, B2 => 
                           dp_ex_stage_alu_n204, C1 => dp_ex_stage_alu_n210, C2
                           => dp_ex_stage_alu_n225, A => dp_ex_stage_alu_n199, 
                           ZN => dp_ex_stage_alu_n102);
   dp_ex_stage_alu_U16 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n32, B2 => 
                           dp_ex_stage_alu_n209, C1 => dp_ex_stage_alu_n212, C2
                           => dp_ex_stage_alu_n230, A => dp_ex_stage_alu_n201, 
                           ZN => dp_ex_stage_alu_n180);
   dp_ex_stage_alu_U15 : AOI221_X1 port map( B1 => dp_ex_stage_muxA_out_14_port
                           , B2 => dp_ex_stage_alu_n209, C1 => 
                           dp_ex_stage_alu_n211, C2 => dp_ex_stage_alu_n233, A 
                           => dp_ex_stage_alu_n200, ZN => dp_ex_stage_alu_n174)
                           ;
   dp_ex_stage_alu_U14 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n29, B2 => 
                           dp_ex_stage_alu_n209, C1 => dp_ex_stage_alu_n212, C2
                           => dp_ex_stage_alu_n234, A => dp_ex_stage_alu_n201, 
                           ZN => dp_ex_stage_alu_n171);
   dp_ex_stage_alu_U13 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n38, B2 => 
                           dp_ex_stage_alu_n209, C1 => dp_ex_stage_alu_n212, C2
                           => dp_ex_stage_alu_n235, A => dp_ex_stage_alu_n201, 
                           ZN => dp_ex_stage_alu_n168);
   dp_ex_stage_alu_U12 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n25, B2 => 
                           dp_ex_stage_alu_n207, C1 => dp_ex_stage_alu_n211, C2
                           => dp_ex_stage_alu_n278, A => dp_ex_stage_alu_n200, 
                           ZN => dp_ex_stage_alu_n153);
   dp_ex_stage_alu_U11 : AOI221_X1 port map( B1 => dp_ex_stage_alu_n240, B2 => 
                           dp_ex_stage_alu_n207, C1 => dp_ex_stage_alu_n211, C2
                           => dp_ex_stage_alu_n39, A => dp_ex_stage_alu_n200, 
                           ZN => dp_ex_stage_alu_n147);
   dp_ex_stage_alu_U10 : AOI221_X1 port map( B1 => dp_ex_stage_muxA_out_24_port
                           , B2 => dp_ex_stage_alu_n207, C1 => 
                           dp_ex_stage_alu_n211, C2 => dp_ex_stage_alu_n243, A 
                           => dp_ex_stage_alu_n200, ZN => dp_ex_stage_alu_n141)
                           ;
   dp_ex_stage_alu_U9 : AOI221_X1 port map( B1 => dp_ex_stage_muxA_out_25_port,
                           B2 => dp_ex_stage_alu_n207, C1 => 
                           dp_ex_stage_alu_n211, C2 => dp_ex_stage_alu_n244, A 
                           => dp_ex_stage_alu_n200, ZN => dp_ex_stage_alu_n138)
                           ;
   dp_ex_stage_alu_U8 : AOI221_X1 port map( B1 => dp_ex_stage_muxA_out_27_port,
                           B2 => dp_ex_stage_alu_n207, C1 => 
                           dp_ex_stage_alu_n211, C2 => dp_ex_stage_alu_n246, A 
                           => dp_ex_stage_alu_n200, ZN => dp_ex_stage_alu_n132)
                           ;
   dp_ex_stage_alu_U7 : AOI221_X1 port map( B1 => dp_ex_stage_muxA_out_31_port,
                           B2 => dp_ex_stage_alu_n204, C1 => 
                           dp_ex_stage_alu_n210, C2 => dp_ex_stage_alu_n249, A 
                           => dp_ex_stage_alu_n199, ZN => dp_ex_stage_alu_n117)
                           ;
   dp_ex_stage_alu_U5 : BUF_X2 port map( A => dp_ex_stage_muxA_out_7_port, Z =>
                           dp_ex_stage_alu_n34);
   dp_ex_stage_alu_U4 : MUX2_X1 port map( A => dp_ex_stage_alu_n255, B => 
                           dp_ex_stage_alu_N19_port, S => dp_ex_stage_alu_n51, 
                           Z => dp_ex_stage_alu_n256);
   dp_ex_stage_alu_U235 : NAND3_X1 port map( A1 => dp_ex_stage_alu_n93, A2 => 
                           dp_ex_stage_alu_n270, A3 => dp_ex_stage_alu_n191, ZN
                           => dp_ex_stage_alu_n206);
   dp_ex_stage_alu_U230 : NAND3_X1 port map( A1 => alu_op_i_4_port, A2 => 
                           dp_ex_stage_alu_n54, A3 => dp_ex_stage_alu_n67, ZN 
                           => dp_ex_stage_alu_n91);
   dp_ex_stage_alu_n13 <= '1';
   dp_ex_stage_alu_n12 <= '0';
   dp_ex_stage_alu_Logic1_port <= '1';
   dp_ex_stage_alu_adder_U53 : OR2_X1 port map( A1 => dp_ex_stage_alu_n20, A2 
                           => dp_ex_stage_alu_adder_n22, ZN => 
                           dp_ex_stage_alu_adder_carries_0_port);
   dp_ex_stage_alu_adder_U52 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22
                           , B => dp_ex_stage_muxB_out_5_port, Z => 
                           dp_ex_stage_alu_adder_n20);
   dp_ex_stage_alu_adder_U51 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n23
                           , B => dp_ex_stage_muxB_out_15_port, Z => 
                           dp_ex_stage_alu_adder_n18);
   dp_ex_stage_alu_adder_U50 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22
                           , B => dp_ex_stage_alu_n45, Z => 
                           dp_ex_stage_alu_adder_n17);
   dp_ex_stage_alu_adder_U49 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_3_port, Z => 
                           dp_ex_stage_alu_adder_n16);
   dp_ex_stage_alu_adder_U48 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_n20, Z => 
                           dp_ex_stage_alu_adder_n14);
   dp_ex_stage_alu_adder_U47 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_6_port, Z => 
                           dp_ex_stage_alu_adder_n10);
   dp_ex_stage_alu_adder_U46 : BUF_X2 port map( A => dp_ex_stage_alu_N23_port, 
                           Z => dp_ex_stage_alu_adder_n15);
   dp_ex_stage_alu_adder_U45 : BUF_X1 port map( A => dp_ex_stage_alu_N23_port, 
                           Z => dp_ex_stage_alu_adder_n21);
   dp_ex_stage_alu_adder_U44 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n13
                           , B => dp_ex_stage_muxB_out_23_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_23_port);
   dp_ex_stage_alu_adder_U43 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_11_port, Z => 
                           dp_ex_stage_alu_adder_n8);
   dp_ex_stage_alu_adder_U42 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_13_port, Z => 
                           dp_ex_stage_alu_adder_n7);
   dp_ex_stage_alu_adder_U41 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_n15, Z => 
                           dp_ex_stage_alu_adder_n11);
   dp_ex_stage_alu_adder_U40 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n13
                           , B => dp_ex_stage_muxB_out_19_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_19_port);
   dp_ex_stage_alu_adder_U39 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_19_port, Z => 
                           dp_ex_stage_alu_adder_n6);
   dp_ex_stage_alu_adder_U38 : CLKBUF_X3 port map( A => 
                           dp_ex_stage_alu_N23_port, Z => 
                           dp_ex_stage_alu_adder_n23);
   dp_ex_stage_alu_adder_U37 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n12
                           , B => dp_ex_stage_muxB_out_15_port, Z => 
                           dp_ex_stage_alu_adder_n5);
   dp_ex_stage_alu_adder_U36 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_14_port, Z => 
                           dp_ex_stage_alu_adder_n4);
   dp_ex_stage_alu_adder_U35 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n9,
                           B => dp_ex_stage_muxB_out_9_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_9_port);
   dp_ex_stage_alu_adder_U34 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_9_port, Z => 
                           dp_ex_stage_alu_adder_n3);
   dp_ex_stage_alu_adder_U30 : BUF_X2 port map( A => dp_ex_stage_alu_adder_n15,
                           Z => dp_ex_stage_alu_adder_n13);
   dp_ex_stage_alu_adder_U27 : CLKBUF_X3 port map( A => 
                           dp_ex_stage_alu_N23_port, Z => 
                           dp_ex_stage_alu_adder_n22);
   dp_ex_stage_alu_adder_U23 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n21
                           , B => dp_ex_stage_muxB_out_7_port, Z => 
                           dp_ex_stage_alu_adder_n19);
   dp_ex_stage_alu_adder_U18 : CLKBUF_X1 port map( A => dp_ex_stage_alu_n231, Z
                           => dp_ex_stage_alu_adder_n2);
   dp_ex_stage_alu_adder_U6 : BUF_X1 port map( A => dp_ex_stage_alu_adder_n15, 
                           Z => dp_ex_stage_alu_adder_n9);
   dp_ex_stage_alu_adder_U4 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n13,
                           B => dp_ex_stage_muxB_out_23_port, Z => 
                           dp_ex_stage_alu_adder_n1);
   dp_ex_stage_alu_adder_U2 : BUF_X2 port map( A => dp_ex_stage_alu_adder_n15, 
                           Z => dp_ex_stage_alu_adder_n12);
   dp_ex_stage_alu_adder_U1 : XOR2_X2 port map( A => dp_ex_stage_alu_adder_n12,
                           B => dp_ex_stage_muxB_out_12_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_12_port);
   dp_ex_stage_alu_adder_U33 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n21
                           , B => dp_ex_stage_alu_n45, Z => 
                           dp_ex_stage_alu_adder_B_xor_0_port);
   dp_ex_stage_alu_adder_U32 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22
                           , B => dp_ex_stage_alu_n35, Z => 
                           dp_ex_stage_alu_adder_B_xor_10_port);
   dp_ex_stage_alu_adder_U31 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22
                           , B => dp_ex_stage_muxB_out_11_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_11_port);
   dp_ex_stage_alu_adder_U29 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n23
                           , B => dp_ex_stage_muxB_out_13_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_13_port);
   dp_ex_stage_alu_adder_U28 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n12
                           , B => dp_ex_stage_muxB_out_14_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_14_port);
   dp_ex_stage_alu_adder_U26 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n11
                           , B => dp_ex_stage_muxB_out_16_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_16_port);
   dp_ex_stage_alu_adder_U25 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n23
                           , B => dp_ex_stage_muxB_out_17_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_17_port);
   dp_ex_stage_alu_adder_U24 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22
                           , B => dp_ex_stage_muxB_out_18_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_18_port);
   dp_ex_stage_alu_adder_U22 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n21
                           , B => dp_ex_stage_alu_n46, Z => 
                           dp_ex_stage_alu_adder_B_xor_1_port);
   dp_ex_stage_alu_adder_U21 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n12
                           , B => dp_ex_stage_muxB_out_20_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_20_port);
   dp_ex_stage_alu_adder_U20 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n23
                           , B => dp_ex_stage_muxB_out_21_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_21_port);
   dp_ex_stage_alu_adder_U19 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n23
                           , B => dp_ex_stage_muxB_out_22_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_22_port);
   dp_ex_stage_alu_adder_U17 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n11
                           , B => dp_ex_stage_muxB_out_24_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_24_port);
   dp_ex_stage_alu_adder_U16 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22
                           , B => dp_ex_stage_muxB_out_25_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_25_port);
   dp_ex_stage_alu_adder_U15 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n23
                           , B => dp_ex_stage_muxB_out_26_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_26_port);
   dp_ex_stage_alu_adder_U14 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n23
                           , B => dp_ex_stage_muxB_out_27_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_27_port);
   dp_ex_stage_alu_adder_U13 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n23
                           , B => dp_ex_stage_muxB_out_28_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_28_port);
   dp_ex_stage_alu_adder_U12 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22
                           , B => dp_ex_stage_muxB_out_29_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_29_port);
   dp_ex_stage_alu_adder_U11 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22
                           , B => dp_ex_stage_alu_n50, Z => 
                           dp_ex_stage_alu_adder_B_xor_2_port);
   dp_ex_stage_alu_adder_U10 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n12
                           , B => dp_ex_stage_muxB_out_30_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_30_port);
   dp_ex_stage_alu_adder_U9 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n13,
                           B => dp_ex_stage_muxB_out_31_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_31_port);
   dp_ex_stage_alu_adder_U8 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n9, 
                           B => dp_ex_stage_alu_n77, Z => 
                           dp_ex_stage_alu_adder_B_xor_3_port);
   dp_ex_stage_alu_adder_U7 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22,
                           B => dp_ex_stage_alu_n222, Z => 
                           dp_ex_stage_alu_adder_B_xor_4_port);
   dp_ex_stage_alu_adder_U5 : XOR2_X1 port map( A => 
                           dp_ex_stage_muxB_out_6_port, B => 
                           dp_ex_stage_alu_adder_n13, Z => 
                           dp_ex_stage_alu_adder_B_xor_6_port);
   dp_ex_stage_alu_adder_U3 : XOR2_X1 port map( A => dp_ex_stage_alu_adder_n22,
                           B => dp_ex_stage_muxB_out_8_port, Z => 
                           dp_ex_stage_alu_adder_B_xor_8_port);
   dp_ex_stage_alu_adder_SparseTree_U6 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_n1, Z => 
                           dp_ex_stage_alu_adder_carries_2_port);
   dp_ex_stage_alu_adder_SparseTree_U5 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_gen_12_9_port, Z =>
                           dp_ex_stage_alu_adder_SparseTree_n4);
   dp_ex_stage_alu_adder_SparseTree_U4 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_gen_24_17_port, Z 
                           => dp_ex_stage_alu_adder_SparseTree_n3);
   dp_ex_stage_alu_adder_SparseTree_U3 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_n9, Z => 
                           dp_ex_stage_alu_adder_carries_1_port);
   dp_ex_stage_alu_adder_SparseTree_U2 : CLKBUF_X2 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_n7, Z => 
                           dp_ex_stage_alu_adder_carries_4_port);
   dp_ex_stage_alu_adder_SparseTree_U1 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_n8, Z => 
                           dp_ex_stage_alu_adder_SparseTree_n1);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_1_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_0_port, A2 => 
                           dp_ex_stage_alu_shifter_N202, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_1_1_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_1_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_0_port, B => 
                           dp_ex_stage_alu_shifter_N202, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_1_1_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_2_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_1_port, A2 => 
                           dp_ex_stage_alu_n76, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_2_2_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_2_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_1_port, B => 
                           dp_ex_stage_alu_n76, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_2_2_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_3_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_2_port, A2 => 
                           dp_ex_stage_alu_n44, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_3_3_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_3_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_2_port, B => 
                           dp_ex_stage_alu_n44, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_3_3_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_4_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_3_port, A2 => 
                           dp_ex_stage_alu_n69, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_4_4_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_4_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_3_port, B => 
                           dp_ex_stage_alu_n69, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_4_4_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_5_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_4_port, A2 => 
                           dp_ex_stage_alu_n52, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_5_5_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_5_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_4_port, B => 
                           dp_ex_stage_alu_n52, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_5_5_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_6_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_n20, A2 => 
                           dp_ex_stage_muxA_out_5_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_6_6_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_6_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_n20, B => 
                           dp_ex_stage_muxA_out_5_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_6_6_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_7_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_6_port, A2 => 
                           dp_ex_stage_alu_n78, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_7_7_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_7_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_6_port, B => 
                           dp_ex_stage_alu_n78, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_7_7_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_8_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_n19, A2 => dp_ex_stage_alu_n34
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_8_8_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_8_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_n19, B => dp_ex_stage_alu_n34,
                           Z => dp_ex_stage_alu_adder_SparseTree_prop_8_8_port)
                           ;
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_9_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_8_port, A2 => 
                           dp_ex_stage_alu_n71, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_9_9_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_9_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_8_port, B => 
                           dp_ex_stage_alu_n71, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_9_9_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_10_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_9_port, A2 => 
                           dp_ex_stage_alu_n72, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_10_10_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_10_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_9_port, B => 
                           dp_ex_stage_alu_n72, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_10_10_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_11_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_10_port, A2 => 
                           dp_ex_stage_alu_n74, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_11_11_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_11_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_10_port, B => 
                           dp_ex_stage_alu_n74, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_11_11_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_12_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_11_port, A2 => 
                           dp_ex_stage_muxA_out_11_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_12_12_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_12_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_11_port, B => 
                           dp_ex_stage_muxA_out_11_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_12_12_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_13_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_12_port, A2 => 
                           dp_ex_stage_alu_n32, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_13_13_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_13_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_12_port, B => 
                           dp_ex_stage_alu_n32, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_13_13_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_14_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_13_port, A2 => 
                           dp_ex_stage_alu_n231, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_14_14_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_14_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_13_port, B => 
                           dp_ex_stage_alu_n231, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_14_14_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_15_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_14_port, A2 => 
                           dp_ex_stage_muxA_out_14_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_15_15_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_15_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_14_port, B => 
                           dp_ex_stage_muxA_out_14_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_15_15_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_16_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_n18, A2 => dp_ex_stage_alu_n29
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_16_16_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_16_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_n18, B => dp_ex_stage_alu_n29,
                           Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_16_16_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_17_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_16_port, A2 => 
                           dp_ex_stage_alu_n38, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_17_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_17_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_16_port, B => 
                           dp_ex_stage_alu_n38, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_17_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_n1, A2 
                           => dp_ex_stage_muxA_out_17_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_18_18_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_U1 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_17_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_n1);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_18_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_17_port, B => 
                           dp_ex_stage_muxA_out_17_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_18_18_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_19_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_18_port, A2 => 
                           dp_ex_stage_muxA_out_18_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_19_19_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_19_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_18_port, B => 
                           dp_ex_stage_muxA_out_18_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_19_19_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_20_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_19_port, A2 => 
                           dp_ex_stage_alu_adder_B_xor_19_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_20_20_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_20_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_19_port, B => 
                           dp_ex_stage_muxA_out_19_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_20_20_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_21_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_20_port, A2 => 
                           dp_ex_stage_alu_n25, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_21_21_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_21_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_20_port, B => 
                           dp_ex_stage_alu_n25, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_21_21_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_n1, A2 
                           => dp_ex_stage_alu_n238, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_22_22_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_U1 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_21_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_n1);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_22_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_21_port, B => 
                           dp_ex_stage_alu_n238, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_22_22_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_23_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_22_port, A2 => 
                           dp_ex_stage_alu_n240, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_23_23_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_23_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_22_port, B => 
                           dp_ex_stage_alu_n240, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_23_23_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_24_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_23_port, A2 => 
                           dp_ex_stage_muxA_out_23_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_24_24_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_24_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_23_port, B => 
                           dp_ex_stage_muxA_out_23_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_24_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_25_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_24_port, A2 => 
                           dp_ex_stage_muxA_out_24_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_25_25_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_25_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_24_port, B => 
                           dp_ex_stage_muxA_out_24_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_25_25_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_26_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_25_port, A2 => 
                           dp_ex_stage_muxA_out_25_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_26_26_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_26_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_25_port, B => 
                           dp_ex_stage_muxA_out_25_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_26_26_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_27_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_26_port, A2 => 
                           dp_ex_stage_muxA_out_26_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_27_27_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_27_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_26_port, B => 
                           dp_ex_stage_muxA_out_26_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_27_27_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_28_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_27_port, A2 => 
                           dp_ex_stage_muxA_out_27_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_28_28_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_28_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_27_port, B => 
                           dp_ex_stage_muxA_out_27_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_28_28_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_29_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_28_port, A2 => 
                           dp_ex_stage_alu_n247, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_29_29_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_29_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_28_port, B => 
                           dp_ex_stage_alu_n247, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_29_29_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_30_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_29_port, A2 => 
                           dp_ex_stage_muxA_out_29_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_30_30_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_30_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_29_port, B => 
                           dp_ex_stage_muxA_out_29_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_30_30_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_31_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_30_port, A2 => 
                           dp_ex_stage_muxA_out_30_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_31_31_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_31_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_30_port, B => 
                           dp_ex_stage_muxA_out_30_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_31_31_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_32_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_31_port, A2 => 
                           dp_ex_stage_muxA_out_31_port, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_32_32_port);
   dp_ex_stage_alu_adder_SparseTree_PG_net_i_32_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_31_port, B => 
                           dp_ex_stage_muxA_out_31_port, Z => 
                           dp_ex_stage_alu_adder_SparseTree_prop_32_32_port);
   dp_ex_stage_alu_adder_SparseTree_G10_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_1_1_port, B2 
                           => dp_ex_stage_alu_adder_carries_0_port, A => 
                           dp_ex_stage_alu_adder_SparseTree_gen_1_1_port, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_G10_n2);
   dp_ex_stage_alu_adder_SparseTree_G10_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G10_n2, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_1_0_port);
   dp_ex_stage_alu_adder_SparseTree_G20_1_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G20_1_n3, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_gen_2_0_port);
   dp_ex_stage_alu_adder_SparseTree_G20_1_U1 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_1_0_port, B2 =>
                           dp_ex_stage_alu_adder_SparseTree_prop_2_2_port, A =>
                           dp_ex_stage_alu_adder_SparseTree_gen_2_2_port, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_G20_1_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_4_4_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_gen_3_3_port, A 
                           => dp_ex_stage_alu_adder_SparseTree_gen_4_4_port, ZN
                           => dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_n2);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_U2 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_3_3_port, A2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_4_4_port, 
                           ZN => dp_ex_stage_alu_adder_SparseTree_prop_4_3_port
                           );
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_0_n2, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_4_3_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_5_5_port, A2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_6_6_port, 
                           ZN => dp_ex_stage_alu_adder_SparseTree_prop_6_5_port
                           );
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_5_5_port, B2 =>
                           dp_ex_stage_alu_adder_SparseTree_prop_6_6_port, A =>
                           dp_ex_stage_alu_adder_SparseTree_gen_6_6_port, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_1_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_6_5_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_8_8_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_gen_7_7_port, A 
                           => dp_ex_stage_alu_adder_SparseTree_gen_8_8_port, ZN
                           => dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_U2 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_7_7_port, A2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_8_8_port, 
                           ZN => dp_ex_stage_alu_adder_SparseTree_prop_8_7_port
                           );
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_2_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_8_7_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_10_10_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_9_9_port, 
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_10_9_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_10_10_port, B2
                           => dp_ex_stage_alu_adder_SparseTree_gen_9_9_port, A 
                           => dp_ex_stage_alu_adder_SparseTree_gen_10_10_port, 
                           ZN => dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_n3)
                           ;
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_3_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_10_9_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_11_11_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_12_12_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_12_11_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_11_11_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_12_12_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_12_12_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_4_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_12_11_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_13_13_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_14_14_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_14_13_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_14_13_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_U1 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_13_13_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_14_14_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_14_14_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_5_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_16_16_port, B2
                           => dp_ex_stage_alu_adder_SparseTree_gen_15_15_port, 
                           A => dp_ex_stage_alu_adder_SparseTree_gen_16_16_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_U2 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_15_15_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_16_16_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_16_15_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_6_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_16_15_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_18_18_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_17_17_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_18_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_17_17_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_18_18_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_18_18_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_7_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_18_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_19_19_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_20_20_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_20_19_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_20_20_port, B2
                           => dp_ex_stage_alu_adder_SparseTree_gen_19_19_port, 
                           A => dp_ex_stage_alu_adder_SparseTree_gen_20_20_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_8_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_20_19_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_22_22_port, B2
                           => dp_ex_stage_alu_adder_SparseTree_gen_21_21_port, 
                           A => dp_ex_stage_alu_adder_SparseTree_gen_22_22_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_22_21_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_9_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_22_22_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_21_21_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_22_21_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_24_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_23_23_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_23_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_24_port, B2
                           => dp_ex_stage_alu_adder_SparseTree_gen_23_23_port, 
                           A => dp_ex_stage_alu_adder_SparseTree_gen_24_24_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_10_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_gen_24_23_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_25_25_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_26_26_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_26_25_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_25_25_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_26_26_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_26_26_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_11_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_gen_26_25_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_27_27_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_28_28_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_28_27_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_27_27_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_28_28_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_28_28_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_12_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_gen_28_27_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_29_29_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_30_30_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_30_30_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_gen_30_29_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_13_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_29_29_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_30_30_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_30_29_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_31_31_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_32_32_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_32_32_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_gen_32_31_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_1_14_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_31_31_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_32_32_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_32_31_port);
   dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_2_0_port, B2 =>
                           dp_ex_stage_alu_adder_SparseTree_prop_4_3_port, A =>
                           dp_ex_stage_alu_adder_SparseTree_gen_4_3_port, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_n3);
   dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G_2exp_0_2_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_n9);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_8_5_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_6_5_port, B2 =>
                           dp_ex_stage_alu_adder_SparseTree_prop_8_7_port, A =>
                           dp_ex_stage_alu_adder_SparseTree_gen_8_7_port, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_0_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_6_5_port, A2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_8_7_port, 
                           ZN => dp_ex_stage_alu_adder_SparseTree_prop_8_5_port
                           );
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_10_9_port, A2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_12_11_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_12_9_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_10_9_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_12_11_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_12_11_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_1_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_12_9_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_14_13_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_16_15_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_16_13_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_14_13_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_16_15_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_16_15_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_2_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_16_13_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_18_17_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_20_19_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_20_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_18_17_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_20_19_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_20_19_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_3_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_20_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_22_21_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_24_23_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_21_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_22_21_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_24_23_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_24_23_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_4_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_24_21_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_26_25_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_28_27_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_28_25_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_26_25_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_28_27_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_28_27_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_5_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_28_25_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_30_29_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_32_31_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_32_31_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_32_29_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_2_6_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_30_29_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_32_31_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_32_29_port);
   dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_n9, B2 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_8_5_port, A =>
                           dp_ex_stage_alu_adder_SparseTree_gen_8_5_port, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_n3);
   dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G_2exp_0_3_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_n8);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_16_9_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_12_9_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_16_13_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_16_13_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_0_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_12_9_port, A2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_16_13_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_16_9_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_U3 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_20_17_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_24_21_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_20_17_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_24_21_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_24_21_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_3_1_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_24_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_28_25_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_32_29_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_32_29_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_n3, ZN =>
                           dp_ex_stage_alu_adder_SparseTree_gen_32_25_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_3_2_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_28_25_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_32_29_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_32_25_port);
   dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_n8, B2 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_16_9_port, A 
                           => dp_ex_stage_alu_adder_SparseTree_gen_16_9_port, 
                           ZN => dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_n3
                           );
   dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G_2exp_0_4_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_n7);
   dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_12_9_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_n1, A => 
                           dp_ex_stage_alu_adder_SparseTree_n4, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_n3);
   dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G_2n_0_4_1_n3, ZN 
                           => dp_ex_stage_alu_adder_carries_3_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_n3, B2 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_32_25_port, A 
                           => dp_ex_stage_alu_adder_SparseTree_gen_32_25_port, 
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_U2 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_17_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_32_25_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_32_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_4_0_0_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_gen_32_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_U3 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_gen_24_17_port, B2 
                           => dp_ex_stage_alu_adder_SparseTree_prop_28_25_port,
                           A => dp_ex_stage_alu_adder_SparseTree_gen_28_25_port
                           , ZN => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_n3);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_n3, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_gen_28_17_port);
   dp_ex_stage_alu_adder_SparseTree_PG_ij_4_1_0_U1 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_17_port, A2
                           => dp_ex_stage_alu_adder_SparseTree_prop_28_25_port,
                           ZN => 
                           dp_ex_stage_alu_adder_SparseTree_prop_28_17_port);
   dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_32_17_port, B2
                           => dp_ex_stage_alu_adder_carries_4_port, A => 
                           dp_ex_stage_alu_adder_SparseTree_gen_32_17_port, ZN 
                           => dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_n3);
   dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G_2exp_0_5_n3, ZN 
                           => dp_ex_stage_alu_adder_Cout);
   dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_n7, B2 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_28_17_port, A 
                           => dp_ex_stage_alu_adder_SparseTree_gen_28_17_port, 
                           ZN => dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_n3
                           );
   dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_1_n3, ZN 
                           => dp_ex_stage_alu_adder_carries_7_port);
   dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_n3, ZN 
                           => dp_ex_stage_alu_adder_carries_6_port);
   dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_U1 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_n7, B2 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_24_17_port, A 
                           => dp_ex_stage_alu_adder_SparseTree_n3, ZN => 
                           dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_2_n3);
   dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_U2 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_adder_SparseTree_n7, B2 => 
                           dp_ex_stage_alu_adder_SparseTree_prop_20_17_port, A 
                           => dp_ex_stage_alu_adder_SparseTree_gen_20_17_port, 
                           ZN => dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_n3
                           );
   dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SparseTree_G_2n_0_5_3_n3, ZN 
                           => dp_ex_stage_alu_adder_carries_5_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Logic0_port <= '0';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Logic1_port <= '1';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_alu_n69, B => 
                           dp_ex_stage_alu_adder_n16, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_alu_n44, B => 
                           dp_ex_stage_alu_adder_B_xor_2_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_alu_n76, B => 
                           dp_ex_stage_alu_adder_B_xor_1_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_shifter_N202, B => 
                           dp_ex_stage_alu_adder_n17, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Logic0_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA0_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_alu_n69, B => 
                           dp_ex_stage_alu_adder_n16, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_alu_n44, B => 
                           dp_ex_stage_alu_adder_B_xor_2_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_alu_n76, B => 
                           dp_ex_stage_alu_adder_B_xor_1_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_shifter_N202, B => 
                           dp_ex_stage_alu_adder_n17, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Logic1_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_RCA1_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U9 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_0_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_0_port
                           , B2 => dp_ex_stage_alu_adder_carries_0_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n9);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U8 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_3_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5,
                           B1 => dp_ex_stage_alu_adder_carries_0_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_3_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n6)
                           ;
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U7 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n6, ZN => 
                           dp_ex_stage_alu_adder_out_3_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U6 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_0_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U5 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_1_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_1_port
                           , B2 => dp_ex_stage_alu_adder_carries_0_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n8);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U4 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n8, ZN => 
                           dp_ex_stage_alu_adder_out_1_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U3 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out0_2_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_rca_out1_2_port
                           , B2 => dp_ex_stage_alu_adder_carries_0_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n7);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n7, ZN => 
                           dp_ex_stage_alu_adder_out_2_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_0_Mux_n9, ZN => 
                           dp_ex_stage_alu_adder_out_0_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Logic0_port <= '0';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Logic1_port <= '1';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_alu_n34, B => 
                           dp_ex_stage_alu_adder_n19, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_alu_n78, B => 
                           dp_ex_stage_alu_adder_n10, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_5_port, B => 
                           dp_ex_stage_alu_adder_n14, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n52, B => 
                           dp_ex_stage_alu_adder_B_xor_4_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Logic0_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA0_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_alu_n34, B => 
                           dp_ex_stage_alu_adder_n19, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_alu_n78, B => 
                           dp_ex_stage_alu_adder_n10, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_5_port, B => 
                           dp_ex_stage_alu_adder_n14, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n52, B => 
                           dp_ex_stage_alu_adder_B_xor_4_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Logic1_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_RCA1_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U9 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_1_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U8 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_0_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_0_port
                           , B2 => dp_ex_stage_alu_adder_carries_1_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n10);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U7 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_1_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_1_port
                           , B2 => dp_ex_stage_alu_adder_carries_1_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n11);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U6 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_2_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_2_port
                           , B2 => dp_ex_stage_alu_adder_carries_1_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n12);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U5 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out0_3_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n5,
                           B1 => dp_ex_stage_alu_adder_carries_1_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_rca_out1_3_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n13
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U4 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n10, ZN => 
                           dp_ex_stage_alu_adder_out_4_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n11, ZN => 
                           dp_ex_stage_alu_adder_out_5_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n12, ZN => 
                           dp_ex_stage_alu_adder_out_6_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_1_Mux_n13, ZN => 
                           dp_ex_stage_alu_adder_out_7_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Logic0_port <= '0';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Logic1_port <= '1';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_11_port, B => 
                           dp_ex_stage_alu_adder_n8, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_alu_n74, B => 
                           dp_ex_stage_alu_adder_B_xor_10_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_alu_n72, B => 
                           dp_ex_stage_alu_adder_n3, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n71, B => 
                           dp_ex_stage_alu_adder_B_xor_8_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Logic0_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA0_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_11_port, B => 
                           dp_ex_stage_alu_adder_n8, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_alu_n74, B => 
                           dp_ex_stage_alu_adder_B_xor_10_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_alu_n72, B => 
                           dp_ex_stage_alu_adder_n3, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n71, B => 
                           dp_ex_stage_alu_adder_B_xor_8_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Logic1_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_RCA1_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U9 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_2_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U8 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_1_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_1_port
                           , B2 => dp_ex_stage_alu_adder_carries_2_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n11);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U7 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_0_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_0_port
                           , B2 => dp_ex_stage_alu_adder_carries_2_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n10);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U6 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_2_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_2_port
                           , B2 => dp_ex_stage_alu_adder_carries_2_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n12);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U5 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out0_3_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n5,
                           B1 => dp_ex_stage_alu_adder_carries_2_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_rca_out1_3_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n13
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U4 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n10, ZN => 
                           dp_ex_stage_alu_adder_out_8_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n13, ZN => 
                           dp_ex_stage_alu_adder_out_11_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n11, ZN => 
                           dp_ex_stage_alu_adder_out_9_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_2_Mux_n12, ZN => 
                           dp_ex_stage_alu_adder_out_10_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Logic0_port <= '0';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Logic1_port <= '1';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_alu_n29, B => 
                           dp_ex_stage_alu_adder_n5, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_14_port, B => 
                           dp_ex_stage_alu_adder_n4, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_alu_adder_n2, B => 
                           dp_ex_stage_alu_adder_n7, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n32, B => 
                           dp_ex_stage_alu_adder_B_xor_12_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Logic0_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA0_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_alu_n29, B => 
                           dp_ex_stage_alu_adder_n5, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_14_port, B => 
                           dp_ex_stage_alu_adder_n4, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_alu_adder_n2, B => 
                           dp_ex_stage_alu_adder_n7, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n32, B => 
                           dp_ex_stage_alu_adder_B_xor_12_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Logic1_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_RCA1_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U9 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_3_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5,
                           B1 => dp_ex_stage_alu_adder_carries_3_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_3_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n13
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U8 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_0_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_0_port
                           , B2 => dp_ex_stage_alu_adder_carries_3_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n10);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U7 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n10, ZN => 
                           dp_ex_stage_alu_adder_out_12_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U6 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n13, ZN => 
                           dp_ex_stage_alu_adder_out_15_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U5 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_1_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_1_port
                           , B2 => dp_ex_stage_alu_adder_carries_3_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n11);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U4 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out0_2_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_rca_out1_2_port
                           , B2 => dp_ex_stage_alu_adder_carries_3_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n12);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n11, ZN => 
                           dp_ex_stage_alu_adder_out_13_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n12, ZN => 
                           dp_ex_stage_alu_adder_out_14_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_3_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_3_Mux_n5);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Logic0_port <= '0';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Logic1_port <= '1';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_19_port, B => 
                           dp_ex_stage_alu_adder_n6, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_18_port, B => 
                           dp_ex_stage_alu_adder_B_xor_18_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_17_port, B => 
                           dp_ex_stage_alu_adder_B_xor_17_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n38, B => 
                           dp_ex_stage_alu_adder_B_xor_16_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Logic0_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA0_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_19_port, B => 
                           dp_ex_stage_alu_adder_n6, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_18_port, B => 
                           dp_ex_stage_alu_adder_B_xor_18_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_17_port, B => 
                           dp_ex_stage_alu_adder_B_xor_17_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n38, B => 
                           dp_ex_stage_alu_adder_B_xor_16_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Logic1_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_RCA1_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U9 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_4_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U8 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_0_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5,
                           B1 => dp_ex_stage_alu_adder_carries_4_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_0_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n10
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U7 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_1_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_1_port
                           , B2 => dp_ex_stage_alu_adder_carries_4_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n11);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U6 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_2_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5,
                           B1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_2_port
                           , B2 => dp_ex_stage_alu_adder_carries_4_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n12);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U5 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out0_3_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n5,
                           B1 => dp_ex_stage_alu_adder_carries_4_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_rca_out1_3_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n13
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U4 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n10, ZN => 
                           dp_ex_stage_alu_adder_out_16_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n11, ZN => 
                           dp_ex_stage_alu_adder_out_17_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n12, ZN => 
                           dp_ex_stage_alu_adder_out_18_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_4_Mux_n13, ZN => 
                           dp_ex_stage_alu_adder_out_19_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Logic0_port <= '0';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Logic1_port <= '1';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_23_port, B => 
                           dp_ex_stage_alu_adder_n1, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_alu_n240, B => 
                           dp_ex_stage_alu_adder_B_xor_22_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_alu_n238, B => 
                           dp_ex_stage_alu_adder_B_xor_21_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n25, B => 
                           dp_ex_stage_alu_adder_B_xor_20_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Logic0_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA0_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_23_port, B => 
                           dp_ex_stage_alu_adder_n1, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_alu_n240, B => 
                           dp_ex_stage_alu_adder_B_xor_22_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_alu_n238, B => 
                           dp_ex_stage_alu_adder_B_xor_21_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n25, B => 
                           dp_ex_stage_alu_adder_B_xor_20_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Logic1_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_RCA1_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U10 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n1, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_0_port
                           , B1 => dp_ex_stage_alu_adder_carries_5_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_0_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n11
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U9 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n11, ZN => 
                           dp_ex_stage_alu_adder_out_20_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U8 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n14, ZN => 
                           dp_ex_stage_alu_adder_out_23_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U7 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_5_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n10);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U6 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_3_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n10
                           , B1 => dp_ex_stage_alu_adder_carries_5_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_3_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n14
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U5 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_2_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n1,
                           B1 => dp_ex_stage_alu_adder_carries_5_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_2_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n13
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U4 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n10, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out0_1_port
                           , B1 => dp_ex_stage_alu_adder_carries_5_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_rca_out1_1_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n12
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n13, ZN => 
                           dp_ex_stage_alu_adder_out_22_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n12, ZN => 
                           dp_ex_stage_alu_adder_out_21_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_5_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_5_Mux_n1);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Logic0_port <= '0';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Logic1_port <= '1';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_27_port, B => 
                           dp_ex_stage_alu_adder_B_xor_27_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_26_port, B => 
                           dp_ex_stage_alu_adder_B_xor_26_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_25_port, B => 
                           dp_ex_stage_alu_adder_B_xor_25_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_24_port, B => 
                           dp_ex_stage_alu_adder_B_xor_24_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Logic0_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA0_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U6 : NAND3_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n2, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n3, A3 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n4, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_3_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U5 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_B_xor_26_port, A2 => 
                           dp_ex_stage_muxA_out_26_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n4);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U4 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_port, 
                           A2 => dp_ex_stage_muxA_out_26_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n3);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U3 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_port, 
                           A2 => dp_ex_stage_alu_adder_B_xor_26_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n2);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U2 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_port, B 
                           => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n1, Z 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_U1 : XOR2_X1 port map( A => 
                           dp_ex_stage_alu_adder_B_xor_26_port, B => 
                           dp_ex_stage_muxA_out_26_port, Z => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_n1);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_27_port, B => 
                           dp_ex_stage_alu_adder_B_xor_27_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_25_port, B => 
                           dp_ex_stage_alu_adder_B_xor_25_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_24_port, B => 
                           dp_ex_stage_alu_adder_B_xor_24_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Logic1_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_RCA1_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U10 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n1, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_3_port
                           , B1 => dp_ex_stage_alu_adder_carries_6_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_3_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n14
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U9 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_2_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n1,
                           B1 => dp_ex_stage_alu_adder_carries_6_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_2_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n13
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U8 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_6_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n10);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U7 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_1_port
                           , A2 => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n10
                           , B1 => dp_ex_stage_alu_adder_carries_6_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_1_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n12
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U6 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n10, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out0_0_port
                           , B1 => dp_ex_stage_alu_adder_carries_6_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_rca_out1_0_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n11
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U5 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n13, ZN => 
                           dp_ex_stage_alu_adder_out_26_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U4 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n11, ZN => 
                           dp_ex_stage_alu_adder_out_24_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n14, ZN => 
                           dp_ex_stage_alu_adder_out_27_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n12, ZN => 
                           dp_ex_stage_alu_adder_out_25_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_6_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_6_Mux_n1);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Logic0_port <= '0';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Logic1_port <= '1';
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_31_port, B => 
                           dp_ex_stage_alu_adder_B_xor_31_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_30_port, B => 
                           dp_ex_stage_alu_adder_B_xor_30_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_29_port, B => 
                           dp_ex_stage_alu_adder_B_xor_29_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n247, B => 
                           dp_ex_stage_alu_adder_B_xor_28_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Logic0_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA0_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_U1_3 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_31_port, B => 
                           dp_ex_stage_alu_adder_B_xor_31_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_3_port, 
                           CO => dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_Co, 
                           S => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_3_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_U1_2 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_30_port, B => 
                           dp_ex_stage_alu_adder_B_xor_30_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_2_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_3_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_2_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_U1_1 : FA_X1 
                           port map( A => dp_ex_stage_muxA_out_29_port, B => 
                           dp_ex_stage_alu_adder_B_xor_29_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_1_port, 
                           CO => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_2_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_1_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_U1_0 : FA_X1 
                           port map( A => dp_ex_stage_alu_n247, B => 
                           dp_ex_stage_alu_adder_B_xor_28_port, CI => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Logic1_port, CO
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_RCA1_add_1_root_add_27_2_carry_1_port, S 
                           => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_0_port
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U10 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n14, ZN => 
                           dp_ex_stage_alu_adder_out_31_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U9 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_7_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n10);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U8 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n1, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_3_port
                           , B1 => dp_ex_stage_alu_adder_carries_7_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_3_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n14
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U7 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n10, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_0_port
                           , B1 => dp_ex_stage_alu_adder_carries_7_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_0_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n11
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U6 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n10, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_1_port
                           , B1 => dp_ex_stage_alu_adder_carries_7_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_1_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n12
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U5 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n1, A2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out0_2_port
                           , B1 => dp_ex_stage_alu_adder_carries_7_port, B2 => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_rca_out1_2_port
                           , ZN => dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n13
                           );
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U4 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n12, ZN => 
                           dp_ex_stage_alu_adder_out_29_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n11, ZN => 
                           dp_ex_stage_alu_adder_out_28_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U2 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n13, ZN => 
                           dp_ex_stage_alu_adder_out_30_port);
   dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_U1 : INV_X1 port map( A => 
                           dp_ex_stage_alu_adder_carries_7_port, ZN => 
                           dp_ex_stage_alu_adder_SumGen_CS_Bn_7_Mux_n1);
   dp_ex_stage_alu_shifter_U150 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N207, A2 => 
                           dp_ex_stage_alu_shifter_n115, B1 => 
                           dp_ex_stage_alu_shifter_N110_port, B2 => 
                           dp_ex_stage_alu_shifter_n112, C1 => 
                           dp_ex_stage_alu_shifter_N142, C2 => 
                           dp_ex_stage_alu_shifter_n109, ZN => 
                           dp_ex_stage_alu_shifter_n36);
   dp_ex_stage_alu_shifter_U149 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n33, A2 => 
                           dp_ex_stage_alu_shifter_n34, ZN => 
                           dp_ex_stage_alu_shifter_out_6_port);
   dp_ex_stage_alu_shifter_U148 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n37, A2 => 
                           dp_ex_stage_alu_shifter_n38, ZN => 
                           dp_ex_stage_alu_shifter_out_4_port);
   dp_ex_stage_alu_shifter_U147 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n35, A2 => 
                           dp_ex_stage_alu_shifter_n36, ZN => 
                           dp_ex_stage_alu_shifter_out_5_port);
   dp_ex_stage_alu_shifter_U146 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N213, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N116_port, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N148, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n86);
   dp_ex_stage_alu_shifter_U145 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N208, A2 => 
                           dp_ex_stage_alu_shifter_n115, B1 => 
                           dp_ex_stage_alu_shifter_N111_port, B2 => 
                           dp_ex_stage_alu_shifter_n112, C1 => 
                           dp_ex_stage_alu_shifter_N143, C2 => 
                           dp_ex_stage_alu_shifter_n109, ZN => 
                           dp_ex_stage_alu_shifter_n34);
   dp_ex_stage_alu_shifter_U144 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N206, A2 => 
                           dp_ex_stage_alu_shifter_n115, B1 => 
                           dp_ex_stage_alu_shifter_N109_port, B2 => 
                           dp_ex_stage_alu_shifter_n112, C1 => 
                           dp_ex_stage_alu_shifter_N141, C2 => 
                           dp_ex_stage_alu_shifter_n109, ZN => 
                           dp_ex_stage_alu_shifter_n38);
   dp_ex_stage_alu_shifter_U143 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N205, A2 => 
                           dp_ex_stage_alu_shifter_n115, B1 => 
                           dp_ex_stage_alu_shifter_N108_port, B2 => 
                           dp_ex_stage_alu_shifter_n112, C1 => 
                           dp_ex_stage_alu_shifter_N140, C2 => 
                           dp_ex_stage_alu_shifter_n109, ZN => 
                           dp_ex_stage_alu_shifter_n40);
   dp_ex_stage_alu_shifter_U142 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n39, A2 => 
                           dp_ex_stage_alu_shifter_n40, ZN => 
                           dp_ex_stage_alu_shifter_out_3_port);
   dp_ex_stage_alu_shifter_U141 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N219, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N122, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N154, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n74);
   dp_ex_stage_alu_shifter_U140 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n73, A2 => 
                           dp_ex_stage_alu_shifter_n74, ZN => 
                           dp_ex_stage_alu_shifter_out_17_port);
   dp_ex_stage_alu_shifter_U139 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N203, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N106_port, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N138, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n68);
   dp_ex_stage_alu_shifter_U138 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n67, A2 => 
                           dp_ex_stage_alu_shifter_n68, ZN => 
                           dp_ex_stage_alu_shifter_out_1_port);
   dp_ex_stage_alu_shifter_U137 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n90, A2 => 
                           dp_ex_stage_alu_shifter_n89, ZN => 
                           dp_ex_stage_alu_shifter_out_0_port);
   dp_ex_stage_alu_shifter_U136 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n45, A2 => 
                           dp_ex_stage_alu_shifter_n46, ZN => 
                           dp_ex_stage_alu_shifter_out_2_port);
   dp_ex_stage_alu_shifter_U135 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N218, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N121, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N153, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n76);
   dp_ex_stage_alu_shifter_U134 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n75, A2 => 
                           dp_ex_stage_alu_shifter_n76, ZN => 
                           dp_ex_stage_alu_shifter_out_16_port);
   dp_ex_stage_alu_shifter_U133 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N221, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N124, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N156, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n70);
   dp_ex_stage_alu_shifter_U132 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n69, A2 => 
                           dp_ex_stage_alu_shifter_n70, ZN => 
                           dp_ex_stage_alu_shifter_out_19_port);
   dp_ex_stage_alu_shifter_U131 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n83, A2 => 
                           dp_ex_stage_alu_shifter_n84, ZN => 
                           dp_ex_stage_alu_shifter_out_12_port);
   dp_ex_stage_alu_shifter_U130 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N212, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N115_port, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N147, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n88);
   dp_ex_stage_alu_shifter_U129 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n87, A2 => 
                           dp_ex_stage_alu_shifter_n88, ZN => 
                           dp_ex_stage_alu_shifter_out_10_port);
   dp_ex_stage_alu_shifter_U128 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N210, A2 => 
                           dp_ex_stage_alu_shifter_n115, B1 => 
                           dp_ex_stage_alu_shifter_N113_port, B2 => 
                           dp_ex_stage_alu_shifter_n112, C1 => 
                           dp_ex_stage_alu_shifter_N145, C2 => 
                           dp_ex_stage_alu_shifter_n109, ZN => 
                           dp_ex_stage_alu_shifter_n30);
   dp_ex_stage_alu_shifter_U127 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n29, A2 => 
                           dp_ex_stage_alu_shifter_n30, ZN => 
                           dp_ex_stage_alu_shifter_out_8_port);
   dp_ex_stage_alu_shifter_U126 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N211, A2 => 
                           dp_ex_stage_alu_shifter_n115, B1 => 
                           dp_ex_stage_alu_shifter_N114_port, B2 => 
                           dp_ex_stage_alu_shifter_n112, C1 => 
                           dp_ex_stage_alu_shifter_N146, C2 => 
                           dp_ex_stage_alu_shifter_n109, ZN => 
                           dp_ex_stage_alu_shifter_n22);
   dp_ex_stage_alu_shifter_U125 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n21, A2 => 
                           dp_ex_stage_alu_shifter_n22, ZN => 
                           dp_ex_stage_alu_shifter_out_9_port);
   dp_ex_stage_alu_shifter_U124 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N220, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N123, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N155, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n72);
   dp_ex_stage_alu_shifter_U123 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n71, A2 => 
                           dp_ex_stage_alu_shifter_n72, ZN => 
                           dp_ex_stage_alu_shifter_out_18_port);
   dp_ex_stage_alu_shifter_U122 : NOR2_X1 port map( A1 => dp_ex_stage_alu_n208,
                           A2 => dp_ex_stage_alu_Logic1_port, ZN => 
                           dp_ex_stage_alu_shifter_n28);
   dp_ex_stage_alu_shifter_U121 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n118, A2 => 
                           dp_ex_stage_alu_Logic1_port, ZN => 
                           dp_ex_stage_alu_shifter_n26);
   dp_ex_stage_alu_shifter_U120 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shift_arith_i, A2 => 
                           dp_ex_stage_alu_Logic1_port, ZN => 
                           dp_ex_stage_alu_shifter_n91);
   dp_ex_stage_alu_shifter_U119 : INV_X1 port map( A => 
                           dp_ex_stage_alu_Logic1_port, ZN => 
                           dp_ex_stage_alu_shifter_n117);
   dp_ex_stage_alu_shifter_U118 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n117, A2 => 
                           dp_ex_stage_alu_shift_arith_i, ZN => 
                           dp_ex_stage_alu_shifter_n92);
   dp_ex_stage_alu_shifter_U117 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n26, Z => 
                           dp_ex_stage_alu_shifter_n106);
   dp_ex_stage_alu_shifter_U116 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n28, Z => 
                           dp_ex_stage_alu_shifter_n100);
   dp_ex_stage_alu_shifter_U115 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n26, Z => 
                           dp_ex_stage_alu_shifter_n104);
   dp_ex_stage_alu_shifter_U114 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n26, Z => 
                           dp_ex_stage_alu_shifter_n105);
   dp_ex_stage_alu_shifter_U113 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n28, Z => 
                           dp_ex_stage_alu_shifter_n98);
   dp_ex_stage_alu_shifter_U112 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n28, Z => 
                           dp_ex_stage_alu_shifter_n99);
   dp_ex_stage_alu_shifter_U111 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n91, A2 => 
                           dp_ex_stage_alu_shifter_n118, ZN => 
                           dp_ex_stage_alu_shifter_n25);
   dp_ex_stage_alu_shifter_U110 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n92, A2 => 
                           dp_ex_stage_alu_shifter_n118, ZN => 
                           dp_ex_stage_alu_shifter_n24);
   dp_ex_stage_alu_shifter_U109 : AND2_X1 port map( A1 => dp_ex_stage_alu_n208,
                           A2 => dp_ex_stage_alu_shifter_n91, ZN => 
                           dp_ex_stage_alu_shifter_n27);
   dp_ex_stage_alu_shifter_U108 : AND2_X1 port map( A1 => dp_ex_stage_alu_n208,
                           A2 => dp_ex_stage_alu_shifter_n92, ZN => 
                           dp_ex_stage_alu_shifter_n23);
   dp_ex_stage_alu_shifter_U107 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N229, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N132, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N164, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n52);
   dp_ex_stage_alu_shifter_U106 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N54_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N249, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N22_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n77);
   dp_ex_stage_alu_shifter_U105 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n77, A2 => 
                           dp_ex_stage_alu_shifter_n78, ZN => 
                           dp_ex_stage_alu_shifter_out_15_port);
   dp_ex_stage_alu_shifter_U104 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N59_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N254, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N27_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n65);
   dp_ex_stage_alu_shifter_U103 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n65, A2 => 
                           dp_ex_stage_alu_shifter_n66, ZN => 
                           dp_ex_stage_alu_shifter_out_20_port);
   dp_ex_stage_alu_shifter_U102 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N62_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N257, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N30_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n59);
   dp_ex_stage_alu_shifter_U101 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n59, A2 => 
                           dp_ex_stage_alu_shifter_n60, ZN => 
                           dp_ex_stage_alu_shifter_out_23_port);
   dp_ex_stage_alu_shifter_U100 : INV_X1 port map( A => dp_ex_stage_alu_n208, 
                           ZN => dp_ex_stage_alu_shifter_n118);
   dp_ex_stage_alu_shifter_U99 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n85, A2 => 
                           dp_ex_stage_alu_shifter_n86, ZN => 
                           dp_ex_stage_alu_shifter_out_11_port);
   dp_ex_stage_alu_shifter_U98 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n25, Z => 
                           dp_ex_stage_alu_shifter_n109);
   dp_ex_stage_alu_shifter_U97 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n24, Z => 
                           dp_ex_stage_alu_shifter_n112);
   dp_ex_stage_alu_shifter_U96 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n23, Z => 
                           dp_ex_stage_alu_shifter_n115);
   dp_ex_stage_alu_shifter_U95 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n23, Z => 
                           dp_ex_stage_alu_shifter_n113);
   dp_ex_stage_alu_shifter_U94 : CLKBUF_X3 port map( A => 
                           dp_ex_stage_muxB_out_4_port, Z => 
                           dp_ex_stage_alu_shifter_n116);
   dp_ex_stage_alu_shifter_U93 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N69_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N264, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N37_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n43);
   dp_ex_stage_alu_shifter_U92 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n43, A2 => 
                           dp_ex_stage_alu_shifter_n44, ZN => 
                           dp_ex_stage_alu_shifter_out_30_port);
   dp_ex_stage_alu_shifter_U91 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N70_port, A2 => 
                           dp_ex_stage_alu_shifter_n106, B1 => 
                           dp_ex_stage_alu_shifter_N265, B2 => 
                           dp_ex_stage_alu_shifter_n103, C1 => 
                           dp_ex_stage_alu_shifter_N38_port, C2 => 
                           dp_ex_stage_alu_shifter_n100, ZN => 
                           dp_ex_stage_alu_shifter_n41);
   dp_ex_stage_alu_shifter_U90 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n41, A2 => 
                           dp_ex_stage_alu_shifter_n42, ZN => 
                           dp_ex_stage_alu_shifter_out_31_port);
   dp_ex_stage_alu_shifter_U89 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N67_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N262, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N35_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n49);
   dp_ex_stage_alu_shifter_U88 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n49, A2 => 
                           dp_ex_stage_alu_shifter_n50, ZN => 
                           dp_ex_stage_alu_shifter_out_28_port);
   dp_ex_stage_alu_shifter_U87 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N68_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N263, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N36_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n47);
   dp_ex_stage_alu_shifter_U86 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n47, A2 => 
                           dp_ex_stage_alu_shifter_n48, ZN => 
                           dp_ex_stage_alu_shifter_out_29_port);
   dp_ex_stage_alu_shifter_U85 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N63_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N258, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N31_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n57);
   dp_ex_stage_alu_shifter_U84 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n57, A2 => 
                           dp_ex_stage_alu_shifter_n58, ZN => 
                           dp_ex_stage_alu_shifter_out_24_port);
   dp_ex_stage_alu_shifter_U83 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N61_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N256, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N29_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n61);
   dp_ex_stage_alu_shifter_U82 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n61, A2 => 
                           dp_ex_stage_alu_shifter_n62, ZN => 
                           dp_ex_stage_alu_shifter_out_22_port);
   dp_ex_stage_alu_shifter_U81 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N65_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N260, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N33_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n53);
   dp_ex_stage_alu_shifter_U80 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n53, A2 => 
                           dp_ex_stage_alu_shifter_n54, ZN => 
                           dp_ex_stage_alu_shifter_out_26_port);
   dp_ex_stage_alu_shifter_U79 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N64_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N259, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N32_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n55);
   dp_ex_stage_alu_shifter_U78 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n55, A2 => 
                           dp_ex_stage_alu_shifter_n56, ZN => 
                           dp_ex_stage_alu_shifter_out_25_port);
   dp_ex_stage_alu_shifter_U77 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N60_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N255, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N28_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n63);
   dp_ex_stage_alu_shifter_U76 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n63, A2 => 
                           dp_ex_stage_alu_shifter_n64, ZN => 
                           dp_ex_stage_alu_shifter_out_21_port);
   dp_ex_stage_alu_shifter_U75 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N66_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N261, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N34_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n51);
   dp_ex_stage_alu_shifter_U74 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n51, A2 => 
                           dp_ex_stage_alu_shifter_n52, ZN => 
                           dp_ex_stage_alu_shifter_out_27_port);
   dp_ex_stage_alu_shifter_U73 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n31, A2 => 
                           dp_ex_stage_alu_shifter_n32, ZN => 
                           dp_ex_stage_alu_shifter_out_7_port);
   dp_ex_stage_alu_shifter_U72 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N52_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N247, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N20_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n81);
   dp_ex_stage_alu_shifter_U71 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n81, A2 => 
                           dp_ex_stage_alu_shifter_n82, ZN => 
                           dp_ex_stage_alu_shifter_out_13_port);
   dp_ex_stage_alu_shifter_U70 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N53_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N248, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N21_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n79);
   dp_ex_stage_alu_shifter_U69 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n79, A2 => 
                           dp_ex_stage_alu_shifter_n80, ZN => 
                           dp_ex_stage_alu_shifter_out_14_port);
   dp_ex_stage_alu_shifter_U68 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n27, Z => 
                           dp_ex_stage_alu_shifter_n103);
   dp_ex_stage_alu_shifter_U67 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n23, Z => 
                           dp_ex_stage_alu_shifter_n114);
   dp_ex_stage_alu_shifter_U66 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n24, Z => 
                           dp_ex_stage_alu_shifter_n111);
   dp_ex_stage_alu_shifter_U65 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n27, Z => 
                           dp_ex_stage_alu_shifter_n101);
   dp_ex_stage_alu_shifter_U64 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n27, Z => 
                           dp_ex_stage_alu_shifter_n102);
   dp_ex_stage_alu_shifter_U63 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N51_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N246, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N19_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n83);
   dp_ex_stage_alu_shifter_U62 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N49_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N244, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N17_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n87);
   dp_ex_stage_alu_shifter_U61 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N56_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N251, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N24_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n73);
   dp_ex_stage_alu_shifter_U60 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N57_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N252, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N25_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n71);
   dp_ex_stage_alu_shifter_U59 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N58_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N253, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N26_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n69);
   dp_ex_stage_alu_shifter_U58 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N55_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N250, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N23_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n75);
   dp_ex_stage_alu_shifter_U57 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N39_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N234, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N7_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n89);
   dp_ex_stage_alu_shifter_U56 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N40_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N235, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N8_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n67);
   dp_ex_stage_alu_shifter_U55 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N41_port, A2 => 
                           dp_ex_stage_alu_shifter_n105, B1 => 
                           dp_ex_stage_alu_shifter_N236, B2 => 
                           dp_ex_stage_alu_shifter_n102, C1 => 
                           dp_ex_stage_alu_shifter_N9_port, C2 => 
                           dp_ex_stage_alu_shifter_n99, ZN => 
                           dp_ex_stage_alu_shifter_n45);
   dp_ex_stage_alu_shifter_U54 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N45_port, A2 => 
                           dp_ex_stage_alu_shifter_n106, B1 => 
                           dp_ex_stage_alu_shifter_N240, B2 => 
                           dp_ex_stage_alu_shifter_n103, C1 => 
                           dp_ex_stage_alu_shifter_N13_port, C2 => 
                           dp_ex_stage_alu_shifter_n100, ZN => 
                           dp_ex_stage_alu_shifter_n33);
   dp_ex_stage_alu_shifter_U53 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N48_port, A2 => 
                           dp_ex_stage_alu_shifter_n106, B1 => 
                           dp_ex_stage_alu_shifter_N243, B2 => 
                           dp_ex_stage_alu_shifter_n103, C1 => 
                           dp_ex_stage_alu_shifter_N16_port, C2 => 
                           dp_ex_stage_alu_shifter_n100, ZN => 
                           dp_ex_stage_alu_shifter_n21);
   dp_ex_stage_alu_shifter_U52 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N47_port, A2 => 
                           dp_ex_stage_alu_shifter_n106, B1 => 
                           dp_ex_stage_alu_shifter_N242, B2 => 
                           dp_ex_stage_alu_shifter_n103, C1 => 
                           dp_ex_stage_alu_shifter_N15_port, C2 => 
                           dp_ex_stage_alu_shifter_n100, ZN => 
                           dp_ex_stage_alu_shifter_n29);
   dp_ex_stage_alu_shifter_U51 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N42_port, A2 => 
                           dp_ex_stage_alu_shifter_n106, B1 => 
                           dp_ex_stage_alu_shifter_N237, B2 => 
                           dp_ex_stage_alu_shifter_n103, C1 => 
                           dp_ex_stage_alu_shifter_N10_port, C2 => 
                           dp_ex_stage_alu_shifter_n100, ZN => 
                           dp_ex_stage_alu_shifter_n39);
   dp_ex_stage_alu_shifter_U50 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N43_port, A2 => 
                           dp_ex_stage_alu_shifter_n106, B1 => 
                           dp_ex_stage_alu_shifter_N238, B2 => 
                           dp_ex_stage_alu_shifter_n103, C1 => 
                           dp_ex_stage_alu_shifter_N11_port, C2 => 
                           dp_ex_stage_alu_shifter_n100, ZN => 
                           dp_ex_stage_alu_shifter_n37);
   dp_ex_stage_alu_shifter_U49 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N44_port, A2 => 
                           dp_ex_stage_alu_shifter_n106, B1 => 
                           dp_ex_stage_alu_shifter_N239, B2 => 
                           dp_ex_stage_alu_shifter_n103, C1 => 
                           dp_ex_stage_alu_shifter_N12_port, C2 => 
                           dp_ex_stage_alu_shifter_n100, ZN => 
                           dp_ex_stage_alu_shifter_n35);
   dp_ex_stage_alu_shifter_U48 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N50_port, A2 => 
                           dp_ex_stage_alu_shifter_n104, B1 => 
                           dp_ex_stage_alu_shifter_N245, B2 => 
                           dp_ex_stage_alu_shifter_n101, C1 => 
                           dp_ex_stage_alu_shifter_N18_port, C2 => 
                           dp_ex_stage_alu_shifter_n98, ZN => 
                           dp_ex_stage_alu_shifter_n85);
   dp_ex_stage_alu_shifter_U47 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N46_port, A2 => 
                           dp_ex_stage_alu_shifter_n106, B1 => 
                           dp_ex_stage_alu_shifter_N241, B2 => 
                           dp_ex_stage_alu_shifter_n103, C1 => 
                           dp_ex_stage_alu_shifter_N14_port, C2 => 
                           dp_ex_stage_alu_shifter_n100, ZN => 
                           dp_ex_stage_alu_shifter_n31);
   dp_ex_stage_alu_shifter_U46 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N217, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N120, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N152, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n78);
   dp_ex_stage_alu_shifter_U45 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N215, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N118_port, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N150, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n82);
   dp_ex_stage_alu_shifter_U44 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N216, A2 => 
                           dp_ex_stage_alu_shifter_n113, B1 => 
                           dp_ex_stage_alu_shifter_N119, B2 => 
                           dp_ex_stage_alu_shifter_n110, C1 => 
                           dp_ex_stage_alu_shifter_N151, C2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n80);
   dp_ex_stage_alu_shifter_U43 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N230, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N133, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N165, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n50);
   dp_ex_stage_alu_shifter_U42 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N232, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N135, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N167, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n44);
   dp_ex_stage_alu_shifter_U41 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N231, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N134, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N166, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n48);
   dp_ex_stage_alu_shifter_U40 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N233, A2 => 
                           dp_ex_stage_alu_shifter_n115, B1 => 
                           dp_ex_stage_alu_shifter_N136, B2 => 
                           dp_ex_stage_alu_shifter_n112, C1 => 
                           dp_ex_stage_alu_shifter_N168, C2 => 
                           dp_ex_stage_alu_shifter_n109, ZN => 
                           dp_ex_stage_alu_shifter_n42);
   dp_ex_stage_alu_shifter_U39 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N209, A2 => 
                           dp_ex_stage_alu_shifter_n115, B1 => 
                           dp_ex_stage_alu_shifter_N112_port, B2 => 
                           dp_ex_stage_alu_shifter_n112, C1 => 
                           dp_ex_stage_alu_shifter_N144, C2 => 
                           dp_ex_stage_alu_shifter_n109, ZN => 
                           dp_ex_stage_alu_shifter_n32);
   dp_ex_stage_alu_shifter_U38 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N227, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N130, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N162, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n56);
   dp_ex_stage_alu_shifter_U37 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N228, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N131, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N163, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n54);
   dp_ex_stage_alu_shifter_U36 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N224, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N127, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N159, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n62);
   dp_ex_stage_alu_shifter_U35 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N223, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N126, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N158, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n64);
   dp_ex_stage_alu_shifter_U34 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N225, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N128, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N160, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n60);
   dp_ex_stage_alu_shifter_U33 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N226, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N129, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N161, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n58);
   dp_ex_stage_alu_shifter_U32 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N222, A2 => 
                           dp_ex_stage_alu_shifter_n114, B1 => 
                           dp_ex_stage_alu_shifter_N125, B2 => 
                           dp_ex_stage_alu_shifter_n111, C1 => 
                           dp_ex_stage_alu_shifter_N157, C2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n66);
   dp_ex_stage_alu_shifter_U31 : AND3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n95, A2 => 
                           dp_ex_stage_alu_shifter_n96, A3 => 
                           dp_ex_stage_alu_shifter_n97, ZN => 
                           dp_ex_stage_alu_shifter_n84);
   dp_ex_stage_alu_shifter_U30 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N149, A2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n97);
   dp_ex_stage_alu_shifter_U29 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N117_port, A2 => 
                           dp_ex_stage_alu_shifter_n110, ZN => 
                           dp_ex_stage_alu_shifter_n96);
   dp_ex_stage_alu_shifter_U28 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N214, A2 => 
                           dp_ex_stage_alu_shifter_n113, ZN => 
                           dp_ex_stage_alu_shifter_n95);
   dp_ex_stage_alu_shifter_U27 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_muxA_out_24_port, Z => 
                           dp_ex_stage_alu_shifter_n94);
   dp_ex_stage_alu_shifter_U26 : NOR3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n93, A2 => 
                           dp_ex_stage_alu_shifter_n20, A3 => 
                           dp_ex_stage_alu_shifter_n19, ZN => 
                           dp_ex_stage_alu_shifter_n90);
   dp_ex_stage_alu_shifter_U25 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N137, A2 => 
                           dp_ex_stage_alu_shifter_n107, ZN => 
                           dp_ex_stage_alu_shifter_n93);
   dp_ex_stage_alu_shifter_U24 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N105_port, A2 => 
                           dp_ex_stage_alu_shifter_n110, ZN => 
                           dp_ex_stage_alu_shifter_n20);
   dp_ex_stage_alu_shifter_U23 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N202, A2 => 
                           dp_ex_stage_alu_shifter_n113, ZN => 
                           dp_ex_stage_alu_shifter_n19);
   dp_ex_stage_alu_shifter_U22 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_muxA_out_27_port, Z => 
                           dp_ex_stage_alu_shifter_n12);
   dp_ex_stage_alu_shifter_U21 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_muxA_out_26_port, Z => 
                           dp_ex_stage_alu_shifter_n11);
   dp_ex_stage_alu_shifter_U20 : AND3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n8, A2 => 
                           dp_ex_stage_alu_shifter_n9, A3 => 
                           dp_ex_stage_alu_shifter_n10, ZN => 
                           dp_ex_stage_alu_shifter_n46);
   dp_ex_stage_alu_shifter_U19 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N139, A2 => 
                           dp_ex_stage_alu_shifter_n108, ZN => 
                           dp_ex_stage_alu_shifter_n10);
   dp_ex_stage_alu_shifter_U18 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N107_port, A2 => 
                           dp_ex_stage_alu_shifter_n111, ZN => 
                           dp_ex_stage_alu_shifter_n9);
   dp_ex_stage_alu_shifter_U17 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N204, A2 => 
                           dp_ex_stage_alu_shifter_n114, ZN => 
                           dp_ex_stage_alu_shifter_n8);
   dp_ex_stage_alu_shifter_U16 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n6, ZN => 
                           dp_ex_stage_alu_shifter_n7);
   dp_ex_stage_alu_shifter_U15 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_25_port, ZN => 
                           dp_ex_stage_alu_shifter_n6);
   dp_ex_stage_alu_shifter_U14 : INV_X2 port map( A => 
                           dp_ex_stage_alu_shifter_n4, ZN => 
                           dp_ex_stage_alu_shifter_n5);
   dp_ex_stage_alu_shifter_U13 : INV_X1 port map( A => dp_ex_stage_alu_n46, ZN 
                           => dp_ex_stage_alu_shifter_n4);
   dp_ex_stage_alu_shifter_U10 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n2, ZN => 
                           dp_ex_stage_alu_shifter_n3);
   dp_ex_stage_alu_shifter_U9 : INV_X1 port map( A => dp_ex_stage_alu_n45, ZN 
                           => dp_ex_stage_alu_shifter_n2);
   dp_ex_stage_alu_shifter_U8 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_muxA_out_31_port, Z => 
                           dp_ex_stage_alu_shifter_n1);
   dp_ex_stage_alu_shifter_U7 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n25, Z => 
                           dp_ex_stage_alu_shifter_n107);
   dp_ex_stage_alu_shifter_U6 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n24, Z => 
                           dp_ex_stage_alu_shifter_n110);
   dp_ex_stage_alu_shifter_U5 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n25, Z => 
                           dp_ex_stage_alu_shifter_n108);
   dp_ex_stage_alu_shifter_n18 <= '0';
   dp_ex_stage_alu_shifter_n17 <= '0';
   dp_ex_stage_alu_shifter_n16 <= '0';
   dp_ex_stage_alu_shifter_n15 <= '0';
   dp_ex_stage_alu_shifter_n14 <= '0';
   dp_ex_stage_alu_shifter_n13 <= '0';
   dp_ex_stage_alu_shifter_sll_48_U59 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N202, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n4, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_0_port);
   dp_ex_stage_alu_shifter_sll_48_U58 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_0_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n8, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_0_port);
   dp_ex_stage_alu_shifter_sll_48_U57 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_1_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n8, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_1_port);
   dp_ex_stage_alu_shifter_sll_48_U56 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_0_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n12, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_0_port);
   dp_ex_stage_alu_shifter_sll_48_U55 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_1_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n12, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_1_port);
   dp_ex_stage_alu_shifter_sll_48_U54 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_2_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n12, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_2_port);
   dp_ex_stage_alu_shifter_sll_48_U53 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_3_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n12, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_3_port);
   dp_ex_stage_alu_shifter_sll_48_U52 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_0_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n34);
   dp_ex_stage_alu_shifter_sll_48_U51 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_1_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n33);
   dp_ex_stage_alu_shifter_sll_48_U50 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_2_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n32);
   dp_ex_stage_alu_shifter_sll_48_U49 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_3_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n31);
   dp_ex_stage_alu_shifter_sll_48_U48 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_4_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n30);
   dp_ex_stage_alu_shifter_sll_48_U47 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_5_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n29);
   dp_ex_stage_alu_shifter_sll_48_U46 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_6_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n28);
   dp_ex_stage_alu_shifter_sll_48_U45 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_7_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n27);
   dp_ex_stage_alu_shifter_sll_48_U44 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_n17, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n34, ZN => 
                           dp_ex_stage_alu_shifter_N234);
   dp_ex_stage_alu_shifter_sll_48_U43 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_10_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_N244);
   dp_ex_stage_alu_shifter_sll_48_U42 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_11_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_N245);
   dp_ex_stage_alu_shifter_sll_48_U41 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_12_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_N246);
   dp_ex_stage_alu_shifter_sll_48_U40 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_13_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_N247);
   dp_ex_stage_alu_shifter_sll_48_U39 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_14_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_N248);
   dp_ex_stage_alu_shifter_sll_48_U38 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_15_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_N249);
   dp_ex_stage_alu_shifter_sll_48_U37 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_n17, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n33, ZN => 
                           dp_ex_stage_alu_shifter_N235);
   dp_ex_stage_alu_shifter_sll_48_U36 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_n17, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n32, ZN => 
                           dp_ex_stage_alu_shifter_N236);
   dp_ex_stage_alu_shifter_sll_48_U35 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_n17, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n31, ZN => 
                           dp_ex_stage_alu_shifter_N237);
   dp_ex_stage_alu_shifter_sll_48_U34 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_n17, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n30, ZN => 
                           dp_ex_stage_alu_shifter_N238);
   dp_ex_stage_alu_shifter_sll_48_U33 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_n17, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n29, ZN => 
                           dp_ex_stage_alu_shifter_N239);
   dp_ex_stage_alu_shifter_sll_48_U32 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_n17, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n28, ZN => 
                           dp_ex_stage_alu_shifter_N240);
   dp_ex_stage_alu_shifter_sll_48_U31 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_n17, A2 => 
                           dp_ex_stage_alu_shifter_sll_48_n27, ZN => 
                           dp_ex_stage_alu_shifter_N241);
   dp_ex_stage_alu_shifter_sll_48_U30 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_8_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_N242);
   dp_ex_stage_alu_shifter_sll_48_U29 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_9_port, A2 
                           => dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_N243);
   dp_ex_stage_alu_shifter_sll_48_U28 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n18);
   dp_ex_stage_alu_shifter_sll_48_U27 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n14);
   dp_ex_stage_alu_shifter_sll_48_U26 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n15, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n13);
   dp_ex_stage_alu_shifter_sll_48_U25 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n49, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n12);
   dp_ex_stage_alu_shifter_sll_48_U24 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n12, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n11);
   dp_ex_stage_alu_shifter_sll_48_U23 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n8, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n7);
   dp_ex_stage_alu_shifter_sll_48_U22 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n4, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n3);
   dp_ex_stage_alu_shifter_sll_48_U21 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n5, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n8);
   dp_ex_stage_alu_shifter_sll_48_U20 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n15);
   dp_ex_stage_alu_shifter_sll_48_U19 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n45, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n4);
   dp_ex_stage_alu_shifter_sll_48_U18 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n4, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n2);
   dp_ex_stage_alu_shifter_sll_48_U17 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n4, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n1);
   dp_ex_stage_alu_shifter_sll_48_U16 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n33, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n23);
   dp_ex_stage_alu_shifter_sll_48_U15 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n32, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n21);
   dp_ex_stage_alu_shifter_sll_48_U14 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n31, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n25);
   dp_ex_stage_alu_shifter_sll_48_U13 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n34, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n19);
   dp_ex_stage_alu_shifter_sll_48_U12 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n28, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n22);
   dp_ex_stage_alu_shifter_sll_48_U11 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n27, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n26);
   dp_ex_stage_alu_shifter_sll_48_U10 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n29, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n24);
   dp_ex_stage_alu_shifter_sll_48_U9 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n30, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n20);
   dp_ex_stage_alu_shifter_sll_48_U8 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n8, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n6);
   dp_ex_stage_alu_shifter_sll_48_U7 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n8, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n5);
   dp_ex_stage_alu_shifter_sll_48_U6 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n12, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n10);
   dp_ex_stage_alu_shifter_sll_48_U5 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n12, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n9);
   dp_ex_stage_alu_shifter_sll_48_U4 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n17);
   dp_ex_stage_alu_shifter_sll_48_U3 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_n18, ZN => 
                           dp_ex_stage_alu_shifter_sll_48_n16);
   dp_ex_stage_alu_shifter_sll_48_M1_0_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n76, B => 
                           dp_ex_stage_alu_shifter_N202, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_1_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n44, B => dp_ex_stage_alu_n76, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_2_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n69, B => dp_ex_stage_alu_n44, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_3_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n52, B => dp_ex_stage_alu_n69, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_4_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n70, B => dp_ex_stage_alu_n52, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_5_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n78, B => dp_ex_stage_alu_n70, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_6_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n34, B => dp_ex_stage_alu_n78, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_7_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n71, B => dp_ex_stage_alu_n34, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_8_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n72, B => dp_ex_stage_alu_n71, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_9_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n74, B => dp_ex_stage_alu_n72, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_10_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n33, B => dp_ex_stage_alu_n74, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_11_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_12_port, B => 
                           dp_ex_stage_alu_n33, S => 
                           dp_ex_stage_alu_shifter_sll_48_n1, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_12_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n231, B => 
                           dp_ex_stage_muxA_out_12_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_13_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_14_port, B => 
                           dp_ex_stage_alu_n231, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_14_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n29, B => 
                           dp_ex_stage_muxA_out_14_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_15_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n38, B => dp_ex_stage_alu_n29, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_16_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_17_port, B => 
                           dp_ex_stage_alu_n38, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_17_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_18_port, B => 
                           dp_ex_stage_muxA_out_17_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_18_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_19_port, B => 
                           dp_ex_stage_muxA_out_18_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_19_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_20_port, B => 
                           dp_ex_stage_muxA_out_19_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_20_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_21_port, B => 
                           dp_ex_stage_muxA_out_20_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_21_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n240, B => 
                           dp_ex_stage_muxA_out_21_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_22_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_23_port, B => 
                           dp_ex_stage_alu_n240, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_23_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n94, B => 
                           dp_ex_stage_muxA_out_23_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n2, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_24_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n7, B => 
                           dp_ex_stage_alu_shifter_n94, S => 
                           dp_ex_stage_alu_shifter_sll_48_n3, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_25_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n11, B => 
                           dp_ex_stage_alu_shifter_n7, S => 
                           dp_ex_stage_alu_shifter_sll_48_n3, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_26_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n12, B => 
                           dp_ex_stage_alu_shifter_n11, S => 
                           dp_ex_stage_alu_shifter_sll_48_n3, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_27_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n1, B => dp_ex_stage_alu_shifter_n12
                           , S => dp_ex_stage_alu_shifter_sll_48_n3, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_28_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_29_port, B => 
                           dp_ex_stage_alu_n1, S => 
                           dp_ex_stage_alu_shifter_sll_48_n3, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_29_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_30_port, B => 
                           dp_ex_stage_muxA_out_29_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n3, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_30_port);
   dp_ex_stage_alu_shifter_sll_48_M1_0_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_31_port, B => 
                           dp_ex_stage_muxA_out_30_port, S => 
                           dp_ex_stage_alu_shifter_sll_48_n3, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_31_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_2_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_0_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_2_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_3_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_1_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_3_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_4_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_2_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_4_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_5_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_3_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_5_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_6_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_4_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_6_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_7_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_5_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_7_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_8_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_6_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_8_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_9_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_7_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_9_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_10_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_8_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_10_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_11_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_9_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_11_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_12_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_10_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_12_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_13_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_11_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n5, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_13_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_14_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_12_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_14_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_15_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_13_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_15_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_16_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_14_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_16_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_17_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_15_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_17_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_18_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_16_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_18_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_19_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_17_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_19_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_20_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_18_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_20_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_21_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_19_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_21_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_22_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_20_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_22_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_23_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_21_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_23_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_24_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_22_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_24_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_25_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_23_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n6, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_25_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_26_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_24_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n7, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_26_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_27_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_25_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n7, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_27_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_28_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_26_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n7, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_28_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_29_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_27_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n7, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_29_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_30_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_28_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n7, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_30_port);
   dp_ex_stage_alu_shifter_sll_48_M1_1_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_1_31_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_1_29_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n7, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_31_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_4_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_0_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_4_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_5_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_1_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_5_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_6_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_2_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_6_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_7_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_3_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_7_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_8_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_4_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_8_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_9_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_5_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_9_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_10_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_6_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_10_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_11_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_7_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_11_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_12_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_8_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_12_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_13_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_9_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_13_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_14_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_10_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_14_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_15_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_11_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n9, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_15_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_16_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_12_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_16_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_17_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_13_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_17_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_18_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_14_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_18_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_19_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_15_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_19_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_20_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_16_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_20_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_21_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_17_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_21_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_22_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_18_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_22_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_23_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_19_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_23_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_24_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_20_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_24_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_25_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_21_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_25_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_26_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_22_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_26_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_27_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_23_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n10, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_27_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_28_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_24_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n11, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_28_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_29_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_25_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n11, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_29_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_30_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_26_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n11, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_30_port);
   dp_ex_stage_alu_shifter_sll_48_M1_2_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_2_31_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_2_27_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n11, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_31_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_8_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_0_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_8_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_9_port, B =>
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_1_port, S =>
                           dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_9_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_10_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_2_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_10_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_11_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_3_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_11_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_12_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_4_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_12_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_13_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_5_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_13_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_14_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_6_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_14_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_15_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_7_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_15_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_16_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_8_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_16_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_17_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_9_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_17_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_18_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_10_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_18_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_19_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_11_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n13, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_19_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_20_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_12_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_20_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_21_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_13_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_21_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_22_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_14_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_22_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_23_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_15_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_23_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_24_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_16_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_24_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_25_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_17_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_25_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_26_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_18_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_26_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_27_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_19_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_27_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_28_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_20_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_28_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_29_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_21_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_29_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_30_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_22_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_30_port);
   dp_ex_stage_alu_shifter_sll_48_M1_3_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_3_31_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_3_23_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n14, Z => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_31_port);
   dp_ex_stage_alu_shifter_sll_48_M1_4_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_16_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_n19, S => 
                           dp_ex_stage_alu_shifter_sll_48_n17, Z => 
                           dp_ex_stage_alu_shifter_N250);
   dp_ex_stage_alu_shifter_sll_48_M1_4_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_17_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_n23, S => 
                           dp_ex_stage_alu_shifter_sll_48_n17, Z => 
                           dp_ex_stage_alu_shifter_N251);
   dp_ex_stage_alu_shifter_sll_48_M1_4_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_18_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_n21, S => 
                           dp_ex_stage_alu_shifter_sll_48_n17, Z => 
                           dp_ex_stage_alu_shifter_N252);
   dp_ex_stage_alu_shifter_sll_48_M1_4_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_19_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_n25, S => 
                           dp_ex_stage_alu_shifter_sll_48_n17, Z => 
                           dp_ex_stage_alu_shifter_N253);
   dp_ex_stage_alu_shifter_sll_48_M1_4_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_20_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_n20, S => 
                           dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N254);
   dp_ex_stage_alu_shifter_sll_48_M1_4_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_21_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_n24, S => 
                           dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N255);
   dp_ex_stage_alu_shifter_sll_48_M1_4_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_22_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_n22, S => 
                           dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N256);
   dp_ex_stage_alu_shifter_sll_48_M1_4_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_23_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_n26, S => 
                           dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N257);
   dp_ex_stage_alu_shifter_sll_48_M1_4_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_24_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_4_8_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N258);
   dp_ex_stage_alu_shifter_sll_48_M1_4_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_25_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_4_9_port, S
                           => dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N259);
   dp_ex_stage_alu_shifter_sll_48_M1_4_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_26_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_4_10_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N260);
   dp_ex_stage_alu_shifter_sll_48_M1_4_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_27_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_4_11_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N261);
   dp_ex_stage_alu_shifter_sll_48_M1_4_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_28_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_4_12_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N262);
   dp_ex_stage_alu_shifter_sll_48_M1_4_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_29_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_4_13_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N263);
   dp_ex_stage_alu_shifter_sll_48_M1_4_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_30_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_4_14_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N264);
   dp_ex_stage_alu_shifter_sll_48_M1_4_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sll_48_ML_int_4_31_port, B 
                           => dp_ex_stage_alu_shifter_sll_48_ML_int_4_15_port, 
                           S => dp_ex_stage_alu_shifter_sll_48_n16, Z => 
                           dp_ex_stage_alu_shifter_N265);
   dp_ex_stage_alu_shifter_sla_46_U225 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n5, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n13, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n95);
   dp_ex_stage_alu_shifter_sla_46_U224 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n45, A2 => 
                           dp_ex_stage_alu_shifter_n5, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n96);
   dp_ex_stage_alu_shifter_sla_46_U223 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n13, A2 => 
                           dp_ex_stage_alu_shifter_n5, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n98);
   dp_ex_stage_alu_shifter_sla_46_U222 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_n45, A2 => 
                           dp_ex_stage_alu_shifter_n5, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n99);
   dp_ex_stage_alu_shifter_sla_46_U221 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n70, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_alu_n78, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n193);
   dp_ex_stage_alu_shifter_sla_46_U220 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n57, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n20, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, A => 
                           dp_ex_stage_alu_shifter_sla_46_n193, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n155);
   dp_ex_stage_alu_shifter_sla_46_U219 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n14, A2 => 
                           dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n133);
   dp_ex_stage_alu_shifter_sla_46_U218 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n72, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n9, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n24, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n12, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n192);
   dp_ex_stage_alu_shifter_sla_46_U217 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n3, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n22, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n21, A => 
                           dp_ex_stage_alu_shifter_sla_46_n192, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n154);
   dp_ex_stage_alu_shifter_sla_46_U216 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n31, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n14, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n137);
   dp_ex_stage_alu_shifter_sla_46_U215 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n31, A2 => 
                           dp_ex_stage_alu_shifter_N202, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n158);
   dp_ex_stage_alu_shifter_sla_46_U214 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n14, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n158, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n139);
   dp_ex_stage_alu_shifter_sla_46_U213 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n137, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n48, A => 
                           dp_ex_stage_alu_shifter_sla_46_n139, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n190);
   dp_ex_stage_alu_shifter_sla_46_U212 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n17, A2 => 
                           dp_ex_stage_alu_shifter_N202, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n80);
   dp_ex_stage_alu_shifter_sla_46_U211 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n17, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n125, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N212);
   dp_ex_stage_alu_shifter_sla_46_U210 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n9, B1 => 
                           dp_ex_stage_alu_n34, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n12, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n189);
   dp_ex_stage_alu_shifter_sla_46_U209 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n3, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n58, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n6, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n57, A => 
                           dp_ex_stage_alu_shifter_sla_46_n189, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n151);
   dp_ex_stage_alu_shifter_sla_46_U208 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n24, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n9, B1 => 
                           dp_ex_stage_alu_n33, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n12, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n188);
   dp_ex_stage_alu_shifter_sla_46_U207 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n3, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n23, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n6, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n22, A => 
                           dp_ex_stage_alu_shifter_sla_46_n188, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n149);
   dp_ex_stage_alu_shifter_sla_46_U206 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n9, A2 => 
                           dp_ex_stage_alu_n44, B1 => dp_ex_stage_alu_n69, B2 
                           => dp_ex_stage_alu_shifter_sla_46_n12, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n187);
   dp_ex_stage_alu_shifter_sla_46_U205 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n56, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n3, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n55, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, A => 
                           dp_ex_stage_alu_shifter_sla_46_n187, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n150);
   dp_ex_stage_alu_shifter_sla_46_U204 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n137, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n150, A => 
                           dp_ex_stage_alu_shifter_sla_46_n139, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n186);
   dp_ex_stage_alu_shifter_sla_46_U203 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n17, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n120, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N213);
   dp_ex_stage_alu_shifter_sla_46_U202 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n34, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_alu_n71, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n12, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n185);
   dp_ex_stage_alu_shifter_sla_46_U201 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n3, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n60, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n6, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n58, A => 
                           dp_ex_stage_alu_shifter_sla_46_n185, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n145);
   dp_ex_stage_alu_shifter_sla_46_U200 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n33, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_muxA_out_12_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n184);
   dp_ex_stage_alu_shifter_sla_46_U199 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n25, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n6, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n23, A => 
                           dp_ex_stage_alu_shifter_sla_46_n184, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n143);
   dp_ex_stage_alu_shifter_sla_46_U198 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n9, A2 => 
                           dp_ex_stage_alu_n69, B1 => dp_ex_stage_alu_n52, B2 
                           => dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n183);
   dp_ex_stage_alu_shifter_sla_46_U197 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n19, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n56, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, A => 
                           dp_ex_stage_alu_shifter_sla_46_n183, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n144);
   dp_ex_stage_alu_shifter_sla_46_U196 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n137, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n144, A => 
                           dp_ex_stage_alu_shifter_sla_46_n139, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n182);
   dp_ex_stage_alu_shifter_sla_46_U195 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n17, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n113, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N214);
   dp_ex_stage_alu_shifter_sla_46_U194 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_N202, B => 
                           dp_ex_stage_alu_n76, S => 
                           dp_ex_stage_alu_shifter_sla_46_n10, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n138);
   dp_ex_stage_alu_shifter_sla_46_U193 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n49, A2 => dp_ex_stage_alu_n31, ZN 
                           => dp_ex_stage_alu_shifter_sla_46_n174);
   dp_ex_stage_alu_shifter_sla_46_U192 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n52, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_alu_n70, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n181);
   dp_ex_stage_alu_shifter_sla_46_U191 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n20, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n6, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n19, A => 
                           dp_ex_stage_alu_shifter_sla_46_n181, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n132);
   dp_ex_stage_alu_shifter_sla_46_U190 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n71, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_alu_n72, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n180);
   dp_ex_stage_alu_shifter_sla_46_U189 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n21, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n60, A => 
                           dp_ex_stage_alu_shifter_sla_46_n180, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n134);
   dp_ex_stage_alu_shifter_sla_46_U188 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_12_port, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n28, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n179);
   dp_ex_stage_alu_shifter_sla_46_U187 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n26, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n25, A => 
                           dp_ex_stage_alu_shifter_sla_46_n179, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n131);
   dp_ex_stage_alu_shifter_sla_46_U186 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n134, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n131, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n178);
   dp_ex_stage_alu_shifter_sla_46_U185 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n138, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n174, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n132, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n137, A => 
                           dp_ex_stage_alu_shifter_sla_46_n59, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n107);
   dp_ex_stage_alu_shifter_sla_46_U184 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n16, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n107, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N215);
   dp_ex_stage_alu_shifter_sla_46_U183 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n28, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n30, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n177);
   dp_ex_stage_alu_shifter_sla_46_U182 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n27, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n26, A => 
                           dp_ex_stage_alu_shifter_sla_46_n177, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n127);
   dp_ex_stage_alu_shifter_sla_46_U181 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n174, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n48, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n137, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n155, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n176);
   dp_ex_stage_alu_shifter_sla_46_U180 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n154, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n127, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n47, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n100);
   dp_ex_stage_alu_shifter_sla_46_U179 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n16, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n100, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N216);
   dp_ex_stage_alu_shifter_sla_46_U178 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n30, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_alu_n29, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n175);
   dp_ex_stage_alu_shifter_sla_46_U177 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n29, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n27, A => 
                           dp_ex_stage_alu_shifter_sla_46_n175, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n122);
   dp_ex_stage_alu_shifter_sla_46_U176 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n174, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n150, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n137, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n151, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n173);
   dp_ex_stage_alu_shifter_sla_46_U175 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n149, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n122, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n54, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n88);
   dp_ex_stage_alu_shifter_sla_46_U174 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n16, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n88, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N217);
   dp_ex_stage_alu_shifter_sla_46_U173 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n87);
   dp_ex_stage_alu_shifter_sla_46_U172 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n29, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n33, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n172);
   dp_ex_stage_alu_shifter_sla_46_U171 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n31, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n29, A => 
                           dp_ex_stage_alu_shifter_sla_46_n172, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n115);
   dp_ex_stage_alu_shifter_sla_46_U170 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n31, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n171);
   dp_ex_stage_alu_shifter_sla_46_U169 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n171, A2 => 
                           dp_ex_stage_alu_n49, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n90);
   dp_ex_stage_alu_shifter_sla_46_U168 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n144, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n145, A => 
                           dp_ex_stage_alu_shifter_sla_46_n53, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n170);
   dp_ex_stage_alu_shifter_sla_46_U167 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n61, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n87, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n62, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, A => 
                           dp_ex_stage_alu_shifter_sla_46_n170, ZN => 
                           dp_ex_stage_alu_shifter_N218);
   dp_ex_stage_alu_shifter_sla_46_U166 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n33, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n35, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n169);
   dp_ex_stage_alu_shifter_sla_46_U165 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n32, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n31, A => 
                           dp_ex_stage_alu_shifter_sla_46_n169, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n109);
   dp_ex_stage_alu_shifter_sla_46_U164 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n55, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n14, A => 
                           dp_ex_stage_alu_shifter_sla_46_n158, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n161);
   dp_ex_stage_alu_shifter_sla_46_U163 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n138, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n161, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n163);
   dp_ex_stage_alu_shifter_sla_46_U162 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n131, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n134, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n132, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n168);
   dp_ex_stage_alu_shifter_sla_46_U161 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n63, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n163, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n168, ZN => 
                           dp_ex_stage_alu_shifter_N219);
   dp_ex_stage_alu_shifter_sla_46_U160 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n35, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_muxA_out_18_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n167);
   dp_ex_stage_alu_shifter_sla_46_U159 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n34, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n32, A => 
                           dp_ex_stage_alu_shifter_sla_46_n167, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n102);
   dp_ex_stage_alu_shifter_sla_46_U158 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n48, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n161, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n106);
   dp_ex_stage_alu_shifter_sla_46_U157 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n127, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n154, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n155, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n166);
   dp_ex_stage_alu_shifter_sla_46_U156 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n64, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n106, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n166, ZN => 
                           dp_ex_stage_alu_shifter_N220);
   dp_ex_stage_alu_shifter_sla_46_U155 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_18_port, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_muxA_out_19_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n165);
   dp_ex_stage_alu_shifter_sla_46_U154 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n36, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n34, A => 
                           dp_ex_stage_alu_shifter_sla_46_n165, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n91);
   dp_ex_stage_alu_shifter_sla_46_U153 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n150, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n161, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n86);
   dp_ex_stage_alu_shifter_sla_46_U152 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n122, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n149, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n151, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n164);
   dp_ex_stage_alu_shifter_sla_46_U151 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n65, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n86, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n164, ZN => 
                           dp_ex_stage_alu_shifter_N221);
   dp_ex_stage_alu_shifter_sla_46_U150 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n16, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n163, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N203);
   dp_ex_stage_alu_shifter_sla_46_U149 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_19_port, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_muxA_out_20_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n162);
   dp_ex_stage_alu_shifter_sla_46_U148 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n37, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n36, A => 
                           dp_ex_stage_alu_shifter_sla_46_n162, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n117);
   dp_ex_stage_alu_shifter_sla_46_U147 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n144, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n161, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n85);
   dp_ex_stage_alu_shifter_sla_46_U146 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n115, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n143, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n145, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n160);
   dp_ex_stage_alu_shifter_sla_46_U145 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n66, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n85, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n160, ZN => 
                           dp_ex_stage_alu_shifter_N222);
   dp_ex_stage_alu_shifter_sla_46_U144 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_20_port, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_muxA_out_21_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n159);
   dp_ex_stage_alu_shifter_sla_46_U143 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n69, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n37, A => 
                           dp_ex_stage_alu_shifter_sla_46_n159, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n111);
   dp_ex_stage_alu_shifter_sla_46_U142 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n109, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n131, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n134, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n157);
   dp_ex_stage_alu_shifter_sla_46_U141 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n67, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n84, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n157, ZN => 
                           dp_ex_stage_alu_shifter_N223);
   dp_ex_stage_alu_shifter_sla_46_U140 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_21_port, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_alu_n240, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n156);
   dp_ex_stage_alu_shifter_sla_46_U139 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n71, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n69, A => 
                           dp_ex_stage_alu_shifter_sla_46_n156, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n104);
   dp_ex_stage_alu_shifter_sla_46_U138 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n102, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n127, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n154, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n153);
   dp_ex_stage_alu_shifter_sla_46_U137 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n68, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n83, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n153, ZN => 
                           dp_ex_stage_alu_shifter_N224);
   dp_ex_stage_alu_shifter_sla_46_U136 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n240, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_muxA_out_23_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n152);
   dp_ex_stage_alu_shifter_sla_46_U135 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n38, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n71, A => 
                           dp_ex_stage_alu_shifter_sla_46_n152, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n94);
   dp_ex_stage_alu_shifter_sla_46_U134 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n91, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n122, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n149, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n148);
   dp_ex_stage_alu_shifter_sla_46_U133 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n70, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n82, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n148, ZN => 
                           dp_ex_stage_alu_shifter_N225);
   dp_ex_stage_alu_shifter_sla_46_U132 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_23_port, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_alu_shifter_n94, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n147);
   dp_ex_stage_alu_shifter_sla_46_U131 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n39, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n38, A => 
                           dp_ex_stage_alu_shifter_sla_46_n147, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n146);
   dp_ex_stage_alu_shifter_sla_46_U130 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n117, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n115, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n143, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n142);
   dp_ex_stage_alu_shifter_sla_46_U129 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n72, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n81, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n142, ZN => 
                           dp_ex_stage_alu_shifter_N226);
   dp_ex_stage_alu_shifter_sla_46_U128 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n94, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_alu_shifter_n7, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n141);
   dp_ex_stage_alu_shifter_sla_46_U127 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n40, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n39, A => 
                           dp_ex_stage_alu_shifter_sla_46_n141, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n140);
   dp_ex_stage_alu_shifter_sla_46_U126 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n137, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n138, A => 
                           dp_ex_stage_alu_shifter_sla_46_n139, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n136);
   dp_ex_stage_alu_shifter_sla_46_U125 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n132, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n134, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n51, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n79);
   dp_ex_stage_alu_shifter_sla_46_U124 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n111, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n109, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n131, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n130);
   dp_ex_stage_alu_shifter_sla_46_U123 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n73, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n79, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n130, ZN => 
                           dp_ex_stage_alu_shifter_N227);
   dp_ex_stage_alu_shifter_sla_46_U122 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n7, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_alu_shifter_n11, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n129);
   dp_ex_stage_alu_shifter_sla_46_U121 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n41, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n40, A => 
                           dp_ex_stage_alu_shifter_sla_46_n129, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n128);
   dp_ex_stage_alu_shifter_sla_46_U120 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n104, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n102, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n127, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n126);
   dp_ex_stage_alu_shifter_sla_46_U119 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n74, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n125, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n126, ZN => 
                           dp_ex_stage_alu_shifter_N228);
   dp_ex_stage_alu_shifter_sla_46_U118 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n11, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_alu_shifter_n12, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n124);
   dp_ex_stage_alu_shifter_sla_46_U117 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n42, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n41, A => 
                           dp_ex_stage_alu_shifter_sla_46_n124, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n123);
   dp_ex_stage_alu_shifter_sla_46_U116 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n78, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n94, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n91, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n122, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n121);
   dp_ex_stage_alu_shifter_sla_46_U115 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n75, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n119, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n120, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n121, ZN => 
                           dp_ex_stage_alu_shifter_N229);
   dp_ex_stage_alu_shifter_sla_46_U114 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_n12, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_alu_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n118);
   dp_ex_stage_alu_shifter_sla_46_U113 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n43, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n42, A => 
                           dp_ex_stage_alu_shifter_sla_46_n118, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n116);
   dp_ex_stage_alu_shifter_sla_46_U112 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n115, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n77, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n116, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n117, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n114);
   dp_ex_stage_alu_shifter_sla_46_U111 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n72, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n87, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n113, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n114, ZN => 
                           dp_ex_stage_alu_shifter_N230);
   dp_ex_stage_alu_shifter_sla_46_U110 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n1, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_muxA_out_29_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n112);
   dp_ex_stage_alu_shifter_sla_46_U109 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n44, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n43, A => 
                           dp_ex_stage_alu_shifter_sla_46_n112, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n110);
   dp_ex_stage_alu_shifter_sla_46_U108 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n109, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n77, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n110, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n111, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n108);
   dp_ex_stage_alu_shifter_sla_46_U107 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n73, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n87, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n107, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n108, ZN => 
                           dp_ex_stage_alu_shifter_N231);
   dp_ex_stage_alu_shifter_sla_46_U106 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n16, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n106, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N204);
   dp_ex_stage_alu_shifter_sla_46_U105 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_29_port, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n7, B1 => 
                           dp_ex_stage_muxA_out_30_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n105);
   dp_ex_stage_alu_shifter_sla_46_U104 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n1, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n45, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n4, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n44, A => 
                           dp_ex_stage_alu_shifter_sla_46_n105, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n103);
   dp_ex_stage_alu_shifter_sla_46_U103 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n102, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n77, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n103, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n104, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n101);
   dp_ex_stage_alu_shifter_sla_46_U102 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n74, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n87, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n100, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n101, ZN => 
                           dp_ex_stage_alu_shifter_N232);
   dp_ex_stage_alu_shifter_sla_46_U101 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_30_port, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n8, B1 => 
                           dp_ex_stage_muxA_out_31_port, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n97);
   dp_ex_stage_alu_shifter_sla_46_U100 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n2, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n76, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n5, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n45, A => 
                           dp_ex_stage_alu_shifter_sla_46_n97, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n92);
   dp_ex_stage_alu_shifter_sla_46_U99 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n90, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n91, B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n77, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n92, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n93, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n94, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n89);
   dp_ex_stage_alu_shifter_sla_46_U98 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n75, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n87, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n88, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, A => 
                           dp_ex_stage_alu_shifter_sla_46_n89, ZN => 
                           dp_ex_stage_alu_shifter_N233);
   dp_ex_stage_alu_shifter_sla_46_U97 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n16, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n86, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N205);
   dp_ex_stage_alu_shifter_sla_46_U96 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n16, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n85, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N206);
   dp_ex_stage_alu_shifter_sla_46_U95 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n15, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n84, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N207);
   dp_ex_stage_alu_shifter_sla_46_U94 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n15, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n83, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N208);
   dp_ex_stage_alu_shifter_sla_46_U93 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n15, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n82, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N209);
   dp_ex_stage_alu_shifter_sla_46_U92 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n15, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n81, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N210);
   dp_ex_stage_alu_shifter_sla_46_U91 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n15, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n79, A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_N211);
   dp_ex_stage_alu_shifter_sla_46_U90 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n1, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n45);
   dp_ex_stage_alu_shifter_sla_46_U89 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n12, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n44);
   dp_ex_stage_alu_shifter_sla_46_U88 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n11, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n43);
   dp_ex_stage_alu_shifter_sla_46_U87 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n7, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n42);
   dp_ex_stage_alu_shifter_sla_46_U86 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n94, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n41);
   dp_ex_stage_alu_shifter_sla_46_U85 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_23_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n40);
   dp_ex_stage_alu_shifter_sla_46_U84 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n240, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n39);
   dp_ex_stage_alu_shifter_sla_46_U83 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_21_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n38);
   dp_ex_stage_alu_shifter_sla_46_U82 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_18_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n37);
   dp_ex_stage_alu_shifter_sla_46_U81 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_17_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n36);
   dp_ex_stage_alu_shifter_sla_46_U80 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n36, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n35);
   dp_ex_stage_alu_shifter_sla_46_U79 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n38, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n34);
   dp_ex_stage_alu_shifter_sla_46_U78 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n34, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n33);
   dp_ex_stage_alu_shifter_sla_46_U77 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n29, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n32);
   dp_ex_stage_alu_shifter_sla_46_U76 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_14_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n31);
   dp_ex_stage_alu_shifter_sla_46_U75 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n31, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n30);
   dp_ex_stage_alu_shifter_sla_46_U74 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n231, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n29);
   dp_ex_stage_alu_shifter_sla_46_U73 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n29, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n28);
   dp_ex_stage_alu_shifter_sla_46_U72 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_12_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n27);
   dp_ex_stage_alu_shifter_sla_46_U71 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n33, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n26);
   dp_ex_stage_alu_shifter_sla_46_U70 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n74, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n25);
   dp_ex_stage_alu_shifter_sla_46_U69 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n25, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n24);
   dp_ex_stage_alu_shifter_sla_46_U68 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n72, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n23);
   dp_ex_stage_alu_shifter_sla_46_U67 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n71, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n22);
   dp_ex_stage_alu_shifter_sla_46_U66 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n34, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n21);
   dp_ex_stage_alu_shifter_sla_46_U65 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n69, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n20);
   dp_ex_stage_alu_shifter_sla_46_U64 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n44, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n19);
   dp_ex_stage_alu_shifter_sla_46_U63 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n49, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n14);
   dp_ex_stage_alu_shifter_sla_46_U62 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n45, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n13);
   dp_ex_stage_alu_shifter_sla_46_U61 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n52, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n57);
   dp_ex_stage_alu_shifter_sla_46_U60 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n78, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n60);
   dp_ex_stage_alu_shifter_sla_46_U59 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_N202, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n55);
   dp_ex_stage_alu_shifter_sla_46_U58 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n70, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n58);
   dp_ex_stage_alu_shifter_sla_46_U57 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n76, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n56);
   dp_ex_stage_alu_shifter_sla_46_U56 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n191, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n48);
   dp_ex_stage_alu_shifter_sla_46_U55 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_20_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n71);
   dp_ex_stage_alu_shifter_sla_46_U54 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_19_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n69);
   dp_ex_stage_alu_shifter_sla_46_U53 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_29_port, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n76);
   dp_ex_stage_alu_shifter_sla_46_U52 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n96, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n6);
   dp_ex_stage_alu_shifter_sla_46_U51 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n99, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n12);
   dp_ex_stage_alu_shifter_sla_46_U50 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n117, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n66);
   dp_ex_stage_alu_shifter_sla_46_U49 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n111, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n67);
   dp_ex_stage_alu_shifter_sla_46_U48 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n178, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n59);
   dp_ex_stage_alu_shifter_sla_46_U47 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n158, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n52);
   dp_ex_stage_alu_shifter_sla_46_U46 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n91, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n65);
   dp_ex_stage_alu_shifter_sla_46_U45 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n96, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n5);
   dp_ex_stage_alu_shifter_sla_46_U44 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n96, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n4);
   dp_ex_stage_alu_shifter_sla_46_U43 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n171, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n14, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n93);
   dp_ex_stage_alu_shifter_sla_46_U42 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n99, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n11);
   dp_ex_stage_alu_shifter_sla_46_U41 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n99, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n10);
   dp_ex_stage_alu_shifter_sla_46_U40 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n80, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n53);
   dp_ex_stage_alu_shifter_sla_46_U39 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n136, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n51);
   dp_ex_stage_alu_shifter_sla_46_U38 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n182, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n50);
   dp_ex_stage_alu_shifter_sla_46_U37 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n190, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n46);
   dp_ex_stage_alu_shifter_sla_46_U36 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n186, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n49);
   dp_ex_stage_alu_shifter_sla_46_U35 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n173, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n54);
   dp_ex_stage_alu_shifter_sla_46_U34 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n176, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n47);
   dp_ex_stage_alu_shifter_sla_46_U33 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n146, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n72);
   dp_ex_stage_alu_shifter_sla_46_U32 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n140, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n73);
   dp_ex_stage_alu_shifter_sla_46_U31 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n128, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n74);
   dp_ex_stage_alu_shifter_sla_46_U30 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n123, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n75);
   dp_ex_stage_alu_shifter_sla_46_U29 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n95, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n3);
   dp_ex_stage_alu_shifter_sla_46_U28 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n104, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n68);
   dp_ex_stage_alu_shifter_sla_46_U27 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n94, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n70);
   dp_ex_stage_alu_shifter_sla_46_U26 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n143, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n61);
   dp_ex_stage_alu_shifter_sla_46_U25 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n115, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n62);
   dp_ex_stage_alu_shifter_sla_46_U24 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n98, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n9);
   dp_ex_stage_alu_shifter_sla_46_U23 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n109, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n63);
   dp_ex_stage_alu_shifter_sla_46_U22 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n102, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n64);
   dp_ex_stage_alu_shifter_sla_46_U21 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n15);
   dp_ex_stage_alu_shifter_sla_46_U20 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n95, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n1);
   dp_ex_stage_alu_shifter_sla_46_U19 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n95, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n2);
   dp_ex_stage_alu_shifter_sla_46_U18 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n98, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n8);
   dp_ex_stage_alu_shifter_sla_46_U17 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n98, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n7);
   dp_ex_stage_alu_shifter_sla_46_U16 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n119, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n77);
   dp_ex_stage_alu_shifter_sla_46_U15 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n87, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n78);
   dp_ex_stage_alu_shifter_sla_46_U14 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sla_46_n15, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n18);
   dp_ex_stage_alu_shifter_sla_46_U13 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n17);
   dp_ex_stage_alu_shifter_sla_46_U12 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_sla_46_n16);
   dp_ex_stage_alu_shifter_sla_46_U11 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n10, A2 => 
                           dp_ex_stage_alu_n44, B1 => dp_ex_stage_alu_n76, B2 
                           => dp_ex_stage_alu_shifter_sla_46_n9, C1 => 
                           dp_ex_stage_alu_shifter_N202, C2 => 
                           dp_ex_stage_alu_shifter_n5, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n191);
   dp_ex_stage_alu_shifter_sla_46_U10 : NOR2_X2 port map( A1 => 
                           dp_ex_stage_alu_n49, A2 => dp_ex_stage_alu_n31, ZN 
                           => dp_ex_stage_alu_shifter_sla_46_n135);
   dp_ex_stage_alu_shifter_sla_46_U9 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n150, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n151, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n52, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n82);
   dp_ex_stage_alu_shifter_sla_46_U8 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n151, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n149, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n49, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n120);
   dp_ex_stage_alu_shifter_sla_46_U7 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n155, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n154, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n46, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n125);
   dp_ex_stage_alu_shifter_sla_46_U6 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n145, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n143, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n50, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n113);
   dp_ex_stage_alu_shifter_sla_46_U5 : NAND2_X2 port map( A1 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A2 => 
                           dp_ex_stage_alu_shifter_sla_46_n18, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n119);
   dp_ex_stage_alu_shifter_sla_46_U4 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n138, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n132, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n52, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n84);
   dp_ex_stage_alu_shifter_sla_46_U3 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n48, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n155, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n52, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n83);
   dp_ex_stage_alu_shifter_sla_46_U2 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sla_46_n144, B2 => 
                           dp_ex_stage_alu_shifter_sla_46_n133, C1 => 
                           dp_ex_stage_alu_shifter_sla_46_n145, C2 => 
                           dp_ex_stage_alu_shifter_sla_46_n135, A => 
                           dp_ex_stage_alu_shifter_sla_46_n52, ZN => 
                           dp_ex_stage_alu_shifter_sla_46_n81);
   dp_ex_stage_alu_shifter_srl_41_U222 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n46, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n3, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n120);
   dp_ex_stage_alu_shifter_srl_41_U221 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n55, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n54, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n189);
   dp_ex_stage_alu_shifter_srl_41_U220 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n24, A2 => 
                           dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n137);
   dp_ex_stage_alu_shifter_srl_41_U219 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n114);
   dp_ex_stage_alu_shifter_srl_41_U218 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_23_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B1 => 
                           dp_ex_stage_alu_n240, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n188);
   dp_ex_stage_alu_shifter_srl_41_U217 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_17_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_n38, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n187);
   dp_ex_stage_alu_shifter_srl_41_U216 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n68, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n45, A => 
                           dp_ex_stage_alu_shifter_srl_41_n187, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n96);
   dp_ex_stage_alu_shifter_srl_41_U215 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n24, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n25, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n164);
   dp_ex_stage_alu_shifter_srl_41_U214 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n24, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n25, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n152);
   dp_ex_stage_alu_shifter_srl_41_U213 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_29_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n186);
   dp_ex_stage_alu_shifter_srl_41_U212 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n25, A2 => 
                           dp_ex_stage_alu_n49, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n140);
   dp_ex_stage_alu_shifter_srl_41_U211 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_25_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_muxA_out_24_port, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n185);
   dp_ex_stage_alu_shifter_srl_41_U210 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n51, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n50, A => 
                           dp_ex_stage_alu_shifter_srl_41_n185, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n138);
   dp_ex_stage_alu_shifter_srl_41_U209 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n152, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n134, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n140, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n138, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n184);
   dp_ex_stage_alu_shifter_srl_41_U208 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n97, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n96, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, A => 
                           dp_ex_stage_alu_shifter_srl_41_n70, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n154);
   dp_ex_stage_alu_shifter_srl_41_U207 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n25, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n28, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n181);
   dp_ex_stage_alu_shifter_srl_41_U206 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n231, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n37, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n183);
   dp_ex_stage_alu_shifter_srl_41_U205 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n42, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n40, A => 
                           dp_ex_stage_alu_shifter_srl_41_n183, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n95);
   dp_ex_stage_alu_shifter_srl_41_U204 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n76, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_shifter_N202, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n182);
   dp_ex_stage_alu_shifter_srl_41_U203 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n31, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n30, A => 
                           dp_ex_stage_alu_shifter_srl_41_n182, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n179);
   dp_ex_stage_alu_shifter_srl_41_U202 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n34, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n33, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n180);
   dp_ex_stage_alu_shifter_srl_41_U201 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n111, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n114, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n154, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n178, ZN => 
                           dp_ex_stage_alu_shifter_N137);
   dp_ex_stage_alu_shifter_srl_41_U200 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n36, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n35, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n177);
   dp_ex_stage_alu_shifter_srl_41_U199 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B2 => 
                           dp_ex_stage_alu_n231, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n37, A => 
                           dp_ex_stage_alu_shifter_srl_41_n177, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n130);
   dp_ex_stage_alu_shifter_srl_41_U198 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_27_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_muxA_out_26_port, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n176);
   dp_ex_stage_alu_shifter_srl_41_U197 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n74, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n52, A => 
                           dp_ex_stage_alu_shifter_srl_41_n176, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n142);
   dp_ex_stage_alu_shifter_srl_41_U196 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n75, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n53, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n126);
   dp_ex_stage_alu_shifter_srl_41_U195 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n142, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n126, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n135);
   dp_ex_stage_alu_shifter_srl_41_U194 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n41, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n39, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n175);
   dp_ex_stage_alu_shifter_srl_41_U193 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n44, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n43, A => 
                           dp_ex_stage_alu_shifter_srl_41_n175, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n106);
   dp_ex_stage_alu_shifter_srl_41_U192 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, A2 => 
                           dp_ex_stage_muxA_out_19_port, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, B2 => 
                           dp_ex_stage_muxA_out_18_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n174);
   dp_ex_stage_alu_shifter_srl_41_U191 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n46, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n69, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, A => 
                           dp_ex_stage_alu_shifter_srl_41_n174, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n107);
   dp_ex_stage_alu_shifter_srl_41_U190 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_23_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_n240, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n173);
   dp_ex_stage_alu_shifter_srl_41_U189 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n49, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n48, A => 
                           dp_ex_stage_alu_shifter_srl_41_n173, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n143);
   dp_ex_stage_alu_shifter_srl_41_U188 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n80, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n106, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n107, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n143, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n172);
   dp_ex_stage_alu_shifter_srl_41_U187 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n130, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n135, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n172, ZN => 
                           dp_ex_stage_alu_shifter_N147);
   dp_ex_stage_alu_shifter_srl_41_U186 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n38, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n41, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n171);
   dp_ex_stage_alu_shifter_srl_41_U185 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n45, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n44, A => 
                           dp_ex_stage_alu_shifter_srl_41_n171, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n101);
   dp_ex_stage_alu_shifter_srl_41_U184 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n38, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n36, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n170);
   dp_ex_stage_alu_shifter_srl_41_U183 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_24_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_muxA_out_23_port, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n169);
   dp_ex_stage_alu_shifter_srl_41_U182 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n50, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n49, A => 
                           dp_ex_stage_alu_shifter_srl_41_n169, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n141);
   dp_ex_stage_alu_shifter_srl_41_U181 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n240, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B1 => 
                           dp_ex_stage_muxA_out_21_port, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n168);
   dp_ex_stage_alu_shifter_srl_41_U180 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n69, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n68, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, A => 
                           dp_ex_stage_alu_shifter_srl_41_n168, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n102);
   dp_ex_stage_alu_shifter_srl_41_U179 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n1, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n19, B1 => 
                           dp_ex_stage_muxA_out_27_port, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n167);
   dp_ex_stage_alu_shifter_srl_41_U178 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n53, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n125);
   dp_ex_stage_alu_shifter_srl_41_U177 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n139, B => 
                           dp_ex_stage_alu_shifter_srl_41_n125, S => 
                           dp_ex_stage_alu_n49, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n150);
   dp_ex_stage_alu_shifter_srl_41_U176 : NOR3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A2 => 
                           dp_ex_stage_alu_n31, A3 => 
                           dp_ex_stage_alu_shifter_srl_41_n73, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n166);
   dp_ex_stage_alu_shifter_srl_41_U175 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n141, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n102, A => 
                           dp_ex_stage_alu_shifter_srl_41_n166, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n165);
   dp_ex_stage_alu_shifter_srl_41_U174 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n64, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n114, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n118, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, A => 
                           dp_ex_stage_alu_shifter_srl_41_n165, ZN => 
                           dp_ex_stage_alu_shifter_N148);
   dp_ex_stage_alu_shifter_srl_41_U173 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n164, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n156);
   dp_ex_stage_alu_shifter_srl_41_U172 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n96, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n80, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n95, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, A => 
                           dp_ex_stage_alu_shifter_srl_41_n2, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n163);
   dp_ex_stage_alu_shifter_srl_41_U171 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_18_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_muxA_out_17_port, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n162);
   dp_ex_stage_alu_shifter_srl_41_U170 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n69, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n68, A => 
                           dp_ex_stage_alu_shifter_srl_41_n162, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n89);
   dp_ex_stage_alu_shifter_srl_41_U169 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n39, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_n231, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n161);
   dp_ex_stage_alu_shifter_srl_41_U168 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n43, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n42, A => 
                           dp_ex_stage_alu_shifter_srl_41_n161, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n87);
   dp_ex_stage_alu_shifter_srl_41_U167 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_26_port, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_muxA_out_25_port, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n160);
   dp_ex_stage_alu_shifter_srl_41_U166 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n52, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n51, A => 
                           dp_ex_stage_alu_shifter_srl_41_n160, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n136);
   dp_ex_stage_alu_shifter_srl_41_U165 : OAI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n75, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n53, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n74, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n133);
   dp_ex_stage_alu_shifter_srl_41_U164 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n240, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_muxA_out_21_port, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n159);
   dp_ex_stage_alu_shifter_srl_41_U163 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n48, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n47, A => 
                           dp_ex_stage_alu_shifter_srl_41_n159, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n91);
   dp_ex_stage_alu_shifter_srl_41_U162 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n136, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n156, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n133, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n91, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n158);
   dp_ex_stage_alu_shifter_srl_41_U161 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n65, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n114, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n62, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, A => 
                           dp_ex_stage_alu_shifter_srl_41_n158, ZN => 
                           dp_ex_stage_alu_shifter_N150);
   dp_ex_stage_alu_shifter_srl_41_U160 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n142, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n156, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n126, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n143, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n157);
   dp_ex_stage_alu_shifter_srl_41_U159 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n66, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n114, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n63, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, A => 
                           dp_ex_stage_alu_shifter_srl_41_n157, ZN => 
                           dp_ex_stage_alu_shifter_N151);
   dp_ex_stage_alu_shifter_srl_41_U158 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n139, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n156, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n125, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n141, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n155);
   dp_ex_stage_alu_shifter_srl_41_U157 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n67, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n114, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n64, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, A => 
                           dp_ex_stage_alu_shifter_srl_41_n155, ZN => 
                           dp_ex_stage_alu_shifter_N152);
   dp_ex_stage_alu_shifter_srl_41_U156 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n28, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n154, ZN => 
                           dp_ex_stage_alu_shifter_N153);
   dp_ex_stage_alu_shifter_srl_41_U155 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n152, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n133, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n140, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n136, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n153);
   dp_ex_stage_alu_shifter_srl_41_U154 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n91, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n89, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, A => 
                           dp_ex_stage_alu_shifter_srl_41_n71, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n144);
   dp_ex_stage_alu_shifter_srl_41_U153 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n27, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n144, ZN => 
                           dp_ex_stage_alu_shifter_N154);
   dp_ex_stage_alu_shifter_srl_41_U152 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n152, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n126, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n140, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n142, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n151);
   dp_ex_stage_alu_shifter_srl_41_U151 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n143, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n107, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, A => 
                           dp_ex_stage_alu_shifter_srl_41_n72, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n127);
   dp_ex_stage_alu_shifter_srl_41_U150 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n27, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n127, ZN => 
                           dp_ex_stage_alu_shifter_N155);
   dp_ex_stage_alu_shifter_srl_41_U149 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n102, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n141, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n150, C2 => 
                           dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n115);
   dp_ex_stage_alu_shifter_srl_41_U148 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n27, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n115, ZN => 
                           dp_ex_stage_alu_shifter_N156);
   dp_ex_stage_alu_shifter_srl_41_U147 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n56, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n55, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n149);
   dp_ex_stage_alu_shifter_srl_41_U146 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n44, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_n76, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n148);
   dp_ex_stage_alu_shifter_srl_41_U145 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n54, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n31, A => 
                           dp_ex_stage_alu_shifter_srl_41_n148, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n146);
   dp_ex_stage_alu_shifter_srl_41_U144 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n35, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n34, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n147);
   dp_ex_stage_alu_shifter_srl_41_U143 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n37, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, C2 => 
                           dp_ex_stage_alu_n33, A => 
                           dp_ex_stage_alu_shifter_srl_41_n147, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n83);
   dp_ex_stage_alu_shifter_srl_41_U142 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n87, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n146, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n58, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n145);
   dp_ex_stage_alu_shifter_srl_41_U141 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n108, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n114, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n144, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n145, ZN => 
                           dp_ex_stage_alu_shifter_N138);
   dp_ex_stage_alu_shifter_srl_41_U140 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n27, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n112, ZN => 
                           dp_ex_stage_alu_shifter_N157);
   dp_ex_stage_alu_shifter_srl_41_U139 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n136, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n133, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n140, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n91, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n109);
   dp_ex_stage_alu_shifter_srl_41_U138 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n27, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n109, ZN => 
                           dp_ex_stage_alu_shifter_N158);
   dp_ex_stage_alu_shifter_srl_41_U137 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n142, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n126, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n140, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n143, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n104);
   dp_ex_stage_alu_shifter_srl_41_U136 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n26, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n104, ZN => 
                           dp_ex_stage_alu_shifter_N159);
   dp_ex_stage_alu_shifter_srl_41_U135 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n26, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n99, ZN => 
                           dp_ex_stage_alu_shifter_N160);
   dp_ex_stage_alu_shifter_srl_41_U134 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n138, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n134, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n93);
   dp_ex_stage_alu_shifter_srl_41_U133 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n26, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n93, ZN => 
                           dp_ex_stage_alu_shifter_N161);
   dp_ex_stage_alu_shifter_srl_41_U132 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n136, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n133, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n85);
   dp_ex_stage_alu_shifter_srl_41_U131 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n26, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n85, ZN => 
                           dp_ex_stage_alu_shifter_N162);
   dp_ex_stage_alu_shifter_srl_41_U130 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n26, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n135, ZN => 
                           dp_ex_stage_alu_shifter_N163);
   dp_ex_stage_alu_shifter_srl_41_U129 : NOR3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n73, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n28, A3 => 
                           dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_shifter_N164);
   dp_ex_stage_alu_shifter_srl_41_U128 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n134, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, ZN => 
                           dp_ex_stage_alu_shifter_N165);
   dp_ex_stage_alu_shifter_srl_41_U127 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n133, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, ZN => 
                           dp_ex_stage_alu_shifter_N166);
   dp_ex_stage_alu_shifter_srl_41_U126 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n32, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n56, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n132);
   dp_ex_stage_alu_shifter_srl_41_U125 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n69, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_n44, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n131);
   dp_ex_stage_alu_shifter_srl_41_U124 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n55, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n22, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n54, A => 
                           dp_ex_stage_alu_shifter_srl_41_n131, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n129);
   dp_ex_stage_alu_shifter_srl_41_U123 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n106, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n129, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n59, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n128);
   dp_ex_stage_alu_shifter_srl_41_U122 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n103, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n114, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n127, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n128, ZN => 
                           dp_ex_stage_alu_shifter_N139);
   dp_ex_stage_alu_shifter_srl_41_U121 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n126, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, ZN => 
                           dp_ex_stage_alu_shifter_N167);
   dp_ex_stage_alu_shifter_srl_41_U120 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n125, ZN => 
                           dp_ex_stage_alu_shifter_N168);
   dp_ex_stage_alu_shifter_srl_41_U119 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n33, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n32, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n124);
   dp_ex_stage_alu_shifter_srl_41_U118 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n52, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n20, B1 => 
                           dp_ex_stage_alu_n69, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n18, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n121);
   dp_ex_stage_alu_shifter_srl_41_U117 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n1, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n56, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n55, A => 
                           dp_ex_stage_alu_shifter_srl_41_n121, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n117);
   dp_ex_stage_alu_shifter_srl_41_U116 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n101, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n117, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n60, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n116);
   dp_ex_stage_alu_shifter_srl_41_U115 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n98, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n114, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n115, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n116, ZN => 
                           dp_ex_stage_alu_shifter_N140);
   dp_ex_stage_alu_shifter_srl_41_U114 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n80, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n57, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n95, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n96, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n113);
   dp_ex_stage_alu_shifter_srl_41_U113 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n111, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n112, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n113, ZN => 
                           dp_ex_stage_alu_shifter_N141);
   dp_ex_stage_alu_shifter_srl_41_U112 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n80, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n58, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n87, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n89, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n110);
   dp_ex_stage_alu_shifter_srl_41_U111 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n108, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n109, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n110, ZN => 
                           dp_ex_stage_alu_shifter_N142);
   dp_ex_stage_alu_shifter_srl_41_U110 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n80, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n59, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n106, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n107, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n105);
   dp_ex_stage_alu_shifter_srl_41_U109 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n103, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n104, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n105, ZN => 
                           dp_ex_stage_alu_shifter_N143);
   dp_ex_stage_alu_shifter_srl_41_U108 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n80, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n60, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n101, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n102, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n100);
   dp_ex_stage_alu_shifter_srl_41_U107 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n98, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n99, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n100, ZN => 
                           dp_ex_stage_alu_shifter_N144);
   dp_ex_stage_alu_shifter_srl_41_U106 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n80, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n95, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n96, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n97, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n94);
   dp_ex_stage_alu_shifter_srl_41_U105 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n92, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n93, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n94, ZN => 
                           dp_ex_stage_alu_shifter_N145);
   dp_ex_stage_alu_shifter_srl_41_U104 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n80, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n87, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n89, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n91, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n86);
   dp_ex_stage_alu_shifter_srl_41_U103 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n83, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n84, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n85, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, A => 
                           dp_ex_stage_alu_shifter_srl_41_n86, ZN => 
                           dp_ex_stage_alu_shifter_N146);
   dp_ex_stage_alu_shifter_srl_41_U102 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_31_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n53);
   dp_ex_stage_alu_shifter_srl_41_U101 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n1, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n52);
   dp_ex_stage_alu_shifter_srl_41_U100 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_27_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n51);
   dp_ex_stage_alu_shifter_srl_41_U99 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_26_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n50);
   dp_ex_stage_alu_shifter_srl_41_U98 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_25_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n49);
   dp_ex_stage_alu_shifter_srl_41_U97 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_24_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n48);
   dp_ex_stage_alu_shifter_srl_41_U96 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_23_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n47);
   dp_ex_stage_alu_shifter_srl_41_U95 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_21_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n46);
   dp_ex_stage_alu_shifter_srl_41_U94 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_18_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n45);
   dp_ex_stage_alu_shifter_srl_41_U93 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_17_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n44);
   dp_ex_stage_alu_shifter_srl_41_U92 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n38, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n43);
   dp_ex_stage_alu_shifter_srl_41_U91 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n29, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n42);
   dp_ex_stage_alu_shifter_srl_41_U90 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n42, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n41);
   dp_ex_stage_alu_shifter_srl_41_U89 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_14_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n40);
   dp_ex_stage_alu_shifter_srl_41_U88 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n40, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n39);
   dp_ex_stage_alu_shifter_srl_41_U87 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_12_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n38);
   dp_ex_stage_alu_shifter_srl_41_U86 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n38, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n37);
   dp_ex_stage_alu_shifter_srl_41_U85 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n33, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n36);
   dp_ex_stage_alu_shifter_srl_41_U84 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n74, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n35);
   dp_ex_stage_alu_shifter_srl_41_U83 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n72, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n34);
   dp_ex_stage_alu_shifter_srl_41_U82 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n71, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n33);
   dp_ex_stage_alu_shifter_srl_41_U81 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n34, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n32);
   dp_ex_stage_alu_shifter_srl_41_U80 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n69, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n31);
   dp_ex_stage_alu_shifter_srl_41_U79 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n44, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n30);
   dp_ex_stage_alu_shifter_srl_41_U78 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n25);
   dp_ex_stage_alu_shifter_srl_41_U77 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n49, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n24);
   dp_ex_stage_alu_shifter_srl_41_U76 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n45, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n23);
   dp_ex_stage_alu_shifter_srl_41_U75 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n23, A2 => 
                           dp_ex_stage_alu_n46, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n122);
   dp_ex_stage_alu_shifter_srl_41_U74 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n163, ZN => 
                           dp_ex_stage_alu_shifter_N149);
   dp_ex_stage_alu_shifter_srl_41_U73 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n52, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n54);
   dp_ex_stage_alu_shifter_srl_41_U72 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n122, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n20);
   dp_ex_stage_alu_shifter_srl_41_U71 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n122, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n19);
   dp_ex_stage_alu_shifter_srl_41_U70 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_n45, A2 => dp_ex_stage_alu_n46, ZN 
                           => dp_ex_stage_alu_shifter_srl_41_n123);
   dp_ex_stage_alu_shifter_srl_41_U69 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n123, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n18);
   dp_ex_stage_alu_shifter_srl_41_U68 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n78, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n56);
   dp_ex_stage_alu_shifter_srl_41_U67 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n70, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n55);
   dp_ex_stage_alu_shifter_srl_41_U66 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_29_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n74);
   dp_ex_stage_alu_shifter_srl_41_U65 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_19_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n68);
   dp_ex_stage_alu_shifter_srl_41_U64 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_30_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n75);
   dp_ex_stage_alu_shifter_srl_41_U63 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_20_port, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n69);
   dp_ex_stage_alu_shifter_srl_41_U62 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n92, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n57);
   dp_ex_stage_alu_shifter_srl_41_U61 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n150, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n73);
   dp_ex_stage_alu_shifter_srl_41_U60 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n107, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n66);
   dp_ex_stage_alu_shifter_srl_41_U59 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n83, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n58);
   dp_ex_stage_alu_shifter_srl_41_U58 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n119, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n79);
   dp_ex_stage_alu_shifter_srl_41_U57 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n184, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n70);
   dp_ex_stage_alu_shifter_srl_41_U56 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n151, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n72);
   dp_ex_stage_alu_shifter_srl_41_U55 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n153, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n71);
   dp_ex_stage_alu_shifter_srl_41_U54 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n89, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n65);
   dp_ex_stage_alu_shifter_srl_41_U53 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n102, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n67);
   dp_ex_stage_alu_shifter_srl_41_U52 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n87, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n62);
   dp_ex_stage_alu_shifter_srl_41_U51 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n106, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n63);
   dp_ex_stage_alu_shifter_srl_41_U50 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n101, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n64);
   dp_ex_stage_alu_shifter_srl_41_U49 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n120, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n22);
   dp_ex_stage_alu_shifter_srl_41_U48 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n118, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n60);
   dp_ex_stage_alu_shifter_srl_41_U47 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n130, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n59);
   dp_ex_stage_alu_shifter_srl_41_U46 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n120, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n77);
   dp_ex_stage_alu_shifter_srl_41_U45 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n114, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n80);
   dp_ex_stage_alu_shifter_srl_41_U44 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n164, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n82);
   dp_ex_stage_alu_shifter_srl_41_U43 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n28, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n29);
   dp_ex_stage_alu_shifter_srl_41_U42 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n84, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n81);
   dp_ex_stage_alu_shifter_srl_41_U41 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n27);
   dp_ex_stage_alu_shifter_srl_41_U40 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n26);
   dp_ex_stage_alu_shifter_srl_41_U39 : INV_X2 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n123, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n76);
   dp_ex_stage_alu_shifter_srl_41_U38 : INV_X2 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n19, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n78);
   dp_ex_stage_alu_shifter_srl_41_U37 : NAND3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n16, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n17, A3 => 
                           dp_ex_stage_alu_shifter_srl_41_n188, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n97);
   dp_ex_stage_alu_shifter_srl_41_U36 : OR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n69, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n76, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n17);
   dp_ex_stage_alu_shifter_srl_41_U35 : OR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n78, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n46, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n16);
   dp_ex_stage_alu_shifter_srl_41_U34 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n97, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n15);
   dp_ex_stage_alu_shifter_srl_41_U33 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n156, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n134, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n14);
   dp_ex_stage_alu_shifter_srl_41_U32 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n138, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n13);
   dp_ex_stage_alu_shifter_srl_41_U31 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, A2 => 
                           dp_ex_stage_alu_n74, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n12);
   dp_ex_stage_alu_shifter_srl_41_U30 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, A2 => 
                           dp_ex_stage_alu_n33, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n11);
   dp_ex_stage_alu_shifter_srl_41_U29 : AND3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n8, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n9, A3 => 
                           dp_ex_stage_alu_shifter_srl_41_n10, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n178);
   dp_ex_stage_alu_shifter_srl_41_U28 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n88, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n57, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n10);
   dp_ex_stage_alu_shifter_srl_41_U27 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n81, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n179, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n9);
   dp_ex_stage_alu_shifter_srl_41_U26 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n90, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n95, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n8);
   dp_ex_stage_alu_shifter_srl_41_U25 : CLKBUF_X3 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n120, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n21);
   dp_ex_stage_alu_shifter_srl_41_U24 : NAND3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n6, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n7, A3 => 
                           dp_ex_stage_alu_shifter_srl_41_n186, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n134);
   dp_ex_stage_alu_shifter_srl_41_U23 : OR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n75, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n7);
   dp_ex_stage_alu_shifter_srl_41_U22 : OR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n53, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n6);
   dp_ex_stage_alu_shifter_srl_41_U21 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n139, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n125, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n140, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n141, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n99);
   dp_ex_stage_alu_shifter_srl_41_U20 : NAND3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n4, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n5, A3 => 
                           dp_ex_stage_alu_shifter_srl_41_n167, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n139);
   dp_ex_stage_alu_shifter_srl_41_U19 : OR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n21, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n74, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n5);
   dp_ex_stage_alu_shifter_srl_41_U18 : OR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n119, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n75, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n4);
   dp_ex_stage_alu_shifter_srl_41_U17 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n45, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n3);
   dp_ex_stage_alu_shifter_srl_41_U16 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n181, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n24, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n88);
   dp_ex_stage_alu_shifter_srl_41_U15 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n138, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n137, B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n134, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n140, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n97, C2 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n112);
   dp_ex_stage_alu_shifter_srl_41_U14 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n49, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n181, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n90);
   dp_ex_stage_alu_shifter_srl_41_U13 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B2 => 
                           dp_ex_stage_alu_shifter_srl_41_n39, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, C2 => 
                           dp_ex_stage_alu_n231, A => 
                           dp_ex_stage_alu_shifter_srl_41_n170, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n118);
   dp_ex_stage_alu_shifter_srl_41_U12 : NAND2_X2 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n82, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n29, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n84);
   dp_ex_stage_alu_shifter_srl_41_U11 : OR3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n13, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n14, A3 => 
                           dp_ex_stage_alu_shifter_srl_41_n15, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n2);
   dp_ex_stage_alu_shifter_srl_41_U10 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_srl_41_n28);
   dp_ex_stage_alu_shifter_srl_41_U9 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n46, A2 => dp_ex_stage_alu_n45, ZN 
                           => dp_ex_stage_alu_shifter_srl_41_n119);
   dp_ex_stage_alu_shifter_srl_41_U8 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_srl_41_n79, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n1);
   dp_ex_stage_alu_shifter_srl_41_U7 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B2 => 
                           dp_ex_stage_alu_n71, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, C2 => 
                           dp_ex_stage_alu_n34, A => 
                           dp_ex_stage_alu_shifter_srl_41_n149, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n108);
   dp_ex_stage_alu_shifter_srl_41_U6 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B2 => 
                           dp_ex_stage_alu_n74, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, C2 => 
                           dp_ex_stage_alu_n72, A => 
                           dp_ex_stage_alu_shifter_srl_41_n124, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n98);
   dp_ex_stage_alu_shifter_srl_41_U5 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B2 => 
                           dp_ex_stage_alu_n34, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, C2 => 
                           dp_ex_stage_alu_n78, A => 
                           dp_ex_stage_alu_shifter_srl_41_n189, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n111);
   dp_ex_stage_alu_shifter_srl_41_U4 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_srl_41_n79, B2 => 
                           dp_ex_stage_alu_n72, C1 => 
                           dp_ex_stage_alu_shifter_srl_41_n77, C2 => 
                           dp_ex_stage_alu_n71, A => 
                           dp_ex_stage_alu_shifter_srl_41_n132, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n103);
   dp_ex_stage_alu_shifter_srl_41_U3 : NOR3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_srl_41_n11, A2 => 
                           dp_ex_stage_alu_shifter_srl_41_n12, A3 => 
                           dp_ex_stage_alu_shifter_srl_41_n180, ZN => 
                           dp_ex_stage_alu_shifter_srl_41_n92);
   dp_ex_stage_alu_shifter_sra_39_U225 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n47, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n46, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n13, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n193);
   dp_ex_stage_alu_shifter_sra_39_U224 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n17, A2 => 
                           dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n131);
   dp_ex_stage_alu_shifter_sra_39_U223 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n107);
   dp_ex_stage_alu_shifter_sra_39_U222 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n240, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n37, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n192);
   dp_ex_stage_alu_shifter_sra_39_U221 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n36, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n63, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n12, A => 
                           dp_ex_stage_alu_shifter_sra_39_n192, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n91);
   dp_ex_stage_alu_shifter_sra_39_U220 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n32, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_alu_n38, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n191);
   dp_ex_stage_alu_shifter_sra_39_U219 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n34, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n62, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, A => 
                           dp_ex_stage_alu_shifter_sra_39_n191, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n90);
   dp_ex_stage_alu_shifter_sra_39_U218 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n49, A2 => dp_ex_stage_alu_n31, ZN 
                           => dp_ex_stage_alu_shifter_sra_39_n155);
   dp_ex_stage_alu_shifter_sra_39_U217 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_29_port, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_alu_n1, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n190);
   dp_ex_stage_alu_shifter_sra_39_U216 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n70, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n45, A => 
                           dp_ex_stage_alu_shifter_sra_39_n190, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n134);
   dp_ex_stage_alu_shifter_sra_39_U215 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n31, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n17, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n141);
   dp_ex_stage_alu_shifter_sra_39_U214 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_25_port, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n14, B1 => 
                           dp_ex_stage_muxA_out_24_port, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n189);
   dp_ex_stage_alu_shifter_sra_39_U213 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n155, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n134, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n141, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n135, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n188);
   dp_ex_stage_alu_shifter_sra_39_U212 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n31, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n22, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n185);
   dp_ex_stage_alu_shifter_sra_39_U211 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n49, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n185, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n85);
   dp_ex_stage_alu_shifter_sra_39_U210 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n231, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n30, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n15, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n187);
   dp_ex_stage_alu_shifter_sra_39_U209 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n76, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n14, B1 => 
                           dp_ex_stage_alu_shifter_N202, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n186);
   dp_ex_stage_alu_shifter_sra_39_U208 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n27, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n26, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n13, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n184);
   dp_ex_stage_alu_shifter_sra_39_U207 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n53, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n77, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n183, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n49, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n182);
   dp_ex_stage_alu_shifter_sra_39_U206 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n104, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n107, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n158, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n182, ZN => 
                           dp_ex_stage_alu_shifter_N105_port);
   dp_ex_stage_alu_shifter_sra_39_U205 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n29, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n28, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n13, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n181);
   dp_ex_stage_alu_shifter_sra_39_U204 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_30_port, B => 
                           dp_ex_stage_alu_shifter_N136, S => 
                           dp_ex_stage_alu_shifter_sra_39_n12, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n142);
   dp_ex_stage_alu_shifter_sra_39_U203 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_27_port, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_muxA_out_26_port, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n180);
   dp_ex_stage_alu_shifter_sra_39_U202 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_N136, A2 => 
                           dp_ex_stage_alu_n31, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n154);
   dp_ex_stage_alu_shifter_sra_39_U201 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n142, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n138, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n71, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n129);
   dp_ex_stage_alu_shifter_sra_39_U200 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n29, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n14, B1 => 
                           dp_ex_stage_muxA_out_14_port, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n15, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n179);
   dp_ex_stage_alu_shifter_sra_39_U199 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_20_port, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n35, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n178);
   dp_ex_stage_alu_shifter_sra_39_U198 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n62, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n34, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n12, A => 
                           dp_ex_stage_alu_shifter_sra_39_n178, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n100);
   dp_ex_stage_alu_shifter_sra_39_U197 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n37, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_alu_n240, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n15, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n177);
   dp_ex_stage_alu_shifter_sra_39_U196 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n39, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n40, A => 
                           dp_ex_stage_alu_shifter_sra_39_n177, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n139);
   dp_ex_stage_alu_shifter_sra_39_U195 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n57, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n100, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n139, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n176);
   dp_ex_stage_alu_shifter_sra_39_U194 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n123, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n129, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n176, ZN => 
                           dp_ex_stage_alu_shifter_N115_port);
   dp_ex_stage_alu_shifter_sra_39_U193 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n31, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n29, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n13, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n175);
   dp_ex_stage_alu_shifter_sra_39_U192 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n1, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n14, B1 => 
                           dp_ex_stage_muxA_out_27_port, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n174);
   dp_ex_stage_alu_shifter_sra_39_U191 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n68, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n70, A => 
                           dp_ex_stage_alu_shifter_sra_39_n174, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n136);
   dp_ex_stage_alu_shifter_sra_39_U190 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n17, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n45, A => 
                           dp_ex_stage_alu_shifter_sra_39_n154, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n162);
   dp_ex_stage_alu_shifter_sra_39_U189 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n136, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n162, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n128);
   dp_ex_stage_alu_shifter_sra_39_U188 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n38, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_alu_n29, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n173);
   dp_ex_stage_alu_shifter_sra_39_U187 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n35, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B1 => 
                           dp_ex_stage_alu_n240, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n172);
   dp_ex_stage_alu_shifter_sra_39_U186 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n63, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n62, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n13, A => 
                           dp_ex_stage_alu_shifter_sra_39_n172, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n96);
   dp_ex_stage_alu_shifter_sra_39_U185 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_24_port, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n14, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n37, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n171);
   dp_ex_stage_alu_shifter_sra_39_U184 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n95, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n96, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n137, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n170);
   dp_ex_stage_alu_shifter_sra_39_U183 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n111, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n128, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n170, ZN => 
                           dp_ex_stage_alu_shifter_N116_port);
   dp_ex_stage_alu_shifter_sra_39_U182 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n7, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n162, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n127);
   dp_ex_stage_alu_shifter_sra_39_U181 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n90, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n91, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n135, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n169);
   dp_ex_stage_alu_shifter_sra_39_U180 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n168, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n127, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n169, ZN => 
                           dp_ex_stage_alu_shifter_N117_port);
   dp_ex_stage_alu_shifter_sra_39_U179 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_14_port, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n14, B1 => 
                           dp_ex_stage_alu_n231, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n15, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n167);
   dp_ex_stage_alu_shifter_sra_39_U178 : OAI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n13, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n68, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n70, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n3, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n45, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n130);
   dp_ex_stage_alu_shifter_sra_39_U177 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n130, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n162, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n126);
   dp_ex_stage_alu_shifter_sra_39_U176 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_18_port, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n14, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n32, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n166);
   dp_ex_stage_alu_shifter_sra_39_U175 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n240, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n14, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n35, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n165);
   dp_ex_stage_alu_shifter_sra_39_U174 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_26_port, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_muxA_out_25_port, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n15, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n164);
   dp_ex_stage_alu_shifter_sra_39_U173 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n42, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n43, A => 
                           dp_ex_stage_alu_shifter_sra_39_n164, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n132);
   dp_ex_stage_alu_shifter_sra_39_U172 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n84, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n86, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n132, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n163);
   dp_ex_stage_alu_shifter_sra_39_U171 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n151, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n126, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n163, ZN => 
                           dp_ex_stage_alu_shifter_N118_port);
   dp_ex_stage_alu_shifter_sra_39_U170 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n142, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n162, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n118);
   dp_ex_stage_alu_shifter_sra_39_U169 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n100, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n139, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n138, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n161);
   dp_ex_stage_alu_shifter_sra_39_U168 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n160, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n118, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n161, ZN => 
                           dp_ex_stage_alu_shifter_N119);
   dp_ex_stage_alu_shifter_sra_39_U167 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n136, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n137, A => 
                           dp_ex_stage_alu_shifter_sra_39_n72, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n159);
   dp_ex_stage_alu_shifter_sra_39_U166 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n61, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n107, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n59, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, A => 
                           dp_ex_stage_alu_shifter_sra_39_n159, ZN => 
                           dp_ex_stage_alu_shifter_N120);
   dp_ex_stage_alu_shifter_sra_39_U165 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n20, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n158, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N121);
   dp_ex_stage_alu_shifter_sra_39_U164 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n155, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n130, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n132, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n141, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n157);
   dp_ex_stage_alu_shifter_sra_39_U163 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n20, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n146, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N122);
   dp_ex_stage_alu_shifter_sra_39_U162 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n139, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n100, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n156);
   dp_ex_stage_alu_shifter_sra_39_U161 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n142, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n155, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n138, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n141, A => 
                           dp_ex_stage_alu_shifter_sra_39_n60, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n120);
   dp_ex_stage_alu_shifter_sra_39_U160 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n20, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n120, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N123);
   dp_ex_stage_alu_shifter_sra_39_U159 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n154, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n17, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n143);
   dp_ex_stage_alu_shifter_sra_39_U158 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n141, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n136, A => 
                           dp_ex_stage_alu_shifter_sra_39_n143, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n153);
   dp_ex_stage_alu_shifter_sra_39_U157 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n19, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n108, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N124);
   dp_ex_stage_alu_shifter_sra_39_U156 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n48, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n47, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n12, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n152);
   dp_ex_stage_alu_shifter_sra_39_U155 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n44, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_alu_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n150);
   dp_ex_stage_alu_shifter_sra_39_U154 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n28, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n27, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n13, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n149);
   dp_ex_stage_alu_shifter_sra_39_U153 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n55, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n77, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n148, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n50, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n147);
   dp_ex_stage_alu_shifter_sra_39_U152 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n101, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n107, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n146, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n147, ZN => 
                           dp_ex_stage_alu_shifter_N106_port);
   dp_ex_stage_alu_shifter_sra_39_U151 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n141, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n134, A => 
                           dp_ex_stage_alu_shifter_sra_39_n143, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n145);
   dp_ex_stage_alu_shifter_sra_39_U150 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n19, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n105, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N125);
   dp_ex_stage_alu_shifter_sra_39_U149 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n141, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n130, A => 
                           dp_ex_stage_alu_shifter_sra_39_n143, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n144);
   dp_ex_stage_alu_shifter_sra_39_U148 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n19, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n102, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N126);
   dp_ex_stage_alu_shifter_sra_39_U147 : AOI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n141, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n142, A => 
                           dp_ex_stage_alu_shifter_sra_39_n143, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n140);
   dp_ex_stage_alu_shifter_sra_39_U146 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n19, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n98, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N127);
   dp_ex_stage_alu_shifter_sra_39_U145 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n19, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n93, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N128);
   dp_ex_stage_alu_shifter_sra_39_U144 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n19, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n88, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N129);
   dp_ex_stage_alu_shifter_sra_39_U143 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n19, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n81, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N130);
   dp_ex_stage_alu_shifter_sra_39_U142 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n18, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n129, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N131);
   dp_ex_stage_alu_shifter_sra_39_U141 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n18, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n128, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N132);
   dp_ex_stage_alu_shifter_sra_39_U140 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n18, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n127, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N133);
   dp_ex_stage_alu_shifter_sra_39_U139 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n18, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n126, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N134);
   dp_ex_stage_alu_shifter_sra_39_U138 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n25, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n48, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n12, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n125);
   dp_ex_stage_alu_shifter_sra_39_U137 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n69, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_alu_n44, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n124);
   dp_ex_stage_alu_shifter_sra_39_U136 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n57, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n77, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n122, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n51, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n121);
   dp_ex_stage_alu_shifter_sra_39_U135 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n97, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n107, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n120, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n121, ZN => 
                           dp_ex_stage_alu_shifter_N107_port);
   dp_ex_stage_alu_shifter_sra_39_U134 : OAI21_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n18, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n118, A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_N135);
   dp_ex_stage_alu_shifter_sra_39_U133 : OAI22_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n26, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n10, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n25, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n13, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n115);
   dp_ex_stage_alu_shifter_sra_39_U132 : AOI22_X1 port map( A1 => 
                           dp_ex_stage_alu_n52, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n73, B1 => 
                           dp_ex_stage_alu_n69, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n75, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n112);
   dp_ex_stage_alu_shifter_sra_39_U131 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n95, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n77, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n110, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n52, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n109);
   dp_ex_stage_alu_shifter_sra_39_U130 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n92, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n107, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n108, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n22, A => 
                           dp_ex_stage_alu_shifter_sra_39_n109, ZN => 
                           dp_ex_stage_alu_shifter_N108_port);
   dp_ex_stage_alu_shifter_sra_39_U129 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n49, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n53, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n90, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n106);
   dp_ex_stage_alu_shifter_sra_39_U128 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n104, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n105, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n22, A => 
                           dp_ex_stage_alu_shifter_sra_39_n106, ZN => 
                           dp_ex_stage_alu_shifter_N109_port);
   dp_ex_stage_alu_shifter_sra_39_U127 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n50, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n55, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n84, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n103);
   dp_ex_stage_alu_shifter_sra_39_U126 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n101, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n102, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n22, A => 
                           dp_ex_stage_alu_shifter_sra_39_n103, ZN => 
                           dp_ex_stage_alu_shifter_N110_port);
   dp_ex_stage_alu_shifter_sra_39_U125 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n51, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n57, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n100, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n99);
   dp_ex_stage_alu_shifter_sra_39_U124 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n97, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n98, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n22, A => 
                           dp_ex_stage_alu_shifter_sra_39_n99, ZN => 
                           dp_ex_stage_alu_shifter_N111_port);
   dp_ex_stage_alu_shifter_sra_39_U123 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n52, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n95, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n96, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n94);
   dp_ex_stage_alu_shifter_sra_39_U122 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n92, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n93, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n22, A => 
                           dp_ex_stage_alu_shifter_sra_39_n94, ZN => 
                           dp_ex_stage_alu_shifter_N112_port);
   dp_ex_stage_alu_shifter_sra_39_U121 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n53, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n90, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n91, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n89);
   dp_ex_stage_alu_shifter_sra_39_U120 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n87, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n88, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n89, ZN => 
                           dp_ex_stage_alu_shifter_N113_port);
   dp_ex_stage_alu_shifter_sra_39_U119 : AOI222_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n78, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n55, B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n83, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n84, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n85, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n86, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n82);
   dp_ex_stage_alu_shifter_sra_39_U118 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n79, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n80, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n81, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, A => 
                           dp_ex_stage_alu_shifter_sra_39_n82, ZN => 
                           dp_ex_stage_alu_shifter_N114_port);
   dp_ex_stage_alu_shifter_sra_39_U117 : INV_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n113, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n76);
   dp_ex_stage_alu_shifter_sra_39_U116 : INV_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n114, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n74);
   dp_ex_stage_alu_shifter_sra_39_U115 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n45, ZN => 
                           dp_ex_stage_alu_shifter_N136);
   dp_ex_stage_alu_shifter_sra_39_U114 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n1, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n43);
   dp_ex_stage_alu_shifter_sra_39_U113 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_27_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n42);
   dp_ex_stage_alu_shifter_sra_39_U112 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_26_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n41);
   dp_ex_stage_alu_shifter_sra_39_U111 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_25_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n40);
   dp_ex_stage_alu_shifter_sra_39_U110 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_24_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n39);
   dp_ex_stage_alu_shifter_sra_39_U109 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_23_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n38);
   dp_ex_stage_alu_shifter_sra_39_U108 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n38, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n37);
   dp_ex_stage_alu_shifter_sra_39_U107 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_21_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n36);
   dp_ex_stage_alu_shifter_sra_39_U106 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n36, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n35);
   dp_ex_stage_alu_shifter_sra_39_U105 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_18_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n34);
   dp_ex_stage_alu_shifter_sra_39_U104 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_17_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n33);
   dp_ex_stage_alu_shifter_sra_39_U103 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n33, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n32);
   dp_ex_stage_alu_shifter_sra_39_U102 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_12_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n31);
   dp_ex_stage_alu_shifter_sra_39_U101 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n31, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n30);
   dp_ex_stage_alu_shifter_sra_39_U100 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n33, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n29);
   dp_ex_stage_alu_shifter_sra_39_U99 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n74, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n28);
   dp_ex_stage_alu_shifter_sra_39_U98 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n72, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n27);
   dp_ex_stage_alu_shifter_sra_39_U97 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n71, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n26);
   dp_ex_stage_alu_shifter_sra_39_U96 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n34, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n25);
   dp_ex_stage_alu_shifter_sra_39_U95 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n69, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n24);
   dp_ex_stage_alu_shifter_sra_39_U94 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n44, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n23);
   dp_ex_stage_alu_shifter_sra_39_U93 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n18, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n22);
   dp_ex_stage_alu_shifter_sra_39_U92 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n49, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n17);
   dp_ex_stage_alu_shifter_sra_39_U91 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n45, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n16);
   dp_ex_stage_alu_shifter_sra_39_U90 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n160, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n57);
   dp_ex_stage_alu_shifter_sra_39_U89 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n168, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n53);
   dp_ex_stage_alu_shifter_sra_39_U88 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n167, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n56);
   dp_ex_stage_alu_shifter_sra_39_U87 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n151, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n55);
   dp_ex_stage_alu_shifter_sra_39_U86 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n179, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n58);
   dp_ex_stage_alu_shifter_sra_39_U85 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n187, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n54);
   dp_ex_stage_alu_shifter_sra_39_U84 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n156, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n60);
   dp_ex_stage_alu_shifter_sra_39_U83 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n153, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n65);
   dp_ex_stage_alu_shifter_sra_39_U82 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n157, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n64);
   dp_ex_stage_alu_shifter_sra_39_U81 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n11, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n15);
   dp_ex_stage_alu_shifter_sra_39_U80 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n52, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n46);
   dp_ex_stage_alu_shifter_sra_39_U79 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n9, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n73);
   dp_ex_stage_alu_shifter_sra_39_U78 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n9, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n14);
   dp_ex_stage_alu_shifter_sra_39_U77 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n16, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n4, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n117);
   dp_ex_stage_alu_shifter_sra_39_U76 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n117, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n12);
   dp_ex_stage_alu_shifter_sra_39_U75 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_n45, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n3, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n116);
   dp_ex_stage_alu_shifter_sra_39_U74 : CLKBUF_X3 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n116, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n10);
   dp_ex_stage_alu_shifter_sra_39_U73 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n78, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n48);
   dp_ex_stage_alu_shifter_sra_39_U72 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n116, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n9);
   dp_ex_stage_alu_shifter_sra_39_U71 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_muxA_out_14_port, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_n29, A => 
                           dp_ex_stage_alu_shifter_sra_39_n54, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n168);
   dp_ex_stage_alu_shifter_sra_39_U70 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n70, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n47);
   dp_ex_stage_alu_shifter_sra_39_U69 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_30_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n70);
   dp_ex_stage_alu_shifter_sra_39_U68 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_20_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n63);
   dp_ex_stage_alu_shifter_sra_39_U67 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_29_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n68);
   dp_ex_stage_alu_shifter_sra_39_U66 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_19_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n62);
   dp_ex_stage_alu_shifter_sra_39_U65 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n38, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n32, A => 
                           dp_ex_stage_alu_shifter_sra_39_n58, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n160);
   dp_ex_stage_alu_shifter_sra_39_U64 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n144, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n67);
   dp_ex_stage_alu_shifter_sra_39_U63 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n140, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n69);
   dp_ex_stage_alu_shifter_sra_39_U62 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n145, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n66);
   dp_ex_stage_alu_shifter_sra_39_U61 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n154, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n71);
   dp_ex_stage_alu_shifter_sra_39_U60 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n95, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n59);
   dp_ex_stage_alu_shifter_sra_39_U59 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n79, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n50);
   dp_ex_stage_alu_shifter_sra_39_U58 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n111, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n52);
   dp_ex_stage_alu_shifter_sra_39_U57 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n87, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n49);
   dp_ex_stage_alu_shifter_sra_39_U56 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_31_port, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n45);
   dp_ex_stage_alu_shifter_sra_39_U55 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n119, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n72);
   dp_ex_stage_alu_shifter_sra_39_U54 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n96, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n61);
   dp_ex_stage_alu_shifter_sra_39_U53 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n123, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n51);
   dp_ex_stage_alu_shifter_sra_39_U52 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n117, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n13);
   dp_ex_stage_alu_shifter_sra_39_U51 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n80, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n77);
   dp_ex_stage_alu_shifter_sra_39_U50 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n107, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n78);
   dp_ex_stage_alu_shifter_sra_39_U49 : INV_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n18, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n21);
   dp_ex_stage_alu_shifter_sra_39_U48 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n20, A2 => 
                           dp_ex_stage_alu_shifter_N136, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n119);
   dp_ex_stage_alu_shifter_sra_39_U47 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n20);
   dp_ex_stage_alu_shifter_sra_39_U46 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n19);
   dp_ex_stage_alu_shifter_sra_39_U45 : BUF_X2 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n18);
   dp_ex_stage_alu_shifter_sra_39_U44 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n135, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n8);
   dp_ex_stage_alu_shifter_sra_39_U43 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n134, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n7);
   dp_ex_stage_alu_shifter_sra_39_U42 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n90, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n6);
   dp_ex_stage_alu_shifter_sra_39_U41 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n91, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n5);
   dp_ex_stage_alu_shifter_sra_39_U40 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n86, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n84, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n64, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n146);
   dp_ex_stage_alu_shifter_sra_39_U39 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n137, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n96, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n65, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n108);
   dp_ex_stage_alu_shifter_sra_39_U38 : OAI221_X4 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n47, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n48, A => 
                           dp_ex_stage_alu_shifter_sra_39_n112, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n110);
   dp_ex_stage_alu_shifter_sra_39_U37 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n46, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n4);
   dp_ex_stage_alu_shifter_sra_39_U36 : INV_X1 port map( A => 
                           dp_ex_stage_alu_n46, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n3);
   dp_ex_stage_alu_shifter_sra_39_U35 : NOR2_X2 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n16, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n3, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n114);
   dp_ex_stage_alu_shifter_sra_39_U34 : AND3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n5, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n6, A3 => 
                           dp_ex_stage_alu_shifter_sra_39_n188, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n158);
   dp_ex_stage_alu_shifter_sra_39_U33 : INV_X2 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n11, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n75);
   dp_ex_stage_alu_shifter_sra_39_U32 : NAND3_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n1, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n2, A3 => 
                           dp_ex_stage_alu_shifter_sra_39_n189, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n135);
   dp_ex_stage_alu_shifter_sra_39_U31 : OR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n42, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n2);
   dp_ex_stage_alu_shifter_sra_39_U30 : OR2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n41, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n1);
   dp_ex_stage_alu_shifter_sra_39_U29 : NOR2_X2 port map( A1 => 
                           dp_ex_stage_alu_n49, A2 => dp_ex_stage_alu_n31, ZN 
                           => dp_ex_stage_alu_shifter_sra_39_n133);
   dp_ex_stage_alu_shifter_sra_39_U28 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n130, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n132, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n71, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n81);
   dp_ex_stage_alu_shifter_sra_39_U27 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n21, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n80);
   dp_ex_stage_alu_shifter_sra_39_U26 : AND2_X1 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n185, A2 => 
                           dp_ex_stage_alu_shifter_sra_39_n17, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n83);
   dp_ex_stage_alu_shifter_sra_39_U25 : NOR2_X2 port map( A1 => 
                           dp_ex_stage_alu_shifter_sra_39_n4, A2 => 
                           dp_ex_stage_alu_n45, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n113);
   dp_ex_stage_alu_shifter_sra_39_U24 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n23, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n24, A => 
                           dp_ex_stage_alu_shifter_sra_39_n186, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n183);
   dp_ex_stage_alu_shifter_sra_39_U23 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n34, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_n71, A => 
                           dp_ex_stage_alu_shifter_sra_39_n152, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n101);
   dp_ex_stage_alu_shifter_sra_39_U22 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n24, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n46, A => 
                           dp_ex_stage_alu_shifter_sra_39_n150, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n148);
   dp_ex_stage_alu_shifter_sra_39_U21 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n46, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n47, A => 
                           dp_ex_stage_alu_shifter_sra_39_n124, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n122);
   dp_ex_stage_alu_shifter_sra_39_U20 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n72, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_n74, A => 
                           dp_ex_stage_alu_shifter_sra_39_n115, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n92);
   dp_ex_stage_alu_shifter_sra_39_U19 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n8, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n91, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n66, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n105);
   dp_ex_stage_alu_shifter_sra_39_U18 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n132, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n86, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n67, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n102);
   dp_ex_stage_alu_shifter_sra_39_U17 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n138, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n139, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n69, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n98);
   dp_ex_stage_alu_shifter_sra_39_U16 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n136, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n137, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n71, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n93);
   dp_ex_stage_alu_shifter_sra_39_U15 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n7, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n131, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n8, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n133, A => 
                           dp_ex_stage_alu_shifter_sra_39_n71, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n88);
   dp_ex_stage_alu_shifter_sra_39_U14 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n231, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_muxA_out_14_port, A => 
                           dp_ex_stage_alu_shifter_sra_39_n175, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n111);
   dp_ex_stage_alu_shifter_sra_39_U13 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n62, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n63, A => 
                           dp_ex_stage_alu_shifter_sra_39_n166, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n84);
   dp_ex_stage_alu_shifter_sra_39_U12 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n33, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n34, A => 
                           dp_ex_stage_alu_shifter_sra_39_n173, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n95);
   dp_ex_stage_alu_shifter_sra_39_U11 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n40, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n41, A => 
                           dp_ex_stage_alu_shifter_sra_39_n171, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n137);
   dp_ex_stage_alu_shifter_sra_39_U10 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n78, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_n34, A => 
                           dp_ex_stage_alu_shifter_sra_39_n193, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n104);
   dp_ex_stage_alu_shifter_sra_39_U9 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n71, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_n72, A => 
                           dp_ex_stage_alu_shifter_sra_39_n125, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n97);
   dp_ex_stage_alu_shifter_sra_39_U8 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n74, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_n33, A => 
                           dp_ex_stage_alu_shifter_sra_39_n184, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n87);
   dp_ex_stage_alu_shifter_sra_39_U7 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n33, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n30, A => 
                           dp_ex_stage_alu_shifter_sra_39_n149, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n79);
   dp_ex_stage_alu_shifter_sra_39_U6 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n30, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_n231, A => 
                           dp_ex_stage_alu_shifter_sra_39_n181, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n123);
   dp_ex_stage_alu_shifter_sra_39_U5 : AOI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n113, B2 => 
                           dp_ex_stage_alu_n29, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n114, C2 => 
                           dp_ex_stage_alu_n38, A => 
                           dp_ex_stage_alu_shifter_sra_39_n56, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n151);
   dp_ex_stage_alu_shifter_sra_39_U4 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n38, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n39, A => 
                           dp_ex_stage_alu_shifter_sra_39_n165, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n86);
   dp_ex_stage_alu_shifter_sra_39_U3 : OAI221_X1 port map( B1 => 
                           dp_ex_stage_alu_shifter_sra_39_n76, B2 => 
                           dp_ex_stage_alu_shifter_sra_39_n43, C1 => 
                           dp_ex_stage_alu_shifter_sra_39_n74, C2 => 
                           dp_ex_stage_alu_shifter_sra_39_n68, A => 
                           dp_ex_stage_alu_shifter_sra_39_n180, ZN => 
                           dp_ex_stage_alu_shifter_sra_39_n138);
   dp_ex_stage_alu_shifter_sra_39_U2 : BUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_sra_39_n117, Z => 
                           dp_ex_stage_alu_shifter_sra_39_n11);
   dp_ex_stage_alu_shifter_rol_32_U16 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n31, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n10);
   dp_ex_stage_alu_shifter_rol_32_U15 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n31, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n11);
   dp_ex_stage_alu_shifter_rol_32_U14 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n31, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n12);
   dp_ex_stage_alu_shifter_rol_32_U13 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n49, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n7);
   dp_ex_stage_alu_shifter_rol_32_U12 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n49, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n8);
   dp_ex_stage_alu_shifter_rol_32_U11 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n49, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n9);
   dp_ex_stage_alu_shifter_rol_32_U10 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n4);
   dp_ex_stage_alu_shifter_rol_32_U9 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n5);
   dp_ex_stage_alu_shifter_rol_32_U8 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n6);
   dp_ex_stage_alu_shifter_rol_32_U7 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n3);
   dp_ex_stage_alu_shifter_rol_32_U6 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n2);
   dp_ex_stage_alu_shifter_rol_32_U5 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n1);
   dp_ex_stage_alu_shifter_rol_32_U4 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n15);
   dp_ex_stage_alu_shifter_rol_32_U3 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n13);
   dp_ex_stage_alu_shifter_rol_32_U2 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_rol_32_n14);
   dp_ex_stage_alu_shifter_rol_32_M0_0_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_N202, B => 
                           dp_ex_stage_alu_shifter_n1, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_0_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n76, B => 
                           dp_ex_stage_alu_shifter_N202, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_1_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n44, B => dp_ex_stage_alu_n76, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_2_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n69, B => dp_ex_stage_alu_n44, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_3_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n52, B => dp_ex_stage_alu_n69, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_4_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n70, B => dp_ex_stage_alu_n52, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_5_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n78, B => dp_ex_stage_alu_n70, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_6_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n34, B => dp_ex_stage_alu_n78, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_7_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n71, B => dp_ex_stage_alu_n34, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_8_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n72, B => dp_ex_stage_alu_n71, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_9_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n74, B => dp_ex_stage_alu_n72, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_10_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n33, B => dp_ex_stage_alu_n74, S => 
                           dp_ex_stage_alu_shifter_rol_32_n1, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_11_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_12_port, B => 
                           dp_ex_stage_alu_n33, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_12_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n231, B => 
                           dp_ex_stage_muxA_out_12_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_13_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_14_port, B => 
                           dp_ex_stage_alu_n231, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_14_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n29, B => 
                           dp_ex_stage_muxA_out_14_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_15_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n38, B => dp_ex_stage_alu_n29, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_16_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_17_port, B => 
                           dp_ex_stage_alu_n38, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_17_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_18_port, B => 
                           dp_ex_stage_muxA_out_17_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_18_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_19_port, B => 
                           dp_ex_stage_muxA_out_18_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_19_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_20_port, B => 
                           dp_ex_stage_muxA_out_19_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_20_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_21_port, B => 
                           dp_ex_stage_muxA_out_20_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_21_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n240, B => 
                           dp_ex_stage_muxA_out_21_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_22_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_23_port, B => 
                           dp_ex_stage_alu_n240, S => 
                           dp_ex_stage_alu_shifter_rol_32_n2, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_23_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n94, B => 
                           dp_ex_stage_muxA_out_23_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_24_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n7, B => 
                           dp_ex_stage_alu_shifter_n94, S => 
                           dp_ex_stage_alu_shifter_rol_32_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_25_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n11, B => 
                           dp_ex_stage_alu_shifter_n7, S => 
                           dp_ex_stage_alu_shifter_rol_32_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_26_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n12, B => 
                           dp_ex_stage_alu_shifter_n11, S => 
                           dp_ex_stage_alu_shifter_rol_32_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_27_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n1, B => dp_ex_stage_alu_shifter_n12
                           , S => dp_ex_stage_alu_shifter_rol_32_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_28_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_29_port, B => 
                           dp_ex_stage_alu_n1, S => 
                           dp_ex_stage_alu_shifter_rol_32_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_29_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_30_port, B => 
                           dp_ex_stage_muxA_out_29_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_30_port);
   dp_ex_stage_alu_shifter_rol_32_M1_0_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n1, B => 
                           dp_ex_stage_muxA_out_30_port, S => 
                           dp_ex_stage_alu_shifter_rol_32_n3, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_31_port);
   dp_ex_stage_alu_shifter_rol_32_M0_1_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_0_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_30_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_0_port);
   dp_ex_stage_alu_shifter_rol_32_M0_1_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_1_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_31_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_1_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_2_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_0_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_2_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_3_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_1_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_3_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_4_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_2_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_4_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_5_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_3_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_5_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_6_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_4_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_6_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_7_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_5_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_7_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_8_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_6_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_8_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_9_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_7_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_9_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_10_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_8_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_10_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_11_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_9_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n4, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_11_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_12_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_10_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_12_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_13_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_11_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_13_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_14_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_12_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_14_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_15_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_13_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_15_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_16_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_14_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_16_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_17_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_15_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_17_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_18_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_16_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_18_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_19_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_17_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_19_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_20_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_18_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_20_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_21_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_19_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_21_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_22_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_20_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_22_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_23_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_21_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n5, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_23_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_24_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_22_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n6, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_24_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_25_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_23_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n6, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_25_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_26_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_24_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n6, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_26_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_27_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_25_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n6, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_27_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_28_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_26_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n6, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_28_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_29_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_27_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n6, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_29_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_30_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_28_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n6, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_30_port);
   dp_ex_stage_alu_shifter_rol_32_M1_1_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_1_31_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_1_29_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n6, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_31_port);
   dp_ex_stage_alu_shifter_rol_32_M0_2_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_0_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_28_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_0_port);
   dp_ex_stage_alu_shifter_rol_32_M0_2_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_1_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_29_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_1_port);
   dp_ex_stage_alu_shifter_rol_32_M0_2_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_2_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_30_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_2_port);
   dp_ex_stage_alu_shifter_rol_32_M0_2_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_3_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_31_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_3_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_4_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_0_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_4_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_5_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_1_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_5_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_6_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_2_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_6_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_7_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_3_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_7_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_8_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_4_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_8_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_9_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_5_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_9_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_10_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_6_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_10_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_11_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_7_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n7, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_11_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_12_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_8_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_12_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_13_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_9_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_13_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_14_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_10_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_14_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_15_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_11_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_15_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_16_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_12_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_16_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_17_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_13_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_17_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_18_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_14_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_18_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_19_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_15_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_19_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_20_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_16_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_20_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_21_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_17_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_21_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_22_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_18_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_22_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_23_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_19_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n8, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_23_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_24_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_20_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n9, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_24_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_25_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_21_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n9, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_25_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_26_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_22_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n9, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_26_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_27_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_23_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n9, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_27_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_28_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_24_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n9, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_28_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_29_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_25_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n9, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_29_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_30_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_26_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n9, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_30_port);
   dp_ex_stage_alu_shifter_rol_32_M1_2_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_2_31_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_2_27_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n9, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_31_port);
   dp_ex_stage_alu_shifter_rol_32_M0_3_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_0_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_24_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_0_port);
   dp_ex_stage_alu_shifter_rol_32_M0_3_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_1_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_25_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_1_port);
   dp_ex_stage_alu_shifter_rol_32_M0_3_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_2_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_26_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_2_port);
   dp_ex_stage_alu_shifter_rol_32_M0_3_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_3_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_27_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_3_port);
   dp_ex_stage_alu_shifter_rol_32_M0_3_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_4_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_28_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_4_port);
   dp_ex_stage_alu_shifter_rol_32_M0_3_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_5_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_29_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_5_port);
   dp_ex_stage_alu_shifter_rol_32_M0_3_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_6_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_30_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_6_port);
   dp_ex_stage_alu_shifter_rol_32_M0_3_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_7_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_31_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_7_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_8_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_0_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_8_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_9_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_1_port, S =>
                           dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_9_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_10_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_2_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_10_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_11_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_3_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n10, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_11_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_12_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_4_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_12_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_13_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_5_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_13_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_14_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_6_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_14_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_15_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_7_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_15_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_16_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_8_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_16_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_17_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_9_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_17_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_18_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_10_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_18_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_19_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_11_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_19_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_20_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_12_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_20_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_21_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_13_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_21_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_22_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_14_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_22_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_23_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_15_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n11, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_23_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_24_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_16_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n12, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_24_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_25_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_17_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n12, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_25_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_26_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_18_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n12, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_26_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_27_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_19_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n12, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_27_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_28_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_20_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n12, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_28_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_29_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_21_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n12, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_29_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_30_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_22_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n12, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_30_port);
   dp_ex_stage_alu_shifter_rol_32_M1_3_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_3_31_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_3_23_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n12, Z => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_31_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_0_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_16_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N39_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_1_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_17_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N40_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_2_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_18_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N41_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_3_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_19_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N42_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_4_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_20_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N43_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_5_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_21_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N44_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_6_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_22_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N45_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_7_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_23_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N46_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_8_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_24_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N47_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_9_port, B =>
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_25_port, S 
                           => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N48_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_10_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_26_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N49_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_11_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_27_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n13, Z => 
                           dp_ex_stage_alu_shifter_N50_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_12_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_28_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N51_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_13_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_29_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N52_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_14_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_30_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N53_port);
   dp_ex_stage_alu_shifter_rol_32_M0_4_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_15_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_31_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N54_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_16_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_0_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N55_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_17_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_1_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N56_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_18_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_2_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N57_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_19_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_3_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N58_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_20_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_4_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N59_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_21_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_5_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N60_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_22_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_6_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N61_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_23_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_7_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n14, Z => 
                           dp_ex_stage_alu_shifter_N62_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_24_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_8_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n15, Z => 
                           dp_ex_stage_alu_shifter_N63_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_25_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_9_port, S
                           => dp_ex_stage_alu_shifter_rol_32_n15, Z => 
                           dp_ex_stage_alu_shifter_N64_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_26_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_10_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n15, Z => 
                           dp_ex_stage_alu_shifter_N65_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_27_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_11_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n15, Z => 
                           dp_ex_stage_alu_shifter_N66_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_28_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_12_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n15, Z => 
                           dp_ex_stage_alu_shifter_N67_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_29_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_13_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n15, Z => 
                           dp_ex_stage_alu_shifter_N68_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_30_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_14_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n15, Z => 
                           dp_ex_stage_alu_shifter_N69_port);
   dp_ex_stage_alu_shifter_rol_32_M1_4_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_rol_32_ML_int_4_31_port, B 
                           => dp_ex_stage_alu_shifter_rol_32_ML_int_4_15_port, 
                           S => dp_ex_stage_alu_shifter_rol_32_n15, Z => 
                           dp_ex_stage_alu_shifter_N70_port);
   dp_ex_stage_alu_shifter_ror_30_U16 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n31, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n10);
   dp_ex_stage_alu_shifter_ror_30_U15 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n31, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n11);
   dp_ex_stage_alu_shifter_ror_30_U14 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n31, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n12);
   dp_ex_stage_alu_shifter_ror_30_U13 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n49, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n7);
   dp_ex_stage_alu_shifter_ror_30_U12 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n49, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n8);
   dp_ex_stage_alu_shifter_ror_30_U11 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_n49, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n9);
   dp_ex_stage_alu_shifter_ror_30_U10 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n4);
   dp_ex_stage_alu_shifter_ror_30_U9 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n5);
   dp_ex_stage_alu_shifter_ror_30_U8 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n6);
   dp_ex_stage_alu_shifter_ror_30_U7 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n3);
   dp_ex_stage_alu_shifter_ror_30_U6 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n1);
   dp_ex_stage_alu_shifter_ror_30_U5 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n2);
   dp_ex_stage_alu_shifter_ror_30_U4 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n15);
   dp_ex_stage_alu_shifter_ror_30_U3 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n13);
   dp_ex_stage_alu_shifter_ror_30_U2 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n116, Z => 
                           dp_ex_stage_alu_shifter_ror_30_n14);
   dp_ex_stage_alu_shifter_ror_30_M1_0_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_N202, B => 
                           dp_ex_stage_alu_n76, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_0_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_1_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n76, B => dp_ex_stage_alu_n44, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_1_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_2_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n44, B => dp_ex_stage_alu_n69, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_2_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_3_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n69, B => dp_ex_stage_alu_n52, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_3_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_4_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n52, B => dp_ex_stage_alu_n70, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_4_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_5_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n70, B => dp_ex_stage_alu_n78, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_5_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_6_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n78, B => dp_ex_stage_alu_n34, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_6_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_7_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n34, B => dp_ex_stage_alu_n71, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_7_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_8_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n71, B => dp_ex_stage_alu_n72, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_8_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_9_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n72, B => dp_ex_stage_alu_n74, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_9_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_10_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n74, B => dp_ex_stage_alu_n33, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_10_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_11_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n33, B => 
                           dp_ex_stage_muxA_out_12_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n1, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_11_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_12_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_12_port, B => 
                           dp_ex_stage_alu_n231, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_12_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_13_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n231, B => 
                           dp_ex_stage_muxA_out_14_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_13_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_14_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_14_port, B => 
                           dp_ex_stage_alu_n29, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_14_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_15_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n29, B => dp_ex_stage_alu_n38, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_15_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_16_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n38, B => 
                           dp_ex_stage_muxA_out_17_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_16_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_17_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_17_port, B => 
                           dp_ex_stage_muxA_out_18_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_17_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_18_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_18_port, B => 
                           dp_ex_stage_muxA_out_19_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_18_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_19_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_19_port, B => 
                           dp_ex_stage_muxA_out_20_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_19_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_20_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_20_port, B => 
                           dp_ex_stage_muxA_out_21_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_20_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_21_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_21_port, B => 
                           dp_ex_stage_alu_n240, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_21_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_22_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n240, B => 
                           dp_ex_stage_muxA_out_23_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_22_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_23_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_23_port, B => 
                           dp_ex_stage_alu_shifter_n94, S => 
                           dp_ex_stage_alu_shifter_ror_30_n2, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_23_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_24_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n94, B => 
                           dp_ex_stage_alu_shifter_n7, S => 
                           dp_ex_stage_alu_shifter_ror_30_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_24_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_25_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n7, B => 
                           dp_ex_stage_alu_shifter_n11, S => 
                           dp_ex_stage_alu_shifter_ror_30_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_25_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_26_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n11, B => 
                           dp_ex_stage_alu_shifter_n12, S => 
                           dp_ex_stage_alu_shifter_ror_30_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_26_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_27_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n12, B => dp_ex_stage_alu_n1
                           , S => dp_ex_stage_alu_shifter_ror_30_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_27_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_28_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_n1, B => 
                           dp_ex_stage_muxA_out_29_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_28_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_29_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_29_port, B => 
                           dp_ex_stage_muxA_out_30_port, S => 
                           dp_ex_stage_alu_shifter_ror_30_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_29_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_30_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_muxA_out_30_port, B => 
                           dp_ex_stage_alu_shifter_n1, S => 
                           dp_ex_stage_alu_shifter_ror_30_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_30_port);
   dp_ex_stage_alu_shifter_ror_30_M1_0_31_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_n1, B => 
                           dp_ex_stage_alu_shifter_N202, S => 
                           dp_ex_stage_alu_shifter_ror_30_n3, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_31_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_0_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_2_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_0_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_1_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_3_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_1_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_2_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_2_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_4_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_2_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_3_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_3_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_5_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_3_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_4_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_4_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_6_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_4_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_5_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_5_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_7_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_5_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_6_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_6_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_8_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_6_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_7_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_7_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_9_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_7_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_8_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_8_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_10_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_8_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_9_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_9_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_11_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_9_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_10_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_10_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_12_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_10_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_11_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_11_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_13_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n4, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_11_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_12_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_12_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_14_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_12_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_13_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_13_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_15_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_13_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_14_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_14_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_16_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_14_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_15_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_15_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_17_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_15_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_16_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_16_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_18_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_16_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_17_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_17_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_19_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_17_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_18_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_18_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_20_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_18_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_19_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_19_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_21_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_19_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_20_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_20_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_22_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_20_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_21_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_21_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_23_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_21_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_22_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_22_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_24_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_22_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_23_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_23_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_25_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n5, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_23_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_24_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_24_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_26_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n6, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_24_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_25_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_25_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_27_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n6, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_25_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_26_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_26_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_28_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n6, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_26_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_27_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_27_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_29_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n6, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_27_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_28_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_28_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_30_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n6, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_28_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_29_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_29_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_31_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n6, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_29_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_30_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_30_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_0_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n6, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_30_port);
   dp_ex_stage_alu_shifter_ror_30_M1_1_31_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_1_31_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_1_1_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n6, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_31_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_0_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_4_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_0_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_1_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_5_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_1_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_2_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_6_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_2_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_3_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_7_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_3_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_4_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_4_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_8_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_4_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_5_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_5_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_9_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_5_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_6_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_6_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_10_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_6_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_7_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_7_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_11_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_7_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_8_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_8_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_12_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_8_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_9_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_9_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_13_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_9_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_10_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_10_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_14_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_10_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_11_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_11_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_15_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n7, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_11_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_12_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_12_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_16_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_12_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_13_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_13_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_17_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_13_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_14_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_14_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_18_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_14_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_15_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_15_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_19_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_15_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_16_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_16_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_20_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_16_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_17_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_17_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_21_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_17_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_18_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_18_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_22_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_18_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_19_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_19_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_23_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_19_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_20_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_20_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_24_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_20_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_21_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_21_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_25_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_21_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_22_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_22_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_26_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_22_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_23_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_23_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_27_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n8, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_23_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_24_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_24_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_28_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n9, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_24_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_25_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_25_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_29_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n9, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_25_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_26_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_26_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_30_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n9, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_26_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_27_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_27_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_31_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n9, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_27_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_28_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_28_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_0_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n9, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_28_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_29_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_29_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_1_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n9, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_29_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_30_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_30_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_2_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n9, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_30_port);
   dp_ex_stage_alu_shifter_ror_30_M1_2_31_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_2_31_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_2_3_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n9, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_31_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_0_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_8_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_0_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_1_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_9_port, S =>
                           dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_1_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_2_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_10_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_2_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_3_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_11_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_3_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_4_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_12_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_4_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_5_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_13_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_5_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_6_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_14_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_6_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_7_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_15_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_7_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_8_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_8_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_16_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_8_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_9_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_9_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_17_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_9_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_10_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_10_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_18_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_10_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_11_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_11_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_19_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n10, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_11_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_12_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_12_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_20_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_12_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_13_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_13_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_21_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_13_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_14_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_14_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_22_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_14_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_15_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_15_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_23_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_15_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_16_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_16_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_24_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_16_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_17_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_17_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_25_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_17_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_18_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_18_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_26_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_18_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_19_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_19_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_27_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_19_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_20_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_20_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_28_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_20_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_21_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_21_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_29_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_21_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_22_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_22_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_30_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_22_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_23_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_23_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_31_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n11, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_23_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_24_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_24_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_0_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n12, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_24_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_25_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_25_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_1_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n12, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_25_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_26_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_26_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_2_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n12, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_26_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_27_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_27_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_3_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n12, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_27_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_28_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_28_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_4_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n12, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_28_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_29_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_29_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_5_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n12, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_29_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_30_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_30_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_6_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n12, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_30_port);
   dp_ex_stage_alu_shifter_ror_30_M1_3_31_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_3_31_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_3_7_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n12, Z => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_31_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_0 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_0_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_16_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N7_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_1 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_1_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_17_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N8_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_2 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_2_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_18_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N9_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_3 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_3_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_19_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N10_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_4 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_4_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_20_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N11_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_5 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_5_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_21_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N12_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_6 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_6_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_22_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N13_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_7 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_7_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_23_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N14_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_8 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_8_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_24_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N15_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_9 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_9_port, B =>
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_25_port, S 
                           => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N16_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_10 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_10_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_26_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N17_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_11 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_11_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_27_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n13, Z => 
                           dp_ex_stage_alu_shifter_N18_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_12 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_12_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_28_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N19_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_13 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_13_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_29_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N20_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_14 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_14_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_30_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N21_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_15 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_15_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_31_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N22_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_16 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_16_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_0_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N23_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_17 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_17_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_1_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N24_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_18 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_18_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_2_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N25_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_19 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_19_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_3_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N26_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_20 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_20_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_4_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N27_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_21 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_21_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_5_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N28_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_22 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_22_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_6_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N29_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_23 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_23_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_7_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n14, Z => 
                           dp_ex_stage_alu_shifter_N30_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_24 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_24_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_8_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n15, Z => 
                           dp_ex_stage_alu_shifter_N31_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_25 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_25_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_9_port, S
                           => dp_ex_stage_alu_shifter_ror_30_n15, Z => 
                           dp_ex_stage_alu_shifter_N32_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_26 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_26_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_10_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n15, Z => 
                           dp_ex_stage_alu_shifter_N33_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_27 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_27_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_11_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n15, Z => 
                           dp_ex_stage_alu_shifter_N34_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_28 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_28_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_12_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n15, Z => 
                           dp_ex_stage_alu_shifter_N35_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_29 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_29_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_13_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n15, Z => 
                           dp_ex_stage_alu_shifter_N36_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_30 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_30_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_14_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n15, Z => 
                           dp_ex_stage_alu_shifter_N37_port);
   dp_ex_stage_alu_shifter_ror_30_M1_4_31 : MUX2_X1 port map( A => 
                           dp_ex_stage_alu_shifter_ror_30_MR_int_4_31_port, B 
                           => dp_ex_stage_alu_shifter_ror_30_MR_int_4_15_port, 
                           S => dp_ex_stage_alu_shifter_ror_30_n15, Z => 
                           dp_ex_stage_alu_shifter_N38_port);
   dp_ex_stage_alu_r61_U225 : INV_X1 port map( A => dp_ex_stage_alu_r61_n91, ZN
                           => dp_ex_stage_alu_r61_n218);
   dp_ex_stage_alu_r61_U224 : INV_X1 port map( A => dp_ex_stage_alu_r61_n51, ZN
                           => dp_ex_stage_alu_r61_n219);
   dp_ex_stage_alu_r61_U223 : INV_X1 port map( A => dp_ex_stage_alu_r61_n45, ZN
                           => dp_ex_stage_alu_r61_n216);
   dp_ex_stage_alu_r61_U222 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r61_n155
                           , A2 => dp_ex_stage_alu_r61_n147, A3 => 
                           dp_ex_stage_alu_r61_n216, ZN => 
                           dp_ex_stage_alu_r61_n212);
   dp_ex_stage_alu_r61_U221 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r61_n211
                           , A2 => dp_ex_stage_alu_r61_n212, A3 => 
                           dp_ex_stage_alu_r61_n213, ZN => 
                           dp_ex_stage_alu_r61_n122);
   dp_ex_stage_alu_r61_U220 : INV_X1 port map( A => dp_ex_stage_alu_r61_n75, ZN
                           => dp_ex_stage_alu_r61_n207);
   dp_ex_stage_alu_r61_U219 : INV_X1 port map( A => dp_ex_stage_alu_r61_n88, ZN
                           => dp_ex_stage_alu_r61_n208);
   dp_ex_stage_alu_r61_U218 : INV_X1 port map( A => dp_ex_stage_alu_r61_n82, ZN
                           => dp_ex_stage_alu_r61_n204);
   dp_ex_stage_alu_r61_U217 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r61_n186
                           , A2 => dp_ex_stage_alu_r61_n193, A3 => 
                           dp_ex_stage_alu_r61_n204, ZN => 
                           dp_ex_stage_alu_r61_n202);
   dp_ex_stage_alu_r61_U216 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r61_n201
                           , A2 => dp_ex_stage_alu_r61_n202, A3 => 
                           dp_ex_stage_alu_r61_n203, ZN => 
                           dp_ex_stage_alu_r61_n166);
   dp_ex_stage_alu_r61_U215 : INV_X1 port map( A => dp_ex_stage_alu_r61_n193, 
                           ZN => dp_ex_stage_alu_r61_n192);
   dp_ex_stage_alu_r61_U214 : INV_X1 port map( A => dp_ex_stage_alu_r61_n161, 
                           ZN => dp_ex_stage_alu_r61_n179);
   dp_ex_stage_alu_r61_U213 : INV_X1 port map( A => dp_ex_stage_alu_r61_n87, ZN
                           => dp_ex_stage_alu_r61_n164);
   dp_ex_stage_alu_r61_U212 : INV_X1 port map( A => dp_ex_stage_alu_r61_n92, ZN
                           => dp_ex_stage_alu_r61_n165);
   dp_ex_stage_alu_r61_U211 : INV_X1 port map( A => dp_ex_stage_alu_r61_n86, ZN
                           => dp_ex_stage_alu_r61_n163);
   dp_ex_stage_alu_r61_U210 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r61_n2, 
                           A2 => dp_ex_stage_alu_r61_n162, A3 => 
                           dp_ex_stage_alu_r61_n163, ZN => 
                           dp_ex_stage_alu_r61_n157);
   dp_ex_stage_alu_r61_U209 : INV_X1 port map( A => dp_ex_stage_alu_r61_n93, ZN
                           => dp_ex_stage_alu_r61_n160);
   dp_ex_stage_alu_r61_U208 : INV_X1 port map( A => dp_ex_stage_alu_r61_n155, 
                           ZN => dp_ex_stage_alu_r61_n154);
   dp_ex_stage_alu_r61_U207 : INV_X1 port map( A => dp_ex_stage_alu_r61_n147, 
                           ZN => dp_ex_stage_alu_r61_n146);
   dp_ex_stage_alu_r61_U206 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r61_n142
                           , A2 => dp_ex_stage_alu_r61_n143, A3 => 
                           dp_ex_stage_alu_r61_n144, ZN => 
                           dp_ex_stage_alu_r61_n141);
   dp_ex_stage_alu_r61_U205 : INV_X1 port map( A => dp_ex_stage_alu_r61_n117, 
                           ZN => dp_ex_stage_alu_r61_n137);
   dp_ex_stage_alu_r61_U204 : INV_X1 port map( A => dp_ex_stage_alu_r61_n118, 
                           ZN => dp_ex_stage_alu_r61_n129);
   dp_ex_stage_alu_r61_U203 : INV_X1 port map( A => dp_ex_stage_alu_r61_n50, ZN
                           => dp_ex_stage_alu_r61_n121);
   dp_ex_stage_alu_r61_U202 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n117
                           , A2 => dp_ex_stage_alu_r61_n121, ZN => 
                           dp_ex_stage_alu_r61_n119);
   dp_ex_stage_alu_r61_U201 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n119
                           , A2 => dp_ex_stage_alu_r61_n120, ZN => 
                           dp_ex_stage_alu_r61_n114);
   dp_ex_stage_alu_r61_U200 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n97,
                           A2 => dp_ex_stage_alu_r61_n98, ZN => 
                           dp_ex_stage_alu_r61_n96);
   dp_ex_stage_alu_r61_U199 : NAND4_X1 port map( A1 => dp_ex_stage_alu_r61_n67,
                           A2 => dp_ex_stage_alu_r61_n68, A3 => 
                           dp_ex_stage_alu_r61_n69, A4 => 
                           dp_ex_stage_alu_r61_n70, ZN => 
                           dp_ex_stage_alu_r61_n34);
   dp_ex_stage_alu_r61_U198 : XNOR2_X1 port map( A => 
                           dp_ex_stage_muxB_out_31_port, B => 
                           dp_ex_stage_alu_r61_n31, ZN => 
                           dp_ex_stage_alu_r61_n60);
   dp_ex_stage_alu_r61_U197 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n60,
                           A2 => dp_ex_stage_alu_r61_n61, ZN => 
                           dp_ex_stage_alu_r61_n59);
   dp_ex_stage_alu_r61_U196 : INV_X1 port map( A => dp_ex_stage_alu_N18_port, 
                           ZN => dp_ex_stage_alu_N19_port);
   dp_ex_stage_alu_r61_U195 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_31_port, ZN => 
                           dp_ex_stage_alu_r61_n32);
   dp_ex_stage_alu_r61_U194 : INV_X1 port map( A => dp_ex_stage_alu_r61_n32, ZN
                           => dp_ex_stage_alu_r61_n31);
   dp_ex_stage_alu_r61_U193 : INV_X1 port map( A => dp_ex_stage_alu_n247, ZN =>
                           dp_ex_stage_alu_r61_n30);
   dp_ex_stage_alu_r61_U192 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_27_port, ZN => 
                           dp_ex_stage_alu_r61_n29);
   dp_ex_stage_alu_r61_U191 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_26_port, ZN => 
                           dp_ex_stage_alu_r61_n28);
   dp_ex_stage_alu_r61_U190 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_25_port, ZN => 
                           dp_ex_stage_alu_r61_n27);
   dp_ex_stage_alu_r61_U189 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_24_port, ZN => 
                           dp_ex_stage_alu_r61_n26);
   dp_ex_stage_alu_r61_U188 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_23_port, ZN => 
                           dp_ex_stage_alu_r61_n25);
   dp_ex_stage_alu_r61_U187 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_22_port, ZN => 
                           dp_ex_stage_alu_r61_n24);
   dp_ex_stage_alu_r61_U186 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_21_port, ZN => 
                           dp_ex_stage_alu_r61_n23);
   dp_ex_stage_alu_r61_U185 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_18_port, ZN => 
                           dp_ex_stage_alu_r61_n22);
   dp_ex_stage_alu_r61_U184 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_17_port, ZN => 
                           dp_ex_stage_alu_r61_n21);
   dp_ex_stage_alu_r61_U183 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_16_port, ZN => 
                           dp_ex_stage_alu_r61_n20);
   dp_ex_stage_alu_r61_U182 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_15_port, ZN => 
                           dp_ex_stage_alu_r61_n19);
   dp_ex_stage_alu_r61_U181 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_14_port, ZN => 
                           dp_ex_stage_alu_r61_n18);
   dp_ex_stage_alu_r61_U180 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_13_port, ZN => 
                           dp_ex_stage_alu_r61_n17);
   dp_ex_stage_alu_r61_U179 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_12_port, ZN => 
                           dp_ex_stage_alu_r61_n16);
   dp_ex_stage_alu_r61_U178 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_11_port, ZN => 
                           dp_ex_stage_alu_r61_n15);
   dp_ex_stage_alu_r61_U177 : INV_X1 port map( A => dp_ex_stage_alu_n30, ZN => 
                           dp_ex_stage_alu_r61_n14);
   dp_ex_stage_alu_r61_U176 : INV_X1 port map( A => dp_ex_stage_muxA_out_9_port
                           , ZN => dp_ex_stage_alu_r61_n13);
   dp_ex_stage_alu_r61_U175 : INV_X1 port map( A => dp_ex_stage_muxA_out_8_port
                           , ZN => dp_ex_stage_alu_r61_n12);
   dp_ex_stage_alu_r61_U174 : INV_X1 port map( A => dp_ex_stage_muxA_out_7_port
                           , ZN => dp_ex_stage_alu_r61_n11);
   dp_ex_stage_alu_r61_U173 : INV_X1 port map( A => dp_ex_stage_muxA_out_3_port
                           , ZN => dp_ex_stage_alu_r61_n10);
   dp_ex_stage_alu_r61_U172 : INV_X1 port map( A => dp_ex_stage_muxA_out_2_port
                           , ZN => dp_ex_stage_alu_r61_n9);
   dp_ex_stage_alu_r61_U171 : INV_X1 port map( A => dp_ex_stage_alu_n22, ZN => 
                           dp_ex_stage_alu_r61_n8);
   dp_ex_stage_alu_r61_U170 : INV_X1 port map( A => dp_ex_stage_alu_n50, ZN => 
                           dp_ex_stage_alu_r61_n7);
   dp_ex_stage_alu_r61_U169 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n77, A2 
                           => dp_ex_stage_alu_r61_n10, ZN => 
                           dp_ex_stage_alu_r61_n76);
   dp_ex_stage_alu_r61_U168 : NOR2_X1 port map( A1 => dp_ex_stage_alu_n77, A2 
                           => dp_ex_stage_alu_r61_n10, ZN => 
                           dp_ex_stage_alu_r61_n187);
   dp_ex_stage_alu_r61_U167 : NOR2_X1 port map( A1 => dp_ex_stage_alu_n46, A2 
                           => dp_ex_stage_alu_r61_n66, ZN => 
                           dp_ex_stage_alu_r61_n199);
   dp_ex_stage_alu_r61_U166 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n46, A2 
                           => dp_ex_stage_alu_r61_n66, ZN => 
                           dp_ex_stage_alu_r61_n200);
   dp_ex_stage_alu_r61_U165 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n46, A2 
                           => dp_ex_stage_alu_r61_n66, ZN => 
                           dp_ex_stage_alu_r61_n63);
   dp_ex_stage_alu_r61_U164 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r61_n167
                           , B2 => dp_ex_stage_alu_r61_n166, A => 
                           dp_ex_stage_alu_r61_n168, ZN => 
                           dp_ex_stage_alu_r61_n139);
   dp_ex_stage_alu_r61_U163 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r61_n139
                           , B2 => dp_ex_stage_alu_r61_n140, A => 
                           dp_ex_stage_alu_r61_n141, ZN => 
                           dp_ex_stage_alu_r61_n123);
   dp_ex_stage_alu_r61_U162 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r61_n123
                           , B2 => dp_ex_stage_alu_r61_n122, A => 
                           dp_ex_stage_alu_r61_n124, ZN => 
                           dp_ex_stage_alu_r61_n107);
   dp_ex_stage_alu_r61_U161 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r61_n107
                           , B2 => dp_ex_stage_alu_r61_n108, A => 
                           dp_ex_stage_alu_r61_n109, ZN => 
                           dp_ex_stage_alu_r61_n102);
   dp_ex_stage_alu_r61_U160 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n30, A2 
                           => dp_ex_stage_alu_r61_n176, ZN => 
                           dp_ex_stage_alu_r61_n173);
   dp_ex_stage_alu_r61_U159 : INV_X1 port map( A => dp_ex_stage_alu_n23, ZN => 
                           dp_ex_stage_alu_r61_n197);
   dp_ex_stage_alu_r61_U158 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n23, A2 
                           => dp_ex_stage_alu_r61_n8, ZN => 
                           dp_ex_stage_alu_r61_n194);
   dp_ex_stage_alu_r61_U157 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n50, A2 
                           => dp_ex_stage_alu_r61_n9, ZN => 
                           dp_ex_stage_alu_r61_n73);
   dp_ex_stage_alu_r61_U156 : INV_X1 port map( A => dp_ex_stage_muxA_out_6_port
                           , ZN => dp_ex_stage_alu_r61_n209);
   dp_ex_stage_alu_r61_U155 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_6_port, A2 => 
                           dp_ex_stage_alu_r61_n206, ZN => 
                           dp_ex_stage_alu_r61_n193);
   dp_ex_stage_alu_r61_U154 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_30_port, A2 => 
                           dp_ex_stage_alu_r61_n62, ZN => 
                           dp_ex_stage_alu_r61_n100);
   dp_ex_stage_alu_r61_U153 : AND3_X1 port map( A1 => dp_ex_stage_alu_r61_n99, 
                           A2 => dp_ex_stage_alu_r61_n100, A3 => 
                           dp_ex_stage_alu_r61_n54, ZN => 
                           dp_ex_stage_alu_r61_n98);
   dp_ex_stage_alu_r61_U152 : INV_X1 port map( A => dp_ex_stage_muxB_out_5_port
                           , ZN => dp_ex_stage_alu_r61_n196);
   dp_ex_stage_alu_r61_U151 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_5_port, A2 => 
                           dp_ex_stage_alu_r61_n196, ZN => 
                           dp_ex_stage_alu_r61_n195);
   dp_ex_stage_alu_r61_U150 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n194
                           , A2 => dp_ex_stage_alu_r61_n195, ZN => 
                           dp_ex_stage_alu_r61_n191);
   dp_ex_stage_alu_r61_U149 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_27_port, ZN => 
                           dp_ex_stage_alu_r61_n113);
   dp_ex_stage_alu_r61_U148 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_26_port, A2 => 
                           dp_ex_stage_alu_r61_n112, ZN => 
                           dp_ex_stage_alu_r61_n111);
   dp_ex_stage_alu_r61_U147 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_27_port, A2 => 
                           dp_ex_stage_alu_r61_n113, ZN => 
                           dp_ex_stage_alu_r61_n110);
   dp_ex_stage_alu_r61_U146 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n110
                           , A2 => dp_ex_stage_alu_r61_n111, ZN => 
                           dp_ex_stage_alu_r61_n109);
   dp_ex_stage_alu_r61_U145 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_10_port, ZN => 
                           dp_ex_stage_alu_r61_n176);
   dp_ex_stage_alu_r61_U144 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_30_port, A2 => 
                           dp_ex_stage_alu_r61_n62, ZN => 
                           dp_ex_stage_alu_r61_n222);
   dp_ex_stage_alu_r61_U143 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_22_port, ZN => 
                           dp_ex_stage_alu_r61_n134);
   dp_ex_stage_alu_r61_U142 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_26_port, ZN => 
                           dp_ex_stage_alu_r61_n112);
   dp_ex_stage_alu_r61_U141 : INV_X1 port map( A => dp_ex_stage_muxA_out_1_port
                           , ZN => dp_ex_stage_alu_r61_n66);
   dp_ex_stage_alu_r61_U140 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_31_port, A2 => 
                           dp_ex_stage_alu_r61_n32, ZN => 
                           dp_ex_stage_alu_r61_n221);
   dp_ex_stage_alu_r61_U139 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n221,
                           A2 => dp_ex_stage_alu_r61_n1, ZN => 
                           dp_ex_stage_alu_r61_n95);
   dp_ex_stage_alu_r61_U138 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_6_port, A2 => 
                           dp_ex_stage_alu_r61_n209, ZN => 
                           dp_ex_stage_alu_r61_n75);
   dp_ex_stage_alu_r61_U137 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_7_port, A2 => 
                           dp_ex_stage_alu_r61_n11, ZN => 
                           dp_ex_stage_alu_r61_n80);
   dp_ex_stage_alu_r61_U136 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_8_port, A2 => 
                           dp_ex_stage_alu_r61_n12, ZN => 
                           dp_ex_stage_alu_r61_n81);
   dp_ex_stage_alu_r61_U135 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_17_port, ZN => 
                           dp_ex_stage_alu_r61_n150);
   dp_ex_stage_alu_r61_U134 : INV_X1 port map( A => dp_ex_stage_alu_n21, ZN => 
                           dp_ex_stage_alu_r61_n65);
   dp_ex_stage_alu_r61_U133 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n145,
                           A2 => dp_ex_stage_alu_r61_n146, ZN => 
                           dp_ex_stage_alu_r61_n144);
   dp_ex_stage_alu_r61_U132 : NAND4_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_14_port, A2 => 
                           dp_ex_stage_alu_r61_n92, A3 => 
                           dp_ex_stage_alu_r61_n93, A4 => 
                           dp_ex_stage_alu_r61_n152, ZN => 
                           dp_ex_stage_alu_r61_n143);
   dp_ex_stage_alu_r61_U131 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r61_n153
                           , B2 => dp_ex_stage_alu_r61_n93, A => 
                           dp_ex_stage_alu_r61_n154, ZN => 
                           dp_ex_stage_alu_r61_n142);
   dp_ex_stage_alu_r61_U130 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n173,
                           A2 => dp_ex_stage_alu_r61_n174, ZN => 
                           dp_ex_stage_alu_r61_n6);
   dp_ex_stage_alu_r61_U129 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n6, 
                           A2 => dp_ex_stage_alu_r61_n162, ZN => 
                           dp_ex_stage_alu_r61_n171);
   dp_ex_stage_alu_r61_U128 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_14_port, ZN => 
                           dp_ex_stage_alu_r61_n152);
   dp_ex_stage_alu_r61_U127 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_16_port, ZN => 
                           dp_ex_stage_alu_r61_n151);
   dp_ex_stage_alu_r61_U126 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_17_port, A2 => 
                           dp_ex_stage_alu_r61_n150, ZN => 
                           dp_ex_stage_alu_r61_n149);
   dp_ex_stage_alu_r61_U125 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_16_port, A2 => 
                           dp_ex_stage_alu_r61_n151, ZN => 
                           dp_ex_stage_alu_r61_n148);
   dp_ex_stage_alu_r61_U124 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n148
                           , A2 => dp_ex_stage_alu_r61_n149, ZN => 
                           dp_ex_stage_alu_r61_n145);
   dp_ex_stage_alu_r61_U123 : INV_X1 port map( A => dp_ex_stage_muxB_out_6_port
                           , ZN => dp_ex_stage_alu_r61_n206);
   dp_ex_stage_alu_r61_U122 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_26_port, A2 => 
                           dp_ex_stage_alu_r61_n28, ZN => 
                           dp_ex_stage_alu_r61_n48);
   dp_ex_stage_alu_r61_U121 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_25_port, A2 => 
                           dp_ex_stage_alu_r61_n27, ZN => 
                           dp_ex_stage_alu_r61_n57);
   dp_ex_stage_alu_r61_U120 : INV_X1 port map( A => dp_ex_stage_muxB_out_7_port
                           , ZN => dp_ex_stage_alu_r61_n210);
   dp_ex_stage_alu_r61_U119 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_7_port, A2 => 
                           dp_ex_stage_alu_r61_n210, ZN => 
                           dp_ex_stage_alu_r61_n186);
   dp_ex_stage_alu_r61_U118 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_18_port, A2 => 
                           dp_ex_stage_alu_r61_n22, ZN => 
                           dp_ex_stage_alu_r61_n91);
   dp_ex_stage_alu_r61_U117 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_24_port, A2 => 
                           dp_ex_stage_alu_r61_n26, ZN => 
                           dp_ex_stage_alu_r61_n50);
   dp_ex_stage_alu_r61_U116 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_29_port, A2 => 
                           dp_ex_stage_alu_r61_n101, ZN => 
                           dp_ex_stage_alu_r61_n54);
   dp_ex_stage_alu_r61_U115 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_30_port, A2 => 
                           dp_ex_stage_alu_r61_n62, ZN => 
                           dp_ex_stage_alu_r61_n61);
   dp_ex_stage_alu_r61_U114 : INV_X1 port map( A => dp_ex_stage_muxA_out_5_port
                           , ZN => dp_ex_stage_alu_r61_n205);
   dp_ex_stage_alu_r61_U113 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_5_port, A2 => 
                           dp_ex_stage_alu_r61_n205, ZN => 
                           dp_ex_stage_alu_r61_n82);
   dp_ex_stage_alu_r61_U112 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_11_port, A2 => 
                           dp_ex_stage_alu_r61_n15, ZN => 
                           dp_ex_stage_alu_r61_n86);
   dp_ex_stage_alu_r61_U111 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_20_port, ZN => 
                           dp_ex_stage_alu_r61_n215);
   dp_ex_stage_alu_r61_U110 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_20_port, A2 => 
                           dp_ex_stage_alu_r61_n215, ZN => 
                           dp_ex_stage_alu_r61_n44);
   dp_ex_stage_alu_r61_U109 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_27_port, A2 => 
                           dp_ex_stage_alu_r61_n29, ZN => 
                           dp_ex_stage_alu_r61_n55);
   dp_ex_stage_alu_r61_U108 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_23_port, A2 => 
                           dp_ex_stage_alu_r61_n25, ZN => 
                           dp_ex_stage_alu_r61_n49);
   dp_ex_stage_alu_r61_U107 : INV_X1 port map( A => dp_ex_stage_muxB_out_8_port
                           , ZN => dp_ex_stage_alu_r61_n177);
   dp_ex_stage_alu_r61_U106 : NAND4_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_8_port, A2 => 
                           dp_ex_stage_alu_r61_n88, A3 => 
                           dp_ex_stage_alu_r61_n79, A4 => 
                           dp_ex_stage_alu_r61_n177, ZN => 
                           dp_ex_stage_alu_r61_n170);
   dp_ex_stage_alu_r61_U105 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_14_port, A2 => 
                           dp_ex_stage_alu_r61_n18, ZN => 
                           dp_ex_stage_alu_r61_n85);
   dp_ex_stage_alu_r61_U104 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_15_port, A2 => 
                           dp_ex_stage_alu_r61_n19, ZN => 
                           dp_ex_stage_alu_r61_n153);
   dp_ex_stage_alu_r61_U103 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_13_port, A2 => 
                           dp_ex_stage_alu_r61_n17, ZN => 
                           dp_ex_stage_alu_r61_n94);
   dp_ex_stage_alu_r61_U102 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_28_port, A2 => 
                           dp_ex_stage_alu_r61_n30, ZN => 
                           dp_ex_stage_alu_r61_n105);
   dp_ex_stage_alu_r61_U101 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_28_port, A2 => 
                           dp_ex_stage_alu_r61_n30, ZN => 
                           dp_ex_stage_alu_r61_n56);
   dp_ex_stage_alu_r61_U100 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_21_port, A2 => 
                           dp_ex_stage_alu_r61_n23, ZN => 
                           dp_ex_stage_alu_r61_n136);
   dp_ex_stage_alu_r61_U99 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r61_n136,
                           B2 => dp_ex_stage_alu_r61_n42, A => 
                           dp_ex_stage_alu_r61_n137, ZN => 
                           dp_ex_stage_alu_r61_n125);
   dp_ex_stage_alu_r61_U98 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_29_port, A2 => 
                           dp_ex_stage_alu_r61_n101, ZN => 
                           dp_ex_stage_alu_r61_n106);
   dp_ex_stage_alu_r61_U97 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_9_port, A2 => 
                           dp_ex_stage_alu_r61_n13, ZN => 
                           dp_ex_stage_alu_r61_n178);
   dp_ex_stage_alu_r61_U96 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r61_n178,
                           B2 => dp_ex_stage_alu_r61_n79, A => 
                           dp_ex_stage_alu_r61_n179, ZN => 
                           dp_ex_stage_alu_r61_n169);
   dp_ex_stage_alu_r61_U95 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_21_port, A2 => 
                           dp_ex_stage_alu_r61_n23, ZN => 
                           dp_ex_stage_alu_r61_n51);
   dp_ex_stage_alu_r61_U94 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n45, A2 
                           => dp_ex_stage_alu_r61_n65, ZN => 
                           dp_ex_stage_alu_r61_n64);
   dp_ex_stage_alu_r61_U93 : NOR2_X1 port map( A1 => dp_ex_stage_alu_n45, A2 =>
                           dp_ex_stage_alu_r61_n65, ZN => 
                           dp_ex_stage_alu_r61_n198);
   dp_ex_stage_alu_r61_U92 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_9_port, A2 => 
                           dp_ex_stage_alu_r61_n13, ZN => 
                           dp_ex_stage_alu_r61_n88);
   dp_ex_stage_alu_r61_U91 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_15_port, A2 => 
                           dp_ex_stage_alu_r61_n19, ZN => 
                           dp_ex_stage_alu_r61_n92);
   dp_ex_stage_alu_r61_U90 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_22_port, A2 => 
                           dp_ex_stage_alu_r61_n24, ZN => 
                           dp_ex_stage_alu_r61_n42);
   dp_ex_stage_alu_r61_U89 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_2_port, A2 => 
                           dp_ex_stage_alu_r61_n76, ZN => 
                           dp_ex_stage_alu_r61_n184);
   dp_ex_stage_alu_r61_U88 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n74, 
                           A2 => dp_ex_stage_alu_r61_n7, ZN => 
                           dp_ex_stage_alu_r61_n183);
   dp_ex_stage_alu_r61_U87 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n187,
                           A2 => dp_ex_stage_alu_r61_n74, ZN => 
                           dp_ex_stage_alu_r61_n185);
   dp_ex_stage_alu_r61_U86 : OAI211_X1 port map( C1 => dp_ex_stage_alu_r61_n183
                           , C2 => dp_ex_stage_alu_r61_n184, A => 
                           dp_ex_stage_alu_r61_n185, B => 
                           dp_ex_stage_alu_r61_n186, ZN => 
                           dp_ex_stage_alu_r61_n182);
   dp_ex_stage_alu_r61_U85 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n22, A2 
                           => dp_ex_stage_alu_r61_n197, ZN => 
                           dp_ex_stage_alu_r61_n74);
   dp_ex_stage_alu_r61_U84 : INV_X1 port map( A => dp_ex_stage_muxB_out_13_port
                           , ZN => dp_ex_stage_alu_r61_n180);
   dp_ex_stage_alu_r61_U83 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n180,
                           A2 => dp_ex_stage_muxA_out_13_port, ZN => 
                           dp_ex_stage_alu_r61_n161);
   dp_ex_stage_alu_r61_U82 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_16_port, A2 => 
                           dp_ex_stage_alu_r61_n20, ZN => 
                           dp_ex_stage_alu_r61_n93);
   dp_ex_stage_alu_r61_U81 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_10_port, A2 => 
                           dp_ex_stage_alu_r61_n14, ZN => 
                           dp_ex_stage_alu_r61_n79);
   dp_ex_stage_alu_r61_U80 : XNOR2_X1 port map( A => 
                           dp_ex_stage_muxB_out_31_port, B => 
                           dp_ex_stage_alu_r61_n31, ZN => 
                           dp_ex_stage_alu_r61_n99);
   dp_ex_stage_alu_r61_U79 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_17_port, A2 => 
                           dp_ex_stage_alu_r61_n21, ZN => 
                           dp_ex_stage_alu_r61_n45);
   dp_ex_stage_alu_r61_U78 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_12_port, A2 => 
                           dp_ex_stage_alu_r61_n16, ZN => 
                           dp_ex_stage_alu_r61_n87);
   dp_ex_stage_alu_r61_U77 : INV_X1 port map( A => dp_ex_stage_muxB_out_23_port
                           , ZN => dp_ex_stage_alu_r61_n133);
   dp_ex_stage_alu_r61_U76 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_23_port, A2 => 
                           dp_ex_stage_alu_r61_n133, ZN => 
                           dp_ex_stage_alu_r61_n132);
   dp_ex_stage_alu_r61_U75 : INV_X1 port map( A => dp_ex_stage_muxB_out_12_port
                           , ZN => dp_ex_stage_alu_r61_n172);
   dp_ex_stage_alu_r61_U74 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_12_port, A2 => 
                           dp_ex_stage_alu_r61_n172, ZN => 
                           dp_ex_stage_alu_r61_n162);
   dp_ex_stage_alu_r61_U73 : INV_X1 port map( A => dp_ex_stage_muxA_out_19_port
                           , ZN => dp_ex_stage_alu_r61_n214);
   dp_ex_stage_alu_r61_U72 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_19_port, A2 => 
                           dp_ex_stage_alu_r61_n214, ZN => 
                           dp_ex_stage_alu_r61_n43);
   dp_ex_stage_alu_r61_U71 : INV_X1 port map( A => dp_ex_stage_muxB_out_18_port
                           , ZN => dp_ex_stage_alu_r61_n217);
   dp_ex_stage_alu_r61_U70 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_18_port, A2 => 
                           dp_ex_stage_alu_r61_n217, ZN => 
                           dp_ex_stage_alu_r61_n147);
   dp_ex_stage_alu_r61_U69 : INV_X1 port map( A => dp_ex_stage_muxB_out_24_port
                           , ZN => dp_ex_stage_alu_r61_n130);
   dp_ex_stage_alu_r61_U68 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_24_port, A2 => 
                           dp_ex_stage_alu_r61_n130, ZN => 
                           dp_ex_stage_alu_r61_n118);
   dp_ex_stage_alu_r61_U67 : INV_X1 port map( A => dp_ex_stage_muxB_out_25_port
                           , ZN => dp_ex_stage_alu_r61_n138);
   dp_ex_stage_alu_r61_U66 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_25_port, A2 => 
                           dp_ex_stage_alu_r61_n138, ZN => 
                           dp_ex_stage_alu_r61_n117);
   dp_ex_stage_alu_r61_U65 : INV_X1 port map( A => dp_ex_stage_muxB_out_11_port
                           , ZN => dp_ex_stage_alu_r61_n175);
   dp_ex_stage_alu_r61_U64 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_11_port, A2 => 
                           dp_ex_stage_alu_r61_n175, ZN => 
                           dp_ex_stage_alu_r61_n174);
   dp_ex_stage_alu_r61_U63 : INV_X1 port map( A => dp_ex_stage_muxA_out_29_port
                           , ZN => dp_ex_stage_alu_r61_n101);
   dp_ex_stage_alu_r61_U62 : INV_X1 port map( A => dp_ex_stage_muxA_out_30_port
                           , ZN => dp_ex_stage_alu_r61_n62);
   dp_ex_stage_alu_r61_U61 : INV_X1 port map( A => dp_ex_stage_muxB_out_19_port
                           , ZN => dp_ex_stage_alu_r61_n220);
   dp_ex_stage_alu_r61_U60 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_19_port, A2 => 
                           dp_ex_stage_alu_r61_n220, ZN => 
                           dp_ex_stage_alu_r61_n155);
   dp_ex_stage_alu_r61_U59 : INV_X1 port map( A => dp_ex_stage_muxB_out_20_port
                           , ZN => dp_ex_stage_alu_r61_n135);
   dp_ex_stage_alu_r61_U58 : NAND4_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_20_port, A2 => 
                           dp_ex_stage_alu_r61_n51, A3 => 
                           dp_ex_stage_alu_r61_n42, A4 => 
                           dp_ex_stage_alu_r61_n135, ZN => 
                           dp_ex_stage_alu_r61_n126);
   dp_ex_stage_alu_r61_U57 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r61_n2, 
                           B2 => dp_ex_stage_alu_r61_n164, A => 
                           dp_ex_stage_alu_r61_n165, ZN => 
                           dp_ex_stage_alu_r61_n156);
   dp_ex_stage_alu_r61_U56 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n159, 
                           A2 => dp_ex_stage_alu_r61_n160, ZN => 
                           dp_ex_stage_alu_r61_n158);
   dp_ex_stage_alu_r61_U55 : AND3_X1 port map( A1 => dp_ex_stage_alu_r61_n156, 
                           A2 => dp_ex_stage_alu_r61_n157, A3 => 
                           dp_ex_stage_alu_r61_n158, ZN => 
                           dp_ex_stage_alu_r61_n140);
   dp_ex_stage_alu_r61_U54 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n34, 
                           A2 => dp_ex_stage_alu_r61_n35, ZN => 
                           dp_ex_stage_alu_r61_n33);
   dp_ex_stage_alu_r61_U53 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n3, 
                           A2 => dp_ex_stage_alu_r61_n33, ZN => 
                           dp_ex_stage_alu_N18_port);
   dp_ex_stage_alu_r61_U52 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n56, 
                           A2 => dp_ex_stage_alu_r61_n57, ZN => 
                           dp_ex_stage_alu_r61_n52);
   dp_ex_stage_alu_r61_U51 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n44, 
                           A2 => dp_ex_stage_alu_r61_n45, ZN => 
                           dp_ex_stage_alu_r61_n40);
   dp_ex_stage_alu_r61_U50 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n54, 
                           A2 => dp_ex_stage_alu_r61_n55, ZN => 
                           dp_ex_stage_alu_r61_n53);
   dp_ex_stage_alu_r61_U49 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n48, 
                           A2 => dp_ex_stage_alu_r61_n49, ZN => 
                           dp_ex_stage_alu_r61_n47);
   dp_ex_stage_alu_r61_U48 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n81, 
                           A2 => dp_ex_stage_alu_r61_n80, ZN => 
                           dp_ex_stage_alu_r61_n5);
   dp_ex_stage_alu_r61_U47 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n5, A2
                           => dp_ex_stage_alu_r61_n79, ZN => 
                           dp_ex_stage_alu_r61_n203);
   dp_ex_stage_alu_r61_U46 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n85, 
                           A2 => dp_ex_stage_alu_r61_n94, ZN => 
                           dp_ex_stage_alu_r61_n159);
   dp_ex_stage_alu_r61_U45 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n50, 
                           A2 => dp_ex_stage_alu_r61_n51, ZN => 
                           dp_ex_stage_alu_r61_n46);
   dp_ex_stage_alu_r61_U44 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n42, 
                           A2 => dp_ex_stage_alu_r61_n43, ZN => 
                           dp_ex_stage_alu_r61_n41);
   dp_ex_stage_alu_r61_U43 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n73, 
                           A2 => dp_ex_stage_alu_r61_n74, ZN => 
                           dp_ex_stage_alu_r61_n72);
   dp_ex_stage_alu_r61_U42 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n75, 
                           A2 => dp_ex_stage_alu_r61_n76, ZN => 
                           dp_ex_stage_alu_r61_n71);
   dp_ex_stage_alu_r61_U41 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n71, 
                           A2 => dp_ex_stage_alu_r61_n72, ZN => 
                           dp_ex_stage_alu_r61_n70);
   dp_ex_stage_alu_r61_U40 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n93, 
                           A2 => dp_ex_stage_alu_r61_n94, ZN => 
                           dp_ex_stage_alu_r61_n89);
   dp_ex_stage_alu_r61_U39 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n91, 
                           A2 => dp_ex_stage_alu_r61_n92, ZN => 
                           dp_ex_stage_alu_r61_n90);
   dp_ex_stage_alu_r61_U38 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n89, 
                           A2 => dp_ex_stage_alu_r61_n90, ZN => 
                           dp_ex_stage_alu_r61_n67);
   dp_ex_stage_alu_r61_U37 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n87, 
                           A2 => dp_ex_stage_alu_r61_n88, ZN => 
                           dp_ex_stage_alu_r61_n83);
   dp_ex_stage_alu_r61_U36 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n85, 
                           A2 => dp_ex_stage_alu_r61_n86, ZN => 
                           dp_ex_stage_alu_r61_n84);
   dp_ex_stage_alu_r61_U35 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n83, 
                           A2 => dp_ex_stage_alu_r61_n84, ZN => 
                           dp_ex_stage_alu_r61_n68);
   dp_ex_stage_alu_r61_U34 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n57, 
                           A2 => dp_ex_stage_alu_r61_n48, ZN => 
                           dp_ex_stage_alu_r61_n120);
   dp_ex_stage_alu_r61_U33 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n81, 
                           A2 => dp_ex_stage_alu_r61_n82, ZN => 
                           dp_ex_stage_alu_r61_n77);
   dp_ex_stage_alu_r61_U32 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n79, 
                           A2 => dp_ex_stage_alu_r61_n80, ZN => 
                           dp_ex_stage_alu_r61_n78);
   dp_ex_stage_alu_r61_U31 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n77, 
                           A2 => dp_ex_stage_alu_r61_n78, ZN => 
                           dp_ex_stage_alu_r61_n69);
   dp_ex_stage_alu_r61_U30 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n44, 
                           A2 => dp_ex_stage_alu_r61_n43, ZN => 
                           dp_ex_stage_alu_r61_n4);
   dp_ex_stage_alu_r61_U29 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n4, A2
                           => dp_ex_stage_alu_r61_n42, ZN => 
                           dp_ex_stage_alu_r61_n213);
   dp_ex_stage_alu_r61_U28 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_22_port, A2 => 
                           dp_ex_stage_alu_r61_n134, ZN => 
                           dp_ex_stage_alu_r61_n131);
   dp_ex_stage_alu_r61_U27 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n131,
                           A2 => dp_ex_stage_alu_r61_n132, ZN => 
                           dp_ex_stage_alu_r61_n128);
   dp_ex_stage_alu_r61_U26 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n128, 
                           A2 => dp_ex_stage_alu_r61_n129, ZN => 
                           dp_ex_stage_alu_r61_n127);
   dp_ex_stage_alu_r61_U25 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n117,
                           A2 => dp_ex_stage_alu_r61_n118, ZN => 
                           dp_ex_stage_alu_r61_n116);
   dp_ex_stage_alu_r61_U24 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n49, 
                           A2 => dp_ex_stage_alu_r61_n116, ZN => 
                           dp_ex_stage_alu_r61_n115);
   dp_ex_stage_alu_r61_U23 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n114, 
                           A2 => dp_ex_stage_alu_r61_n115, ZN => 
                           dp_ex_stage_alu_r61_n108);
   dp_ex_stage_alu_r61_U22 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n55, 
                           A2 => dp_ex_stage_alu_r61_n56, ZN => 
                           dp_ex_stage_alu_r61_n103);
   dp_ex_stage_alu_r61_U21 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n105, 
                           A2 => dp_ex_stage_alu_r61_n106, ZN => 
                           dp_ex_stage_alu_r61_n104);
   dp_ex_stage_alu_r61_U20 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r61_n102,
                           B2 => dp_ex_stage_alu_r61_n103, A => 
                           dp_ex_stage_alu_r61_n104, ZN => 
                           dp_ex_stage_alu_r61_n97);
   dp_ex_stage_alu_r61_U19 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n63, 
                           A2 => dp_ex_stage_alu_r61_n64, ZN => 
                           dp_ex_stage_alu_r61_n58);
   dp_ex_stage_alu_r61_U18 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n58, 
                           A2 => dp_ex_stage_alu_r61_n59, ZN => 
                           dp_ex_stage_alu_r61_n36);
   dp_ex_stage_alu_r61_U17 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r61_n186,
                           B2 => dp_ex_stage_alu_r61_n207, A => 
                           dp_ex_stage_alu_r61_n208, ZN => 
                           dp_ex_stage_alu_r61_n201);
   dp_ex_stage_alu_r61_U16 : OAI211_X1 port map( C1 => dp_ex_stage_alu_r61_n198
                           , C2 => dp_ex_stage_alu_r61_n199, A => 
                           dp_ex_stage_alu_r61_n200, B => 
                           dp_ex_stage_alu_r61_n73, ZN => 
                           dp_ex_stage_alu_r61_n188);
   dp_ex_stage_alu_r61_U15 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n191, 
                           A2 => dp_ex_stage_alu_r61_n192, ZN => 
                           dp_ex_stage_alu_r61_n190);
   dp_ex_stage_alu_r61_U14 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r61_n76, 
                           A2 => dp_ex_stage_alu_r61_n74, ZN => 
                           dp_ex_stage_alu_r61_n189);
   dp_ex_stage_alu_r61_U13 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r61_n188,
                           B2 => dp_ex_stage_alu_r61_n189, A => 
                           dp_ex_stage_alu_r61_n190, ZN => 
                           dp_ex_stage_alu_r61_n181);
   dp_ex_stage_alu_r61_U12 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r61_n155,
                           B2 => dp_ex_stage_alu_r61_n218, A => 
                           dp_ex_stage_alu_r61_n219, ZN => 
                           dp_ex_stage_alu_r61_n211);
   dp_ex_stage_alu_r61_U11 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n181, 
                           A2 => dp_ex_stage_alu_r61_n182, ZN => 
                           dp_ex_stage_alu_r61_n167);
   dp_ex_stage_alu_r61_U10 : AND3_X1 port map( A1 => dp_ex_stage_alu_r61_n169, 
                           A2 => dp_ex_stage_alu_r61_n170, A3 => 
                           dp_ex_stage_alu_r61_n171, ZN => 
                           dp_ex_stage_alu_r61_n168);
   dp_ex_stage_alu_r61_U9 : AND3_X1 port map( A1 => dp_ex_stage_alu_r61_n125, 
                           A2 => dp_ex_stage_alu_r61_n126, A3 => 
                           dp_ex_stage_alu_r61_n127, ZN => 
                           dp_ex_stage_alu_r61_n124);
   dp_ex_stage_alu_r61_U8 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n52, A2
                           => dp_ex_stage_alu_r61_n53, ZN => 
                           dp_ex_stage_alu_r61_n37);
   dp_ex_stage_alu_r61_U7 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n46, A2
                           => dp_ex_stage_alu_r61_n47, ZN => 
                           dp_ex_stage_alu_r61_n38);
   dp_ex_stage_alu_r61_U6 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r61_n40, A2
                           => dp_ex_stage_alu_r61_n41, ZN => 
                           dp_ex_stage_alu_r61_n39);
   dp_ex_stage_alu_r61_U5 : NAND4_X1 port map( A1 => dp_ex_stage_alu_r61_n36, 
                           A2 => dp_ex_stage_alu_r61_n37, A3 => 
                           dp_ex_stage_alu_r61_n38, A4 => 
                           dp_ex_stage_alu_r61_n39, ZN => 
                           dp_ex_stage_alu_r61_n35);
   dp_ex_stage_alu_r61_U4 : BUF_X1 port map( A => dp_ex_stage_alu_r61_n161, Z 
                           => dp_ex_stage_alu_r61_n2);
   dp_ex_stage_alu_r61_U3 : INV_X1 port map( A => dp_ex_stage_alu_r61_n3, ZN =>
                           dp_ex_stage_alu_N21_port);
   dp_ex_stage_alu_r61_U2 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n222, 
                           A2 => dp_ex_stage_alu_r61_n99, ZN => 
                           dp_ex_stage_alu_r61_n1);
   dp_ex_stage_alu_r61_U1 : AND2_X1 port map( A1 => dp_ex_stage_alu_r61_n95, A2
                           => dp_ex_stage_alu_r61_n96, ZN => 
                           dp_ex_stage_alu_r61_n3);
   dp_ex_stage_alu_r60_U318 : INV_X1 port map( A => dp_ex_stage_alu_r60_n4, ZN 
                           => dp_ex_stage_alu_r60_n306);
   dp_ex_stage_alu_r60_U317 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n306,
                           A2 => dp_ex_stage_alu_r60_n20, ZN => 
                           dp_ex_stage_alu_r60_n305);
   dp_ex_stage_alu_r60_U316 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r60_n304
                           , A2 => dp_ex_stage_alu_r60_n4, A3 => 
                           dp_ex_stage_alu_r60_n25, ZN => 
                           dp_ex_stage_alu_r60_n301);
   dp_ex_stage_alu_r60_U315 : INV_X1 port map( A => dp_ex_stage_alu_r60_n121, 
                           ZN => dp_ex_stage_alu_r60_n183);
   dp_ex_stage_alu_r60_U314 : INV_X1 port map( A => dp_ex_stage_alu_r60_n122, 
                           ZN => dp_ex_stage_alu_r60_n303);
   dp_ex_stage_alu_r60_U313 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n183,
                           A2 => dp_ex_stage_alu_r60_n303, ZN => 
                           dp_ex_stage_alu_r60_n302);
   dp_ex_stage_alu_r60_U312 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n19,
                           A2 => dp_ex_stage_alu_r60_n162, ZN => 
                           dp_ex_stage_alu_r60_n296);
   dp_ex_stage_alu_r60_U311 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r60_n285
                           , A2 => dp_ex_stage_alu_r60_n158, A3 => 
                           dp_ex_stage_alu_r60_n271, ZN => 
                           dp_ex_stage_alu_r60_n284);
   dp_ex_stage_alu_r60_U310 : INV_X1 port map( A => dp_ex_stage_alu_r60_n151, 
                           ZN => dp_ex_stage_alu_r60_n278);
   dp_ex_stage_alu_r60_U309 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n13, 
                           A2 => dp_ex_stage_alu_r60_n278, ZN => 
                           dp_ex_stage_alu_r60_n277);
   dp_ex_stage_alu_r60_U308 : INV_X1 port map( A => dp_ex_stage_alu_r60_n271, 
                           ZN => dp_ex_stage_alu_r60_n272);
   dp_ex_stage_alu_r60_U307 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n272,
                           A2 => dp_ex_stage_alu_r60_n14, ZN => 
                           dp_ex_stage_alu_r60_n270);
   dp_ex_stage_alu_r60_U306 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r60_n262
                           , A2 => dp_ex_stage_alu_r60_n135, A3 => 
                           dp_ex_stage_alu_r60_n263, ZN => 
                           dp_ex_stage_alu_r60_n261);
   dp_ex_stage_alu_r60_U305 : INV_X1 port map( A => dp_ex_stage_alu_r60_n252, 
                           ZN => dp_ex_stage_alu_r60_n251);
   dp_ex_stage_alu_r60_U304 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n251
                           , A2 => dp_ex_stage_alu_r60_n121, ZN => 
                           dp_ex_stage_alu_r60_n249);
   dp_ex_stage_alu_r60_U303 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r60_n245
                           , A2 => dp_ex_stage_alu_r60_n109, A3 => 
                           dp_ex_stage_alu_r60_n232, ZN => 
                           dp_ex_stage_alu_r60_n244);
   dp_ex_stage_alu_r60_U302 : INV_X1 port map( A => dp_ex_stage_alu_r60_n99, ZN
                           => dp_ex_stage_alu_r60_n93);
   dp_ex_stage_alu_r60_U301 : INV_X1 port map( A => dp_ex_stage_alu_r60_n226, 
                           ZN => dp_ex_stage_alu_r60_n225);
   dp_ex_stage_alu_r60_U300 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n225
                           , A2 => dp_ex_stage_alu_r60_n99, ZN => 
                           dp_ex_stage_alu_r60_n218);
   dp_ex_stage_alu_r60_U299 : INV_X1 port map( A => dp_ex_stage_alu_r60_n80, ZN
                           => dp_ex_stage_alu_r60_n220);
   dp_ex_stage_alu_r60_U298 : INV_X1 port map( A => dp_ex_stage_alu_r60_n222, 
                           ZN => dp_ex_stage_alu_r60_n221);
   dp_ex_stage_alu_r60_U297 : OAI211_X1 port map( C1 => dp_ex_stage_alu_r60_n12
                           , C2 => dp_ex_stage_alu_r60_n218, A => 
                           dp_ex_stage_alu_r60_n10, B => 
                           dp_ex_stage_alu_r60_n219, ZN => 
                           dp_ex_stage_alu_r60_n217);
   dp_ex_stage_alu_r60_U296 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n21,
                           A2 => dp_ex_stage_alu_r60_n84, ZN => 
                           dp_ex_stage_alu_r60_n209);
   dp_ex_stage_alu_r60_U295 : INV_X1 port map( A => dp_ex_stage_alu_r60_n213, 
                           ZN => dp_ex_stage_alu_r60_n211);
   dp_ex_stage_alu_r60_U294 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n22,
                           A2 => dp_ex_stage_alu_r60_n73, ZN => 
                           dp_ex_stage_alu_r60_n196);
   dp_ex_stage_alu_r60_U293 : INV_X1 port map( A => dp_ex_stage_alu_r60_n201, 
                           ZN => dp_ex_stage_alu_r60_n198);
   dp_ex_stage_alu_r60_U292 : INV_X1 port map( A => dp_ex_stage_alu_r60_n60, ZN
                           => dp_ex_stage_alu_r60_n199);
   dp_ex_stage_alu_r60_U291 : INV_X1 port map( A => dp_ex_stage_alu_r60_n187, 
                           ZN => dp_ex_stage_alu_r60_n58);
   dp_ex_stage_alu_r60_U290 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n67,
                           A2 => dp_ex_stage_alu_r60_n61, ZN => 
                           dp_ex_stage_alu_r60_n193);
   dp_ex_stage_alu_r60_U289 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n191
                           , A2 => dp_ex_stage_alu_r60_n192, ZN => 
                           dp_ex_stage_alu_r60_n190);
   dp_ex_stage_alu_r60_U288 : INV_X1 port map( A => dp_ex_stage_alu_r60_n123, 
                           ZN => dp_ex_stage_alu_r60_n182);
   dp_ex_stage_alu_r60_U287 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n182,
                           A2 => dp_ex_stage_alu_r60_n183, ZN => 
                           dp_ex_stage_alu_r60_n180);
   dp_ex_stage_alu_r60_U286 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r60_n121
                           , A2 => dp_ex_stage_alu_r60_n123, A3 => 
                           dp_ex_stage_alu_r60_n20, ZN => 
                           dp_ex_stage_alu_r60_n177);
   dp_ex_stage_alu_r60_U285 : NAND4_X1 port map( A1 => dp_ex_stage_alu_r60_n174
                           , A2 => dp_ex_stage_alu_r60_n175, A3 => 
                           dp_ex_stage_alu_r60_n176, A4 => 
                           dp_ex_stage_alu_r60_n177, ZN => 
                           dp_ex_stage_alu_r60_n100);
   dp_ex_stage_alu_r60_U284 : INV_X1 port map( A => dp_ex_stage_alu_r60_n155, 
                           ZN => dp_ex_stage_alu_r60_n169);
   dp_ex_stage_alu_r60_U283 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n169
                           , A2 => dp_ex_stage_alu_r60_n170, ZN => 
                           dp_ex_stage_alu_r60_n145);
   dp_ex_stage_alu_r60_U282 : INV_X1 port map( A => dp_ex_stage_alu_r60_n158, 
                           ZN => dp_ex_stage_alu_r60_n156);
   dp_ex_stage_alu_r60_U281 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r60_n143
                           , A2 => dp_ex_stage_alu_r60_n11, A3 => 
                           dp_ex_stage_alu_r60_n14, ZN => 
                           dp_ex_stage_alu_r60_n142);
   dp_ex_stage_alu_r60_U280 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n141
                           , A2 => dp_ex_stage_alu_r60_n142, ZN => 
                           dp_ex_stage_alu_r60_n130);
   dp_ex_stage_alu_r60_U279 : INV_X1 port map( A => dp_ex_stage_alu_r60_n11, ZN
                           => dp_ex_stage_alu_r60_n139);
   dp_ex_stage_alu_r60_U278 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n139,
                           A2 => dp_ex_stage_alu_r60_n13, ZN => 
                           dp_ex_stage_alu_r60_n137);
   dp_ex_stage_alu_r60_U277 : INV_X1 port map( A => dp_ex_stage_alu_r60_n136, 
                           ZN => dp_ex_stage_alu_r60_n134);
   dp_ex_stage_alu_r60_U276 : INV_X1 port map( A => dp_ex_stage_alu_r60_n135, 
                           ZN => dp_ex_stage_alu_r60_n128);
   dp_ex_stage_alu_r60_U275 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n134,
                           A2 => dp_ex_stage_alu_r60_n128, ZN => 
                           dp_ex_stage_alu_r60_n133);
   dp_ex_stage_alu_r60_U274 : INV_X1 port map( A => dp_ex_stage_alu_r60_n127, 
                           ZN => dp_ex_stage_alu_r60_n125);
   dp_ex_stage_alu_r60_U273 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n126
                           , A2 => dp_ex_stage_alu_r60_n125, ZN => 
                           dp_ex_stage_alu_r60_n116);
   dp_ex_stage_alu_r60_U272 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n125
                           , A2 => dp_ex_stage_alu_r60_n25, ZN => 
                           dp_ex_stage_alu_r60_n117);
   dp_ex_stage_alu_r60_U271 : NAND3_X1 port map( A1 => dp_ex_stage_alu_r60_n116
                           , A2 => dp_ex_stage_alu_r60_n117, A3 => 
                           dp_ex_stage_alu_r60_n118, ZN => 
                           dp_ex_stage_alu_r60_n115);
   dp_ex_stage_alu_r60_U270 : INV_X1 port map( A => dp_ex_stage_alu_r60_n110, 
                           ZN => dp_ex_stage_alu_r60_n108);
   dp_ex_stage_alu_r60_U269 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n108
                           , A2 => dp_ex_stage_alu_r60_n109, ZN => 
                           dp_ex_stage_alu_r60_n106);
   dp_ex_stage_alu_r60_U268 : INV_X1 port map( A => dp_ex_stage_alu_r60_n12, ZN
                           => dp_ex_stage_alu_r60_n97);
   dp_ex_stage_alu_r60_U267 : INV_X1 port map( A => dp_ex_stage_alu_r60_n94, ZN
                           => dp_ex_stage_alu_r60_n92);
   dp_ex_stage_alu_r60_U266 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n92, 
                           A2 => dp_ex_stage_alu_r60_n93, ZN => 
                           dp_ex_stage_alu_r60_n90);
   dp_ex_stage_alu_r60_U265 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n21,
                           A2 => dp_ex_stage_alu_r60_n80, ZN => 
                           dp_ex_stage_alu_r60_n76);
   dp_ex_stage_alu_r60_U264 : INV_X1 port map( A => dp_ex_stage_alu_r60_n79, ZN
                           => dp_ex_stage_alu_r60_n78);
   dp_ex_stage_alu_r60_U263 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n22,
                           A2 => dp_ex_stage_alu_r60_n69, ZN => 
                           dp_ex_stage_alu_r60_n63);
   dp_ex_stage_alu_r60_U262 : INV_X1 port map( A => dp_ex_stage_alu_r60_n68, ZN
                           => dp_ex_stage_alu_r60_n65);
   dp_ex_stage_alu_r60_U261 : INV_X1 port map( A => dp_ex_stage_alu_r60_n67, ZN
                           => dp_ex_stage_alu_r60_n66);
   dp_ex_stage_alu_r60_U260 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n60,
                           A2 => dp_ex_stage_alu_r60_n61, ZN => 
                           dp_ex_stage_alu_r60_n59);
   dp_ex_stage_alu_r60_U259 : INV_X1 port map( A => dp_ex_stage_alu_N22_port, 
                           ZN => dp_ex_stage_alu_N16_port);
   dp_ex_stage_alu_r60_U258 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_31_port, ZN => 
                           dp_ex_stage_alu_r60_n53);
   dp_ex_stage_alu_r60_U257 : INV_X1 port map( A => dp_ex_stage_alu_n247, ZN =>
                           dp_ex_stage_alu_r60_n52);
   dp_ex_stage_alu_r60_U256 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_27_port, ZN => 
                           dp_ex_stage_alu_r60_n51);
   dp_ex_stage_alu_r60_U255 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_26_port, ZN => 
                           dp_ex_stage_alu_r60_n50);
   dp_ex_stage_alu_r60_U254 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_25_port, ZN => 
                           dp_ex_stage_alu_r60_n49);
   dp_ex_stage_alu_r60_U253 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_24_port, ZN => 
                           dp_ex_stage_alu_r60_n48);
   dp_ex_stage_alu_r60_U252 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_23_port, ZN => 
                           dp_ex_stage_alu_r60_n47);
   dp_ex_stage_alu_r60_U251 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_22_port, ZN => 
                           dp_ex_stage_alu_r60_n46);
   dp_ex_stage_alu_r60_U250 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_21_port, ZN => 
                           dp_ex_stage_alu_r60_n45);
   dp_ex_stage_alu_r60_U249 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_18_port, ZN => 
                           dp_ex_stage_alu_r60_n44);
   dp_ex_stage_alu_r60_U248 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_17_port, ZN => 
                           dp_ex_stage_alu_r60_n43);
   dp_ex_stage_alu_r60_U247 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_16_port, ZN => 
                           dp_ex_stage_alu_r60_n42);
   dp_ex_stage_alu_r60_U246 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_15_port, ZN => 
                           dp_ex_stage_alu_r60_n41);
   dp_ex_stage_alu_r60_U245 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_14_port, ZN => 
                           dp_ex_stage_alu_r60_n40);
   dp_ex_stage_alu_r60_U244 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_13_port, ZN => 
                           dp_ex_stage_alu_r60_n39);
   dp_ex_stage_alu_r60_U243 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_12_port, ZN => 
                           dp_ex_stage_alu_r60_n38);
   dp_ex_stage_alu_r60_U242 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_11_port, ZN => 
                           dp_ex_stage_alu_r60_n37);
   dp_ex_stage_alu_r60_U241 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_10_port, ZN => 
                           dp_ex_stage_alu_r60_n36);
   dp_ex_stage_alu_r60_U240 : INV_X1 port map( A => dp_ex_stage_muxA_out_9_port
                           , ZN => dp_ex_stage_alu_r60_n35);
   dp_ex_stage_alu_r60_U239 : INV_X1 port map( A => dp_ex_stage_muxA_out_8_port
                           , ZN => dp_ex_stage_alu_r60_n34);
   dp_ex_stage_alu_r60_U238 : INV_X1 port map( A => dp_ex_stage_muxA_out_7_port
                           , ZN => dp_ex_stage_alu_r60_n33);
   dp_ex_stage_alu_r60_U237 : INV_X1 port map( A => dp_ex_stage_muxA_out_3_port
                           , ZN => dp_ex_stage_alu_r60_n32);
   dp_ex_stage_alu_r60_U236 : INV_X1 port map( A => dp_ex_stage_muxA_out_2_port
                           , ZN => dp_ex_stage_alu_r60_n31);
   dp_ex_stage_alu_r60_U235 : INV_X1 port map( A => dp_ex_stage_muxB_out_4_port
                           , ZN => dp_ex_stage_alu_r60_n30);
   dp_ex_stage_alu_r60_U234 : INV_X1 port map( A => dp_ex_stage_alu_n77, ZN => 
                           dp_ex_stage_alu_r60_n29);
   dp_ex_stage_alu_r60_U233 : INV_X1 port map( A => dp_ex_stage_alu_n73, ZN => 
                           dp_ex_stage_alu_r60_n28);
   dp_ex_stage_alu_r60_U232 : INV_X1 port map( A => dp_ex_stage_alu_n46, ZN => 
                           dp_ex_stage_alu_r60_n27);
   dp_ex_stage_alu_r60_U231 : INV_X1 port map( A => dp_ex_stage_alu_n45, ZN => 
                           dp_ex_stage_alu_r60_n26);
   dp_ex_stage_alu_r60_U230 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n32,
                           A2 => dp_ex_stage_alu_n77, ZN => 
                           dp_ex_stage_alu_r60_n162);
   dp_ex_stage_alu_r60_U229 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n266,
                           A2 => dp_ex_stage_alu_r60_n267, ZN => 
                           dp_ex_stage_alu_r60_n254);
   dp_ex_stage_alu_r60_U228 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n256
                           , A2 => dp_ex_stage_alu_r60_n257, ZN => 
                           dp_ex_stage_alu_r60_n255);
   dp_ex_stage_alu_r60_U227 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r60_n253
                           , B2 => dp_ex_stage_alu_r60_n254, A => 
                           dp_ex_stage_alu_r60_n255, ZN => 
                           dp_ex_stage_alu_r60_n240);
   dp_ex_stage_alu_r60_U226 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n240
                           , B2 => dp_ex_stage_alu_r60_n239, A => 
                           dp_ex_stage_alu_r60_n241, ZN => 
                           dp_ex_stage_alu_r60_n215);
   dp_ex_stage_alu_r60_U225 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r60_n215
                           , B2 => dp_ex_stage_alu_r60_n216, A => 
                           dp_ex_stage_alu_r60_n217, ZN => 
                           dp_ex_stage_alu_r60_n208);
   dp_ex_stage_alu_r60_U224 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n46, A2 
                           => dp_ex_stage_alu_r60_n291, ZN => 
                           dp_ex_stage_alu_r60_n290);
   dp_ex_stage_alu_r60_U223 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n208
                           , B2 => dp_ex_stage_alu_r60_n209, A => 
                           dp_ex_stage_alu_r60_n210, ZN => 
                           dp_ex_stage_alu_r60_n204);
   dp_ex_stage_alu_r60_U222 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n195
                           , B2 => dp_ex_stage_alu_r60_n196, A => 
                           dp_ex_stage_alu_r60_n197, ZN => 
                           dp_ex_stage_alu_r60_n191);
   dp_ex_stage_alu_r60_U221 : INV_X1 port map( A => dp_ex_stage_muxA_out_4_port
                           , ZN => dp_ex_stage_alu_r60_n298);
   dp_ex_stage_alu_r60_U220 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_4_port, A2 => 
                           dp_ex_stage_alu_r60_n30, ZN => 
                           dp_ex_stage_alu_r60_n285);
   dp_ex_stage_alu_r60_U219 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n7, 
                           A2 => dp_ex_stage_alu_r60_n31, ZN => 
                           dp_ex_stage_alu_r60_n163);
   dp_ex_stage_alu_r60_U218 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_6_port, A2 => 
                           dp_ex_stage_alu_r60_n286, ZN => 
                           dp_ex_stage_alu_r60_n271);
   dp_ex_stage_alu_r60_U217 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_10_port, A2 => 
                           dp_ex_stage_alu_r60_n274, ZN => 
                           dp_ex_stage_alu_r60_n262);
   dp_ex_stage_alu_r60_U216 : NOR3_X1 port map( A1 => dp_ex_stage_alu_r60_n144,
                           A2 => dp_ex_stage_alu_r60_n13, A3 => 
                           dp_ex_stage_alu_r60_n259, ZN => 
                           dp_ex_stage_alu_r60_n258);
   dp_ex_stage_alu_r60_U215 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n258,
                           A2 => dp_ex_stage_alu_r60_n20, ZN => 
                           dp_ex_stage_alu_r60_n257);
   dp_ex_stage_alu_r60_U214 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r60_n204
                           , B2 => dp_ex_stage_alu_r60_n203, A => 
                           dp_ex_stage_alu_r60_n205, ZN => 
                           dp_ex_stage_alu_r60_n195);
   dp_ex_stage_alu_r60_U213 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_31_port, ZN => 
                           dp_ex_stage_alu_r60_n315);
   dp_ex_stage_alu_r60_U212 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_31_port, A2 => 
                           dp_ex_stage_alu_r60_n53, ZN => 
                           dp_ex_stage_alu_r60_n185);
   dp_ex_stage_alu_r60_U211 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n56,
                           A2 => dp_ex_stage_alu_r60_n57, ZN => 
                           dp_ex_stage_alu_r60_n55);
   dp_ex_stage_alu_r60_U210 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n185,
                           A2 => dp_ex_stage_alu_r60_n3, ZN => 
                           dp_ex_stage_alu_r60_n54);
   dp_ex_stage_alu_r60_U209 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n54,
                           A2 => dp_ex_stage_alu_r60_n55, ZN => 
                           dp_ex_stage_alu_N22_port);
   dp_ex_stage_alu_r60_U208 : INV_X1 port map( A => dp_ex_stage_muxA_out_1_port
                           , ZN => dp_ex_stage_alu_r60_n291);
   dp_ex_stage_alu_r60_U207 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_10_port, ZN => 
                           dp_ex_stage_alu_r60_n274);
   dp_ex_stage_alu_r60_U206 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_30_port, ZN => 
                           dp_ex_stage_alu_r60_n314);
   dp_ex_stage_alu_r60_U205 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_30_port, A2 => 
                           dp_ex_stage_alu_r60_n314, ZN => 
                           dp_ex_stage_alu_r60_n313);
   dp_ex_stage_alu_r60_U204 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_30_port, ZN => 
                           dp_ex_stage_alu_r60_n188);
   dp_ex_stage_alu_r60_U203 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_30_port, A2 => 
                           dp_ex_stage_alu_r60_n188, ZN => 
                           dp_ex_stage_alu_r60_n186);
   dp_ex_stage_alu_r60_U202 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_10_port, A2 => 
                           dp_ex_stage_alu_r60_n36, ZN => 
                           dp_ex_stage_alu_r60_n129);
   dp_ex_stage_alu_r60_U201 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n1, 
                           A2 => dp_ex_stage_alu_r60_n298, ZN => 
                           dp_ex_stage_alu_r60_n157);
   dp_ex_stage_alu_r60_U200 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n28,
                           A2 => dp_ex_stage_muxA_out_2_port, ZN => 
                           dp_ex_stage_alu_r60_n293);
   dp_ex_stage_alu_r60_U199 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_8_port, A2 => 
                           dp_ex_stage_alu_r60_n34, ZN => 
                           dp_ex_stage_alu_r60_n140);
   dp_ex_stage_alu_r60_U198 : AND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_11_port, A2 => 
                           dp_ex_stage_alu_r60_n37, ZN => 
                           dp_ex_stage_alu_r60_n25);
   dp_ex_stage_alu_r60_U197 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n15,
                           A2 => dp_ex_stage_alu_r60_n27, ZN => 
                           dp_ex_stage_alu_r60_n168);
   dp_ex_stage_alu_r60_U196 : INV_X1 port map( A => dp_ex_stage_muxB_out_9_port
                           , ZN => dp_ex_stage_alu_r60_n265);
   dp_ex_stage_alu_r60_U195 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_9_port, A2 => 
                           dp_ex_stage_alu_r60_n265, ZN => 
                           dp_ex_stage_alu_r60_n136);
   dp_ex_stage_alu_r60_U194 : INV_X1 port map( A => dp_ex_stage_muxB_out_8_port
                           , ZN => dp_ex_stage_alu_r60_n275);
   dp_ex_stage_alu_r60_U193 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_8_port, A2 => 
                           dp_ex_stage_alu_r60_n275, ZN => 
                           dp_ex_stage_alu_r60_n259);
   dp_ex_stage_alu_r60_U192 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n29,
                           A2 => dp_ex_stage_muxA_out_3_port, ZN => 
                           dp_ex_stage_alu_r60_n173);
   dp_ex_stage_alu_r60_U191 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_29_port, ZN => 
                           dp_ex_stage_alu_r60_n194);
   dp_ex_stage_alu_r60_U190 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_29_port, A2 => 
                           dp_ex_stage_alu_r60_n194, ZN => 
                           dp_ex_stage_alu_r60_n67);
   dp_ex_stage_alu_r60_U189 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_0_port, A2 => 
                           dp_ex_stage_alu_r60_n26, ZN => 
                           dp_ex_stage_alu_r60_n166);
   dp_ex_stage_alu_r60_U188 : INV_X1 port map( A => dp_ex_stage_muxB_out_5_port
                           , ZN => dp_ex_stage_alu_r60_n287);
   dp_ex_stage_alu_r60_U187 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_5_port, A2 => 
                           dp_ex_stage_alu_r60_n287, ZN => 
                           dp_ex_stage_alu_r60_n158);
   dp_ex_stage_alu_r60_U186 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_23_port, A2 => 
                           dp_ex_stage_alu_r60_n47, ZN => 
                           dp_ex_stage_alu_r60_n84);
   dp_ex_stage_alu_r60_U185 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n15, 
                           A2 => dp_ex_stage_alu_r60_n27, ZN => 
                           dp_ex_stage_alu_r60_n167);
   dp_ex_stage_alu_r60_U184 : INV_X1 port map( A => dp_ex_stage_muxB_out_7_port
                           , ZN => dp_ex_stage_alu_r60_n297);
   dp_ex_stage_alu_r60_U183 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_7_port, A2 => 
                           dp_ex_stage_alu_r60_n297, ZN => 
                           dp_ex_stage_alu_r60_n273);
   dp_ex_stage_alu_r60_U182 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_13_port, A2 => 
                           dp_ex_stage_alu_r60_n39, ZN => 
                           dp_ex_stage_alu_r60_n122);
   dp_ex_stage_alu_r60_U181 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_7_port, A2 => 
                           dp_ex_stage_alu_r60_n33, ZN => 
                           dp_ex_stage_alu_r60_n151);
   dp_ex_stage_alu_r60_U180 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_24_port, A2 => 
                           dp_ex_stage_alu_r60_n48, ZN => 
                           dp_ex_stage_alu_r60_n79);
   dp_ex_stage_alu_r60_U179 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_16_port, A2 => 
                           dp_ex_stage_alu_r60_n42, ZN => 
                           dp_ex_stage_alu_r60_n110);
   dp_ex_stage_alu_r60_U178 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_28_port, A2 => 
                           dp_ex_stage_alu_r60_n52, ZN => 
                           dp_ex_stage_alu_r60_n68);
   dp_ex_stage_alu_r60_U177 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_26_port, A2 => 
                           dp_ex_stage_alu_r60_n50, ZN => 
                           dp_ex_stage_alu_r60_n74);
   dp_ex_stage_alu_r60_U176 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_22_port, A2 => 
                           dp_ex_stage_alu_r60_n46, ZN => 
                           dp_ex_stage_alu_r60_n85);
   dp_ex_stage_alu_r60_U175 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_17_port, A2 => 
                           dp_ex_stage_alu_r60_n43, ZN => 
                           dp_ex_stage_alu_r60_n107);
   dp_ex_stage_alu_r60_U174 : INV_X1 port map( A => dp_ex_stage_muxA_out_5_port
                           , ZN => dp_ex_stage_alu_r60_n279);
   dp_ex_stage_alu_r60_U173 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_5_port, A2 => 
                           dp_ex_stage_alu_r60_n279, ZN => 
                           dp_ex_stage_alu_r60_n159);
   dp_ex_stage_alu_r60_U172 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_12_port, A2 => 
                           dp_ex_stage_alu_r60_n38, ZN => 
                           dp_ex_stage_alu_r60_n124);
   dp_ex_stage_alu_r60_U171 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n44,
                           A2 => dp_ex_stage_muxB_out_18_port, ZN => 
                           dp_ex_stage_alu_r60_n112);
   dp_ex_stage_alu_r60_U170 : AND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_25_port, A2 => 
                           dp_ex_stage_alu_r60_n49, ZN => 
                           dp_ex_stage_alu_r60_n24);
   dp_ex_stage_alu_r60_U169 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_13_port, ZN => 
                           dp_ex_stage_alu_r60_n307);
   dp_ex_stage_alu_r60_U168 : AND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_25_port, A2 => 
                           dp_ex_stage_alu_r60_n212, ZN => 
                           dp_ex_stage_alu_r60_n23);
   dp_ex_stage_alu_r60_U167 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_15_port, A2 => 
                           dp_ex_stage_alu_r60_n41, ZN => 
                           dp_ex_stage_alu_r60_n121);
   dp_ex_stage_alu_r60_U166 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_22_port, ZN => 
                           dp_ex_stage_alu_r60_n233);
   dp_ex_stage_alu_r60_U165 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_22_port, A2 => 
                           dp_ex_stage_alu_r60_n233, ZN => 
                           dp_ex_stage_alu_r60_n222);
   dp_ex_stage_alu_r60_U164 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_21_port, A2 => 
                           dp_ex_stage_alu_r60_n45, ZN => 
                           dp_ex_stage_alu_r60_n99);
   dp_ex_stage_alu_r60_U163 : INV_X1 port map( A => dp_ex_stage_muxA_out_0_port
                           , ZN => dp_ex_stage_alu_r60_n292);
   dp_ex_stage_alu_r60_U162 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_14_port, A2 => 
                           dp_ex_stage_alu_r60_n40, ZN => 
                           dp_ex_stage_alu_r60_n123);
   dp_ex_stage_alu_r60_U161 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_20_port, ZN => 
                           dp_ex_stage_alu_r60_n234);
   dp_ex_stage_alu_r60_U160 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_20_port, A2 => 
                           dp_ex_stage_alu_r60_n234, ZN => 
                           dp_ex_stage_alu_r60_n94);
   dp_ex_stage_alu_r60_U159 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_27_port, A2 => 
                           dp_ex_stage_alu_r60_n51, ZN => 
                           dp_ex_stage_alu_r60_n73);
   dp_ex_stage_alu_r60_U158 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_23_port, ZN => 
                           dp_ex_stage_alu_r60_n223);
   dp_ex_stage_alu_r60_U157 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_23_port, A2 => 
                           dp_ex_stage_alu_r60_n223, ZN => 
                           dp_ex_stage_alu_r60_n80);
   dp_ex_stage_alu_r60_U156 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_28_port, ZN => 
                           dp_ex_stage_alu_r60_n202);
   dp_ex_stage_alu_r60_U155 : NAND2_X1 port map( A1 => dp_ex_stage_alu_n247, A2
                           => dp_ex_stage_alu_r60_n202, ZN => 
                           dp_ex_stage_alu_r60_n201);
   dp_ex_stage_alu_r60_U154 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_27_port, ZN => 
                           dp_ex_stage_alu_r60_n207);
   dp_ex_stage_alu_r60_U153 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_27_port, A2 => 
                           dp_ex_stage_alu_r60_n207, ZN => 
                           dp_ex_stage_alu_r60_n69);
   dp_ex_stage_alu_r60_U152 : XNOR2_X1 port map( A => 
                           dp_ex_stage_muxA_out_31_port, B => 
                           dp_ex_stage_muxB_out_31_port, ZN => 
                           dp_ex_stage_alu_r60_n187);
   dp_ex_stage_alu_r60_U151 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_24_port, ZN => 
                           dp_ex_stage_alu_r60_n214);
   dp_ex_stage_alu_r60_U150 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_24_port, A2 => 
                           dp_ex_stage_alu_r60_n214, ZN => 
                           dp_ex_stage_alu_r60_n213);
   dp_ex_stage_alu_r60_U149 : INV_X1 port map( A => 
                           dp_ex_stage_muxA_out_19_port, ZN => 
                           dp_ex_stage_alu_r60_n238);
   dp_ex_stage_alu_r60_U148 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxB_out_19_port, A2 => 
                           dp_ex_stage_alu_r60_n238, ZN => 
                           dp_ex_stage_alu_r60_n111);
   dp_ex_stage_alu_r60_U147 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_17_port, ZN => 
                           dp_ex_stage_alu_r60_n247);
   dp_ex_stage_alu_r60_U146 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_17_port, A2 => 
                           dp_ex_stage_alu_r60_n247, ZN => 
                           dp_ex_stage_alu_r60_n109);
   dp_ex_stage_alu_r60_U145 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_26_port, ZN => 
                           dp_ex_stage_alu_r60_n311);
   dp_ex_stage_alu_r60_U144 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_26_port, A2 => 
                           dp_ex_stage_alu_r60_n311, ZN => 
                           dp_ex_stage_alu_r60_n206);
   dp_ex_stage_alu_r60_U143 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_21_port, ZN => 
                           dp_ex_stage_alu_r60_n224);
   dp_ex_stage_alu_r60_U142 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_21_port, A2 => 
                           dp_ex_stage_alu_r60_n224, ZN => 
                           dp_ex_stage_alu_r60_n89);
   dp_ex_stage_alu_r60_U141 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_15_port, ZN => 
                           dp_ex_stage_alu_r60_n248);
   dp_ex_stage_alu_r60_U140 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_15_port, A2 => 
                           dp_ex_stage_alu_r60_n248, ZN => 
                           dp_ex_stage_alu_r60_n179);
   dp_ex_stage_alu_r60_U139 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_11_port, ZN => 
                           dp_ex_stage_alu_r60_n264);
   dp_ex_stage_alu_r60_U138 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_11_port, A2 => 
                           dp_ex_stage_alu_r60_n264, ZN => 
                           dp_ex_stage_alu_r60_n135);
   dp_ex_stage_alu_r60_U137 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_16_port, ZN => 
                           dp_ex_stage_alu_r60_n309);
   dp_ex_stage_alu_r60_U136 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_16_port, A2 => 
                           dp_ex_stage_alu_r60_n309, ZN => 
                           dp_ex_stage_alu_r60_n245);
   dp_ex_stage_alu_r60_U135 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_14_port, ZN => 
                           dp_ex_stage_alu_r60_n310);
   dp_ex_stage_alu_r60_U134 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_14_port, A2 => 
                           dp_ex_stage_alu_r60_n310, ZN => 
                           dp_ex_stage_alu_r60_n252);
   dp_ex_stage_alu_r60_U133 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_12_port, ZN => 
                           dp_ex_stage_alu_r60_n308);
   dp_ex_stage_alu_r60_U132 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_12_port, A2 => 
                           dp_ex_stage_alu_r60_n308, ZN => 
                           dp_ex_stage_alu_r60_n263);
   dp_ex_stage_alu_r60_U131 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_29_port, ZN => 
                           dp_ex_stage_alu_r60_n200);
   dp_ex_stage_alu_r60_U130 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_29_port, A2 => 
                           dp_ex_stage_alu_r60_n200, ZN => 
                           dp_ex_stage_alu_r60_n60);
   dp_ex_stage_alu_r60_U129 : INV_X1 port map( A => dp_ex_stage_muxB_out_6_port
                           , ZN => dp_ex_stage_alu_r60_n286);
   dp_ex_stage_alu_r60_U128 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_20_port, ZN => 
                           dp_ex_stage_alu_r60_n235);
   dp_ex_stage_alu_r60_U127 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_20_port, A2 => 
                           dp_ex_stage_alu_r60_n235, ZN => 
                           dp_ex_stage_alu_r60_n226);
   dp_ex_stage_alu_r60_U126 : XNOR2_X1 port map( A => 
                           dp_ex_stage_muxA_out_30_port, B => 
                           dp_ex_stage_muxB_out_30_port, ZN => 
                           dp_ex_stage_alu_r60_n61);
   dp_ex_stage_alu_r60_U125 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_18_port, ZN => 
                           dp_ex_stage_alu_r60_n246);
   dp_ex_stage_alu_r60_U124 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_18_port, A2 => 
                           dp_ex_stage_alu_r60_n246, ZN => 
                           dp_ex_stage_alu_r60_n232);
   dp_ex_stage_alu_r60_U123 : INV_X1 port map( A => 
                           dp_ex_stage_muxB_out_19_port, ZN => 
                           dp_ex_stage_alu_r60_n250);
   dp_ex_stage_alu_r60_U122 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_19_port, A2 => 
                           dp_ex_stage_alu_r60_n250, ZN => 
                           dp_ex_stage_alu_r60_n95);
   dp_ex_stage_alu_r60_U121 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n220,
                           A2 => dp_ex_stage_alu_r60_n221, ZN => 
                           dp_ex_stage_alu_r60_n219);
   dp_ex_stage_alu_r60_U120 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n180
                           , A2 => dp_ex_stage_alu_r60_n181, ZN => 
                           dp_ex_stage_alu_r60_n174);
   dp_ex_stage_alu_r60_U119 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n137
                           , A2 => dp_ex_stage_alu_r60_n138, ZN => 
                           dp_ex_stage_alu_r60_n132);
   dp_ex_stage_alu_r60_U118 : NOR2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_31_port, A2 => 
                           dp_ex_stage_alu_r60_n315, ZN => 
                           dp_ex_stage_alu_r60_n312);
   dp_ex_stage_alu_r60_U117 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n312,
                           A2 => dp_ex_stage_alu_r60_n2, ZN => 
                           dp_ex_stage_alu_r60_n189);
   dp_ex_stage_alu_r60_U116 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n190
                           , A2 => dp_ex_stage_alu_r60_n189, ZN => 
                           dp_ex_stage_alu_N20_port);
   dp_ex_stage_alu_r60_U115 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n90,
                           A2 => dp_ex_stage_alu_r60_n91, ZN => 
                           dp_ex_stage_alu_r60_n88);
   dp_ex_stage_alu_r60_U114 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n260,
                           A2 => dp_ex_stage_alu_r60_n261, ZN => 
                           dp_ex_stage_alu_r60_n256);
   dp_ex_stage_alu_r60_U113 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n305
                           , A2 => dp_ex_stage_alu_r60_n127, ZN => 
                           dp_ex_stage_alu_r60_n300);
   dp_ex_stage_alu_r60_U112 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n143
                           , A2 => dp_ex_stage_alu_r60_n151, ZN => 
                           dp_ex_stage_alu_r60_n150);
   dp_ex_stage_alu_r60_U111 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n73,
                           A2 => dp_ex_stage_alu_r60_n74, ZN => 
                           dp_ex_stage_alu_r60_n72);
   dp_ex_stage_alu_r60_U110 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n84,
                           A2 => dp_ex_stage_alu_r60_n85, ZN => 
                           dp_ex_stage_alu_r60_n83);
   dp_ex_stage_alu_r60_U109 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n121
                           , A2 => dp_ex_stage_alu_r60_n122, ZN => 
                           dp_ex_stage_alu_r60_n120);
   dp_ex_stage_alu_r60_U108 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n232,
                           A2 => dp_ex_stage_alu_r60_n95, ZN => 
                           dp_ex_stage_alu_r60_n231);
   dp_ex_stage_alu_r60_U107 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n11,
                           A2 => dp_ex_stage_alu_r60_n152, ZN => 
                           dp_ex_stage_alu_r60_n149);
   dp_ex_stage_alu_r60_U106 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n123
                           , A2 => dp_ex_stage_alu_r60_n124, ZN => 
                           dp_ex_stage_alu_r60_n119);
   dp_ex_stage_alu_r60_U105 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n270
                           , A2 => dp_ex_stage_alu_r60_n155, ZN => 
                           dp_ex_stage_alu_r60_n269);
   dp_ex_stage_alu_r60_U104 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n69,
                           A2 => dp_ex_stage_alu_r60_n206, ZN => 
                           dp_ex_stage_alu_r60_n205);
   dp_ex_stage_alu_r60_U103 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n201,
                           A2 => dp_ex_stage_alu_r60_n68, ZN => 
                           dp_ex_stage_alu_r60_n22);
   dp_ex_stage_alu_r60_U102 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n213,
                           A2 => dp_ex_stage_alu_r60_n79, ZN => 
                           dp_ex_stage_alu_r60_n21);
   dp_ex_stage_alu_r60_U101 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n128,
                           A2 => dp_ex_stage_alu_r60_n129, ZN => 
                           dp_ex_stage_alu_r60_n126);
   dp_ex_stage_alu_r60_U100 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n24, 
                           A2 => dp_ex_stage_alu_r60_n184, ZN => 
                           dp_ex_stage_alu_r60_n203);
   dp_ex_stage_alu_r60_U99 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n95, 
                           A2 => dp_ex_stage_alu_r60_n232, ZN => 
                           dp_ex_stage_alu_r60_n236);
   dp_ex_stage_alu_r60_U98 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n229,
                           A2 => dp_ex_stage_alu_r60_n230, ZN => 
                           dp_ex_stage_alu_r60_n228);
   dp_ex_stage_alu_r60_U97 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n107,
                           B2 => dp_ex_stage_alu_r60_n236, A => 
                           dp_ex_stage_alu_r60_n237, ZN => 
                           dp_ex_stage_alu_r60_n227);
   dp_ex_stage_alu_r60_U96 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n227, 
                           A2 => dp_ex_stage_alu_r60_n228, ZN => 
                           dp_ex_stage_alu_r60_n216);
   dp_ex_stage_alu_r60_U95 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n58, 
                           A2 => dp_ex_stage_alu_r60_n193, ZN => 
                           dp_ex_stage_alu_r60_n192);
   dp_ex_stage_alu_r60_U94 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n158,
                           A2 => dp_ex_stage_alu_r60_n173, ZN => 
                           dp_ex_stage_alu_r60_n172);
   dp_ex_stage_alu_r60_U93 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n171, 
                           A2 => dp_ex_stage_alu_r60_n172, ZN => 
                           dp_ex_stage_alu_r60_n170);
   dp_ex_stage_alu_r60_U92 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n259,
                           A2 => dp_ex_stage_alu_r60_n140, ZN => 
                           dp_ex_stage_alu_r60_n138);
   dp_ex_stage_alu_r60_U91 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n295, 
                           A2 => dp_ex_stage_alu_r60_n294, ZN => 
                           dp_ex_stage_alu_r60_n280);
   dp_ex_stage_alu_r60_U90 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r60_n282,
                           B2 => dp_ex_stage_alu_r60_n283, A => 
                           dp_ex_stage_alu_r60_n284, ZN => 
                           dp_ex_stage_alu_r60_n281);
   dp_ex_stage_alu_r60_U89 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n281,
                           A2 => dp_ex_stage_alu_r60_n280, ZN => 
                           dp_ex_stage_alu_r60_n253);
   dp_ex_stage_alu_r60_U88 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n119, 
                           A2 => dp_ex_stage_alu_r60_n120, ZN => 
                           dp_ex_stage_alu_r60_n118);
   dp_ex_stage_alu_r60_U87 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n23, 
                           A2 => dp_ex_stage_alu_r60_n184, ZN => 
                           dp_ex_stage_alu_r60_n70);
   dp_ex_stage_alu_r60_U86 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n293,
                           A2 => dp_ex_stage_alu_r60_n163, ZN => 
                           dp_ex_stage_alu_r60_n164);
   dp_ex_stage_alu_r60_U85 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n206,
                           A2 => dp_ex_stage_alu_r60_n74, ZN => 
                           dp_ex_stage_alu_r60_n184);
   dp_ex_stage_alu_r60_U84 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n166,
                           B2 => dp_ex_stage_alu_r60_n167, A => 
                           dp_ex_stage_alu_r60_n168, ZN => 
                           dp_ex_stage_alu_r60_n165);
   dp_ex_stage_alu_r60_U83 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n6, A2
                           => dp_ex_stage_alu_r60_n165, ZN => 
                           dp_ex_stage_alu_r60_n160);
   dp_ex_stage_alu_r60_U82 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n162,
                           A2 => dp_ex_stage_alu_r60_n163, ZN => 
                           dp_ex_stage_alu_r60_n161);
   dp_ex_stage_alu_r60_U81 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n160, 
                           A2 => dp_ex_stage_alu_r60_n161, ZN => 
                           dp_ex_stage_alu_r60_n146);
   dp_ex_stage_alu_r60_U80 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n5, A2
                           => dp_ex_stage_alu_r60_n136, ZN => 
                           dp_ex_stage_alu_r60_n260);
   dp_ex_stage_alu_r60_U79 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n171, 
                           A2 => dp_ex_stage_alu_r60_n173, ZN => 
                           dp_ex_stage_alu_r60_n294);
   dp_ex_stage_alu_r60_U78 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n159, 
                           A2 => dp_ex_stage_alu_r60_n9, ZN => 
                           dp_ex_stage_alu_r60_n153);
   dp_ex_stage_alu_r60_U77 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n58, 
                           A2 => dp_ex_stage_alu_r60_n59, ZN => 
                           dp_ex_stage_alu_r60_n57);
   dp_ex_stage_alu_r60_U76 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n290,
                           A2 => dp_ex_stage_alu_r60_n162, ZN => 
                           dp_ex_stage_alu_r60_n289);
   dp_ex_stage_alu_r60_U75 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n288, 
                           A2 => dp_ex_stage_alu_r60_n289, ZN => 
                           dp_ex_stage_alu_r60_n283);
   dp_ex_stage_alu_r60_U74 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n179, 
                           A2 => dp_ex_stage_alu_r60_n109, ZN => 
                           dp_ex_stage_alu_r60_n175);
   dp_ex_stage_alu_r60_U73 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n99, 
                           A2 => dp_ex_stage_alu_r60_n94, ZN => 
                           dp_ex_stage_alu_r60_n96);
   dp_ex_stage_alu_r60_U72 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n88, 
                           A2 => dp_ex_stage_alu_r60_n89, ZN => 
                           dp_ex_stage_alu_r60_n87);
   dp_ex_stage_alu_r60_U71 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n95, 
                           B2 => dp_ex_stage_alu_r60_n96, A => 
                           dp_ex_stage_alu_r60_n97, ZN => 
                           dp_ex_stage_alu_r60_n86);
   dp_ex_stage_alu_r60_U70 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n86, 
                           A2 => dp_ex_stage_alu_r60_n87, ZN => 
                           dp_ex_stage_alu_r60_n82);
   dp_ex_stage_alu_r60_U69 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n252,
                           A2 => dp_ex_stage_alu_r60_n123, ZN => 
                           dp_ex_stage_alu_r60_n181);
   dp_ex_stage_alu_r60_U68 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n273,
                           A2 => dp_ex_stage_alu_r60_n8, ZN => 
                           dp_ex_stage_alu_r60_n276);
   dp_ex_stage_alu_r60_U67 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n269,
                           A2 => dp_ex_stage_alu_r60_n268, ZN => 
                           dp_ex_stage_alu_r60_n267);
   dp_ex_stage_alu_r60_U66 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n159,
                           B2 => dp_ex_stage_alu_r60_n276, A => 
                           dp_ex_stage_alu_r60_n277, ZN => 
                           dp_ex_stage_alu_r60_n266);
   dp_ex_stage_alu_r60_U65 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n226,
                           A2 => dp_ex_stage_alu_r60_n94, ZN => 
                           dp_ex_stage_alu_r60_n91);
   dp_ex_stage_alu_r60_U64 : NAND4_X1 port map( A1 => dp_ex_stage_alu_r60_n99, 
                           A2 => dp_ex_stage_alu_r60_n111, A3 => 
                           dp_ex_stage_alu_r60_n94, A4 => 
                           dp_ex_stage_alu_r60_n112, ZN => 
                           dp_ex_stage_alu_r60_n103);
   dp_ex_stage_alu_r60_U63 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n178, 
                           A2 => dp_ex_stage_alu_r60_n179, ZN => 
                           dp_ex_stage_alu_r60_n243);
   dp_ex_stage_alu_r60_U62 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r60_n70, 
                           B2 => dp_ex_stage_alu_r60_n71, A => 
                           dp_ex_stage_alu_r60_n72, ZN => 
                           dp_ex_stage_alu_r60_n62);
   dp_ex_stage_alu_r60_U61 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n65, 
                           A2 => dp_ex_stage_alu_r60_n66, ZN => 
                           dp_ex_stage_alu_r60_n64);
   dp_ex_stage_alu_r60_U60 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n62, 
                           B2 => dp_ex_stage_alu_r60_n63, A => 
                           dp_ex_stage_alu_r60_n64, ZN => 
                           dp_ex_stage_alu_r60_n56);
   dp_ex_stage_alu_r60_U59 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n4, 
                           A2 => dp_ex_stage_alu_r60_n124, ZN => 
                           dp_ex_stage_alu_r60_n127);
   dp_ex_stage_alu_r60_U58 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n222,
                           A2 => dp_ex_stage_alu_r60_n85, ZN => 
                           dp_ex_stage_alu_r60_n98);
   dp_ex_stage_alu_r60_U57 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n296,
                           B2 => dp_ex_stage_alu_r60_n171, A => 
                           dp_ex_stage_alu_r60_n273, ZN => 
                           dp_ex_stage_alu_r60_n295);
   dp_ex_stage_alu_r60_U56 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r60_n81, 
                           B2 => dp_ex_stage_alu_r60_n82, A => 
                           dp_ex_stage_alu_r60_n83, ZN => 
                           dp_ex_stage_alu_r60_n75);
   dp_ex_stage_alu_r60_U55 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n78, 
                           A2 => dp_ex_stage_alu_r60_n24, ZN => 
                           dp_ex_stage_alu_r60_n77);
   dp_ex_stage_alu_r60_U54 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n75, 
                           B2 => dp_ex_stage_alu_r60_n76, A => 
                           dp_ex_stage_alu_r60_n77, ZN => 
                           dp_ex_stage_alu_r60_n71);
   dp_ex_stage_alu_r60_U53 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n198, 
                           A2 => dp_ex_stage_alu_r60_n199, ZN => 
                           dp_ex_stage_alu_r60_n197);
   dp_ex_stage_alu_r60_U52 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n178,
                           B2 => dp_ex_stage_alu_r60_n249, A => 
                           dp_ex_stage_alu_r60_n95, ZN => 
                           dp_ex_stage_alu_r60_n242);
   dp_ex_stage_alu_r60_U51 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n211, 
                           A2 => dp_ex_stage_alu_r60_n23, ZN => 
                           dp_ex_stage_alu_r60_n210);
   dp_ex_stage_alu_r60_U50 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n262,
                           A2 => dp_ex_stage_alu_r60_n129, ZN => 
                           dp_ex_stage_alu_r60_n144);
   dp_ex_stage_alu_r60_U49 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n271,
                           A2 => dp_ex_stage_alu_r60_n152, ZN => 
                           dp_ex_stage_alu_r60_n155);
   dp_ex_stage_alu_r60_U48 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n285,
                           A2 => dp_ex_stage_alu_r60_n157, ZN => 
                           dp_ex_stage_alu_r60_n171);
   dp_ex_stage_alu_r60_U47 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n245,
                           A2 => dp_ex_stage_alu_r60_n110, ZN => 
                           dp_ex_stage_alu_r60_n178);
   dp_ex_stage_alu_r60_U46 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n112,
                           A2 => dp_ex_stage_alu_r60_n232, ZN => 
                           dp_ex_stage_alu_r60_n105);
   dp_ex_stage_alu_r60_U45 : NOR3_X1 port map( A1 => dp_ex_stage_alu_r60_n156, 
                           A2 => dp_ex_stage_alu_r60_n155, A3 => 
                           dp_ex_stage_alu_r60_n157, ZN => 
                           dp_ex_stage_alu_r60_n154);
   dp_ex_stage_alu_r60_U44 : OAI22_X1 port map( A1 => dp_ex_stage_alu_r60_n105,
                           A2 => dp_ex_stage_alu_r60_n106, B1 => 
                           dp_ex_stage_alu_r60_n107, B2 => 
                           dp_ex_stage_alu_r60_n105, ZN => 
                           dp_ex_stage_alu_r60_n104);
   dp_ex_stage_alu_r60_U43 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n127, 
                           A2 => dp_ex_stage_alu_r60_n5, ZN => 
                           dp_ex_stage_alu_r60_n141);
   dp_ex_stage_alu_r60_U42 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n105, 
                           A2 => dp_ex_stage_alu_r60_n178, ZN => 
                           dp_ex_stage_alu_r60_n176);
   dp_ex_stage_alu_r60_U41 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n181, 
                           A2 => dp_ex_stage_alu_r60_n178, ZN => 
                           dp_ex_stage_alu_r60_n299);
   dp_ex_stage_alu_r60_U40 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n138, 
                           A2 => dp_ex_stage_alu_r60_n144, ZN => 
                           dp_ex_stage_alu_r60_n268);
   dp_ex_stage_alu_r60_U39 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n91, 
                           A2 => dp_ex_stage_alu_r60_n98, ZN => 
                           dp_ex_stage_alu_r60_n229);
   dp_ex_stage_alu_r60_U38 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n164, 
                           A2 => dp_ex_stage_alu_r60_n171, ZN => 
                           dp_ex_stage_alu_r60_n282);
   dp_ex_stage_alu_r60_U37 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n132,
                           A2 => dp_ex_stage_alu_r60_n133, ZN => 
                           dp_ex_stage_alu_r60_n131);
   dp_ex_stage_alu_r60_U36 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n130, 
                           A2 => dp_ex_stage_alu_r60_n131, ZN => 
                           dp_ex_stage_alu_r60_n114);
   dp_ex_stage_alu_r60_U35 : AOI21_X1 port map( B1 => dp_ex_stage_alu_r60_n113,
                           B2 => dp_ex_stage_alu_r60_n114, A => 
                           dp_ex_stage_alu_r60_n115, ZN => 
                           dp_ex_stage_alu_r60_n101);
   dp_ex_stage_alu_r60_U34 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n103, 
                           A2 => dp_ex_stage_alu_r60_n104, ZN => 
                           dp_ex_stage_alu_r60_n102);
   dp_ex_stage_alu_r60_U33 : OAI21_X1 port map( B1 => dp_ex_stage_alu_r60_n100,
                           B2 => dp_ex_stage_alu_r60_n101, A => 
                           dp_ex_stage_alu_r60_n102, ZN => 
                           dp_ex_stage_alu_r60_n81);
   dp_ex_stage_alu_r60_U32 : NAND4_X1 port map( A1 => dp_ex_stage_alu_r60_n299,
                           A2 => dp_ex_stage_alu_r60_n300, A3 => 
                           dp_ex_stage_alu_r60_n301, A4 => 
                           dp_ex_stage_alu_r60_n302, ZN => 
                           dp_ex_stage_alu_r60_n239);
   dp_ex_stage_alu_r60_U31 : NOR3_X1 port map( A1 => dp_ex_stage_alu_r60_n242, 
                           A2 => dp_ex_stage_alu_r60_n243, A3 => 
                           dp_ex_stage_alu_r60_n244, ZN => 
                           dp_ex_stage_alu_r60_n241);
   dp_ex_stage_alu_r60_U30 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n153, 
                           A2 => dp_ex_stage_alu_r60_n154, ZN => 
                           dp_ex_stage_alu_r60_n147);
   dp_ex_stage_alu_r60_U29 : NOR2_X1 port map( A1 => dp_ex_stage_alu_r60_n149, 
                           A2 => dp_ex_stage_alu_r60_n150, ZN => 
                           dp_ex_stage_alu_r60_n148);
   dp_ex_stage_alu_r60_U28 : OAI211_X1 port map( C1 => dp_ex_stage_alu_r60_n145
                           , C2 => dp_ex_stage_alu_r60_n146, A => 
                           dp_ex_stage_alu_r60_n147, B => 
                           dp_ex_stage_alu_r60_n148, ZN => 
                           dp_ex_stage_alu_r60_n113);
   dp_ex_stage_alu_r60_U27 : AND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_13_port, A2 => 
                           dp_ex_stage_alu_r60_n307, ZN => 
                           dp_ex_stage_alu_r60_n20);
   dp_ex_stage_alu_r60_U26 : AND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_2_port, A2 => 
                           dp_ex_stage_alu_r60_n28, ZN => 
                           dp_ex_stage_alu_r60_n19);
   dp_ex_stage_alu_r60_U25 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n190, 
                           A2 => dp_ex_stage_alu_r60_n189, ZN => 
                           dp_ex_stage_alu_N17_port);
   dp_ex_stage_alu_r60_U24 : OR2_X1 port map( A1 => dp_ex_stage_alu_n46, A2 => 
                           dp_ex_stage_alu_r60_n291, ZN => 
                           dp_ex_stage_alu_r60_n17);
   dp_ex_stage_alu_r60_U23 : OR2_X1 port map( A1 => dp_ex_stage_alu_n45, A2 => 
                           dp_ex_stage_alu_r60_n292, ZN => 
                           dp_ex_stage_alu_r60_n16);
   dp_ex_stage_alu_r60_U22 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n16, 
                           A2 => dp_ex_stage_alu_r60_n17, ZN => 
                           dp_ex_stage_alu_r60_n288);
   dp_ex_stage_alu_r60_U21 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_muxA_out_1_port, Z => 
                           dp_ex_stage_alu_r60_n15);
   dp_ex_stage_alu_r60_U20 : AND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_7_port, A2 => 
                           dp_ex_stage_alu_r60_n297, ZN => 
                           dp_ex_stage_alu_r60_n14);
   dp_ex_stage_alu_r60_U19 : AND2_X2 port map( A1 => 
                           dp_ex_stage_muxB_out_9_port, A2 => 
                           dp_ex_stage_alu_r60_n35, ZN => 
                           dp_ex_stage_alu_r60_n13);
   dp_ex_stage_alu_r60_U18 : OR2_X1 port map( A1 => dp_ex_stage_alu_r60_n286, 
                           A2 => dp_ex_stage_muxA_out_6_port, ZN => 
                           dp_ex_stage_alu_r60_n152);
   dp_ex_stage_alu_r60_U17 : CLKBUF_X1 port map( A => dp_ex_stage_alu_r60_n98, 
                           Z => dp_ex_stage_alu_r60_n12);
   dp_ex_stage_alu_r60_U16 : CLKBUF_X1 port map( A => dp_ex_stage_alu_r60_n140,
                           Z => dp_ex_stage_alu_r60_n11);
   dp_ex_stage_alu_r60_U15 : OR2_X1 port map( A1 => dp_ex_stage_alu_r60_n98, A2
                           => dp_ex_stage_alu_r60_n89, ZN => 
                           dp_ex_stage_alu_r60_n10);
   dp_ex_stage_alu_r60_U14 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n99, 
                           A2 => dp_ex_stage_alu_r60_n111, ZN => 
                           dp_ex_stage_alu_r60_n237);
   dp_ex_stage_alu_r60_U13 : INV_X1 port map( A => dp_ex_stage_alu_r60_n169, ZN
                           => dp_ex_stage_alu_r60_n9);
   dp_ex_stage_alu_r60_U12 : BUF_X1 port map( A => dp_ex_stage_alu_r60_n271, Z 
                           => dp_ex_stage_alu_r60_n8);
   dp_ex_stage_alu_r60_U11 : CLKBUF_X1 port map( A => dp_ex_stage_alu_r60_n164,
                           Z => dp_ex_stage_alu_r60_n6);
   dp_ex_stage_alu_r60_U10 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n262,
                           A2 => dp_ex_stage_alu_r60_n129, ZN => 
                           dp_ex_stage_alu_r60_n5);
   dp_ex_stage_alu_r60_U9 : NAND2_X1 port map( A1 => 
                           dp_ex_stage_muxA_out_12_port, A2 => 
                           dp_ex_stage_alu_r60_n308, ZN => 
                           dp_ex_stage_alu_r60_n4);
   dp_ex_stage_alu_r60_U8 : CLKBUF_X1 port map( A => dp_ex_stage_alu_n73, Z => 
                           dp_ex_stage_alu_r60_n7);
   dp_ex_stage_alu_r60_U7 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n186, 
                           A2 => dp_ex_stage_alu_r60_n187, ZN => 
                           dp_ex_stage_alu_r60_n3);
   dp_ex_stage_alu_r60_U6 : AND2_X1 port map( A1 => dp_ex_stage_alu_r60_n313, 
                           A2 => dp_ex_stage_alu_r60_n187, ZN => 
                           dp_ex_stage_alu_r60_n2);
   dp_ex_stage_alu_r60_U5 : INV_X1 port map( A => dp_ex_stage_muxB_out_25_port,
                           ZN => dp_ex_stage_alu_r60_n212);
   dp_ex_stage_alu_r60_U4 : NAND2_X1 port map( A1 => dp_ex_stage_alu_r60_n231, 
                           A2 => dp_ex_stage_alu_r60_n105, ZN => 
                           dp_ex_stage_alu_r60_n230);
   dp_ex_stage_alu_r60_U3 : INV_X1 port map( A => dp_ex_stage_alu_r60_n13, ZN 
                           => dp_ex_stage_alu_r60_n143);
   dp_ex_stage_alu_r60_U2 : INV_X1 port map( A => dp_ex_stage_alu_r60_n20, ZN 
                           => dp_ex_stage_alu_r60_n304);
   dp_ex_stage_alu_r60_U1 : CLKBUF_X1 port map( A => 
                           dp_ex_stage_muxB_out_4_port, Z => 
                           dp_ex_stage_alu_r60_n1);

end SYN_dlx_rtl;
